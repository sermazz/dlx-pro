

    module DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW_sra_0 ( 
        A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  AOI21_X1 U2 ( .B1(n217), .B2(n218), .A(n50), .ZN(n113) );
  AOI21_X1 U3 ( .B1(n189), .B2(n190), .A(n50), .ZN(n149) );
  AOI21_X1 U4 ( .B1(n203), .B2(n204), .A(n50), .ZN(n97) );
  AOI21_X1 U5 ( .B1(n234), .B2(n235), .A(n50), .ZN(n226) );
  NAND2_X1 U50 ( .A1(n45), .A2(n46), .ZN(B[9]) );
  AOI21_X1 U51 ( .B1(n47), .B2(n48), .A(n49), .ZN(n46) );
  OAI21_X1 U52 ( .B1(n260), .B2(n50), .A(n51), .ZN(n49) );
  NAND2_X1 U53 ( .A1(n288), .A2(n52), .ZN(n51) );
  AOI22_X1 U54 ( .A1(n54), .A2(n55), .B1(SH[4]), .B2(n56), .ZN(n45) );
  NAND2_X1 U55 ( .A1(n57), .A2(n58), .ZN(B[8]) );
  AOI21_X1 U56 ( .B1(n47), .B2(n59), .A(n60), .ZN(n58) );
  OAI21_X1 U57 ( .B1(n276), .B2(n61), .A(n62), .ZN(n60) );
  NAND2_X1 U58 ( .A1(n287), .A2(n63), .ZN(n62) );
  AOI22_X1 U59 ( .A1(n54), .A2(n64), .B1(SH[4]), .B2(n277), .ZN(n57) );
  NAND2_X1 U60 ( .A1(n66), .A2(n67), .ZN(B[7]) );
  AOI21_X1 U61 ( .B1(n248), .B2(n68), .A(n69), .ZN(n67) );
  OAI21_X1 U62 ( .B1(n269), .B2(n50), .A(n70), .ZN(n69) );
  NAND2_X1 U63 ( .A1(n288), .A2(n71), .ZN(n70) );
  AOI22_X1 U64 ( .A1(n250), .A2(n72), .B1(n255), .B2(n73), .ZN(n66) );
  NAND2_X1 U65 ( .A1(n74), .A2(n75), .ZN(B[6]) );
  AOI21_X1 U66 ( .B1(n248), .B2(n76), .A(n77), .ZN(n75) );
  OAI21_X1 U67 ( .B1(n282), .B2(n50), .A(n78), .ZN(n77) );
  NAND2_X1 U68 ( .A1(n288), .A2(n79), .ZN(n78) );
  AOI22_X1 U69 ( .A1(n250), .A2(n80), .B1(n255), .B2(n81), .ZN(n74) );
  NAND2_X1 U70 ( .A1(n82), .A2(n83), .ZN(B[5]) );
  AOI21_X1 U71 ( .B1(n47), .B2(n55), .A(n84), .ZN(n83) );
  OAI21_X1 U72 ( .B1(n265), .B2(n50), .A(n85), .ZN(n84) );
  NAND2_X1 U73 ( .A1(n288), .A2(n48), .ZN(n85) );
  AOI22_X1 U74 ( .A1(n54), .A2(n86), .B1(SH[4]), .B2(n87), .ZN(n82) );
  NAND2_X1 U75 ( .A1(n88), .A2(n89), .ZN(B[4]) );
  AOI21_X1 U76 ( .B1(n47), .B2(n64), .A(n90), .ZN(n89) );
  OAI21_X1 U77 ( .B1(n276), .B2(n50), .A(n91), .ZN(n90) );
  NAND2_X1 U78 ( .A1(n288), .A2(n59), .ZN(n91) );
  AOI22_X1 U79 ( .A1(n54), .A2(n93), .B1(SH[4]), .B2(n94), .ZN(n88) );
  NAND2_X1 U80 ( .A1(n95), .A2(n96), .ZN(B[3]) );
  NOR3_X1 U81 ( .A1(n97), .A2(n98), .A3(n99), .ZN(n96) );
  AOI21_X1 U83 ( .B1(n100), .B2(n101), .A(n290), .ZN(n98) );
  AOI22_X1 U84 ( .A1(A[5]), .A2(n254), .B1(A[6]), .B2(n253), .ZN(n101) );
  AOI22_X1 U85 ( .A1(A[4]), .A2(n252), .B1(A[3]), .B2(n251), .ZN(n100) );
  AOI22_X1 U86 ( .A1(n248), .A2(n72), .B1(n255), .B2(n106), .ZN(n95) );
  NAND2_X1 U87 ( .A1(n107), .A2(n108), .ZN(n72) );
  AOI22_X1 U88 ( .A1(A[9]), .A2(n254), .B1(A[10]), .B2(n103), .ZN(n108) );
  AOI22_X1 U89 ( .A1(A[8]), .A2(n252), .B1(A[7]), .B2(n105), .ZN(n107) );
  OAI21_X1 U90 ( .B1(n255), .B2(n109), .A(n110), .ZN(B[30]) );
  NAND2_X1 U91 ( .A1(n111), .A2(n112), .ZN(B[2]) );
  NOR3_X1 U92 ( .A1(n113), .A2(n114), .A3(n115), .ZN(n112) );
  AOI21_X1 U94 ( .B1(n116), .B2(n117), .A(n290), .ZN(n114) );
  AOI22_X1 U95 ( .A1(A[4]), .A2(n254), .B1(A[5]), .B2(n103), .ZN(n117) );
  AOI22_X1 U96 ( .A1(A[3]), .A2(n104), .B1(A[2]), .B2(n105), .ZN(n116) );
  AOI22_X1 U97 ( .A1(n248), .A2(n80), .B1(n255), .B2(n118), .ZN(n111) );
  NAND2_X1 U98 ( .A1(n119), .A2(n120), .ZN(n80) );
  AOI22_X1 U99 ( .A1(A[8]), .A2(n254), .B1(A[9]), .B2(n103), .ZN(n120) );
  AOI22_X1 U100 ( .A1(A[7]), .A2(n252), .B1(A[6]), .B2(n105), .ZN(n119) );
  OAI21_X1 U101 ( .B1(n255), .B2(n121), .A(n110), .ZN(B[29]) );
  OAI21_X1 U102 ( .B1(n255), .B2(n122), .A(n110), .ZN(B[28]) );
  OAI21_X1 U103 ( .B1(n255), .B2(n123), .A(n110), .ZN(B[27]) );
  OAI21_X1 U104 ( .B1(n255), .B2(n280), .A(n110), .ZN(B[26]) );
  OAI21_X1 U105 ( .B1(n255), .B2(n263), .A(n110), .ZN(B[25]) );
  OAI21_X1 U106 ( .B1(n264), .B2(n291), .A(n125), .ZN(n56) );
  AOI21_X1 U107 ( .B1(n126), .B2(n127), .A(n286), .ZN(n125) );
  OAI21_X1 U108 ( .B1(n255), .B2(n65), .A(n110), .ZN(B[24]) );
  AOI21_X1 U109 ( .B1(n128), .B2(n129), .A(n130), .ZN(n65) );
  OAI21_X1 U110 ( .B1(n289), .B2(n278), .A(n131), .ZN(n130) );
  OAI21_X1 U111 ( .B1(n255), .B2(n266), .A(n110), .ZN(B[23]) );
  OAI21_X1 U112 ( .B1(n267), .B2(n291), .A(n133), .ZN(n73) );
  AOI21_X1 U113 ( .B1(n126), .B2(n134), .A(n286), .ZN(n133) );
  OAI21_X1 U114 ( .B1(n255), .B2(n272), .A(n110), .ZN(B[22]) );
  NAND2_X1 U115 ( .A1(n135), .A2(n136), .ZN(n81) );
  AOI21_X1 U116 ( .B1(n137), .B2(n138), .A(n139), .ZN(n136) );
  AOI22_X1 U117 ( .A1(n126), .A2(n140), .B1(n249), .B2(n141), .ZN(n135) );
  OAI21_X1 U118 ( .B1(n255), .B2(n262), .A(n110), .ZN(B[21]) );
  NAND2_X1 U119 ( .A1(n142), .A2(n143), .ZN(n87) );
  AOI21_X1 U120 ( .B1(n137), .B2(n127), .A(n139), .ZN(n143) );
  AOI22_X1 U121 ( .A1(n126), .A2(n144), .B1(n249), .B2(n53), .ZN(n142) );
  OAI21_X1 U122 ( .B1(n255), .B2(n275), .A(n110), .ZN(B[20]) );
  NAND2_X1 U123 ( .A1(n145), .A2(n146), .ZN(n94) );
  AOI21_X1 U124 ( .B1(n137), .B2(n132), .A(n139), .ZN(n146) );
  AOI22_X1 U125 ( .A1(n126), .A2(n128), .B1(n249), .B2(n63), .ZN(n145) );
  NAND2_X1 U126 ( .A1(n147), .A2(n148), .ZN(B[1]) );
  NOR3_X1 U127 ( .A1(n149), .A2(n150), .A3(n151), .ZN(n148) );
  NAND2_X1 U129 ( .A1(n152), .A2(n153), .ZN(n55) );
  AOI22_X1 U130 ( .A1(A[11]), .A2(n254), .B1(A[12]), .B2(n103), .ZN(n153) );
  AOI22_X1 U131 ( .A1(A[10]), .A2(n104), .B1(A[9]), .B2(n105), .ZN(n152) );
  AOI21_X1 U132 ( .B1(n154), .B2(n155), .A(n290), .ZN(n150) );
  AOI22_X1 U133 ( .A1(A[3]), .A2(n254), .B1(A[4]), .B2(n103), .ZN(n155) );
  AOI22_X1 U134 ( .A1(A[2]), .A2(n252), .B1(A[1]), .B2(n105), .ZN(n154) );
  AOI22_X1 U135 ( .A1(n47), .A2(n86), .B1(SH[4]), .B2(n156), .ZN(n147) );
  NAND2_X1 U136 ( .A1(n157), .A2(n158), .ZN(n86) );
  AOI22_X1 U137 ( .A1(A[7]), .A2(n254), .B1(A[8]), .B2(n103), .ZN(n158) );
  AOI22_X1 U138 ( .A1(A[6]), .A2(n104), .B1(A[5]), .B2(n105), .ZN(n157) );
  OAI21_X1 U139 ( .B1(n255), .B2(n268), .A(n110), .ZN(B[19]) );
  NAND2_X1 U140 ( .A1(n159), .A2(n160), .ZN(n106) );
  AOI21_X1 U141 ( .B1(n137), .B2(n134), .A(n139), .ZN(n160) );
  NOR2_X1 U142 ( .A1(n131), .A2(n257), .ZN(n139) );
  AOI22_X1 U143 ( .A1(n126), .A2(n161), .B1(n249), .B2(n162), .ZN(n159) );
  OAI21_X1 U144 ( .B1(n255), .B2(n271), .A(n110), .ZN(B[18]) );
  NAND2_X1 U145 ( .A1(n163), .A2(n164), .ZN(n118) );
  AOI22_X1 U146 ( .A1(n165), .A2(n138), .B1(n137), .B2(n140), .ZN(n164) );
  AOI22_X1 U147 ( .A1(n126), .A2(n141), .B1(n249), .B2(n166), .ZN(n163) );
  OAI21_X1 U148 ( .B1(n255), .B2(n261), .A(n110), .ZN(B[17]) );
  NAND2_X1 U149 ( .A1(n167), .A2(n168), .ZN(n156) );
  AOI22_X1 U150 ( .A1(n165), .A2(n127), .B1(n137), .B2(n144), .ZN(n168) );
  AOI22_X1 U151 ( .A1(n126), .A2(n53), .B1(n249), .B2(n52), .ZN(n167) );
  OAI21_X1 U152 ( .B1(n255), .B2(n274), .A(n110), .ZN(B[16]) );
  NAND2_X1 U153 ( .A1(n170), .A2(n171), .ZN(B[15]) );
  AOI21_X1 U154 ( .B1(n287), .B2(n134), .A(n172), .ZN(n171) );
  OAI21_X1 U155 ( .B1(n267), .B2(n61), .A(n110), .ZN(n172) );
  NAND2_X1 U156 ( .A1(n255), .A2(\A[31] ), .ZN(n110) );
  AOI22_X1 U157 ( .A1(n47), .A2(n162), .B1(n250), .B2(n71), .ZN(n170) );
  NAND2_X1 U158 ( .A1(n173), .A2(n174), .ZN(B[14]) );
  AOI21_X1 U159 ( .B1(n248), .B2(n166), .A(n175), .ZN(n174) );
  OAI21_X1 U160 ( .B1(n281), .B2(n50), .A(n176), .ZN(n175) );
  NAND2_X1 U161 ( .A1(n288), .A2(n141), .ZN(n176) );
  AOI22_X1 U162 ( .A1(n250), .A2(n79), .B1(SH[4]), .B2(n284), .ZN(n173) );
  AOI21_X1 U163 ( .B1(n138), .B2(n129), .A(n177), .ZN(n109) );
  NAND2_X1 U164 ( .A1(n178), .A2(n179), .ZN(B[13]) );
  AOI21_X1 U165 ( .B1(n248), .B2(n52), .A(n180), .ZN(n179) );
  OAI21_X1 U166 ( .B1(n264), .B2(n50), .A(n181), .ZN(n180) );
  NAND2_X1 U167 ( .A1(n288), .A2(n53), .ZN(n181) );
  NAND2_X1 U168 ( .A1(n182), .A2(n183), .ZN(n53) );
  AOI22_X1 U169 ( .A1(A[23]), .A2(n254), .B1(A[24]), .B2(n103), .ZN(n183) );
  AOI22_X1 U170 ( .A1(A[22]), .A2(n252), .B1(A[21]), .B2(n105), .ZN(n182) );
  NAND2_X1 U171 ( .A1(n184), .A2(n185), .ZN(n144) );
  AOI22_X1 U172 ( .A1(A[27]), .A2(n254), .B1(A[28]), .B2(n103), .ZN(n185) );
  AOI22_X1 U173 ( .A1(A[26]), .A2(n252), .B1(A[25]), .B2(n251), .ZN(n184) );
  NAND2_X1 U174 ( .A1(n186), .A2(n187), .ZN(n52) );
  AOI22_X1 U175 ( .A1(A[19]), .A2(n254), .B1(A[20]), .B2(n103), .ZN(n187) );
  AOI22_X1 U176 ( .A1(A[18]), .A2(n252), .B1(A[17]), .B2(n105), .ZN(n186) );
  AOI22_X1 U177 ( .A1(n250), .A2(n48), .B1(n255), .B2(n283), .ZN(n178) );
  AOI21_X1 U178 ( .B1(n127), .B2(n249), .A(n177), .ZN(n121) );
  OAI21_X1 U179 ( .B1(n258), .B2(n285), .A(n188), .ZN(n127) );
  AOI22_X1 U180 ( .A1(A[30]), .A2(n252), .B1(A[29]), .B2(n105), .ZN(n188) );
  NAND2_X1 U181 ( .A1(n189), .A2(n190), .ZN(n48) );
  AOI22_X1 U182 ( .A1(A[15]), .A2(n254), .B1(A[16]), .B2(n103), .ZN(n190) );
  AOI22_X1 U183 ( .A1(A[14]), .A2(n104), .B1(A[13]), .B2(n105), .ZN(n189) );
  NAND2_X1 U184 ( .A1(n191), .A2(n192), .ZN(B[12]) );
  AOI21_X1 U185 ( .B1(n47), .B2(n92), .A(n193), .ZN(n192) );
  OAI21_X1 U186 ( .B1(n273), .B2(n61), .A(n194), .ZN(n193) );
  NAND2_X1 U187 ( .A1(n287), .A2(n128), .ZN(n194) );
  AOI22_X1 U188 ( .A1(n54), .A2(n59), .B1(SH[4]), .B2(n279), .ZN(n191) );
  AOI21_X1 U189 ( .B1(n132), .B2(n249), .A(n177), .ZN(n122) );
  NAND2_X1 U190 ( .A1(n195), .A2(n196), .ZN(B[11]) );
  AOI21_X1 U191 ( .B1(n47), .B2(n71), .A(n197), .ZN(n196) );
  OAI21_X1 U192 ( .B1(n269), .B2(n61), .A(n198), .ZN(n197) );
  NAND2_X1 U193 ( .A1(n287), .A2(n161), .ZN(n198) );
  NAND2_X1 U194 ( .A1(n199), .A2(n200), .ZN(n161) );
  AOI22_X1 U195 ( .A1(A[25]), .A2(n254), .B1(A[26]), .B2(n253), .ZN(n200) );
  AOI22_X1 U196 ( .A1(A[24]), .A2(n104), .B1(A[23]), .B2(n105), .ZN(n199) );
  NAND2_X1 U197 ( .A1(n201), .A2(n202), .ZN(n162) );
  AOI22_X1 U198 ( .A1(A[21]), .A2(n102), .B1(A[22]), .B2(n253), .ZN(n202) );
  AOI22_X1 U199 ( .A1(n104), .A2(A[20]), .B1(n251), .B2(A[19]), .ZN(n201) );
  NAND2_X1 U200 ( .A1(n203), .A2(n204), .ZN(n71) );
  AOI22_X1 U201 ( .A1(A[17]), .A2(n254), .B1(A[18]), .B2(n253), .ZN(n204) );
  AOI22_X1 U202 ( .A1(A[16]), .A2(n252), .B1(A[15]), .B2(n251), .ZN(n203) );
  AOI22_X1 U203 ( .A1(n54), .A2(n68), .B1(SH[4]), .B2(n270), .ZN(n195) );
  AOI21_X1 U204 ( .B1(n134), .B2(n249), .A(n177), .ZN(n123) );
  OAI21_X1 U205 ( .B1(n257), .B2(n285), .A(n131), .ZN(n177) );
  NAND2_X1 U206 ( .A1(n205), .A2(n206), .ZN(n134) );
  AOI22_X1 U207 ( .A1(A[29]), .A2(n102), .B1(A[30]), .B2(n253), .ZN(n206) );
  AOI22_X1 U208 ( .A1(A[28]), .A2(n252), .B1(A[27]), .B2(n251), .ZN(n205) );
  NAND2_X1 U209 ( .A1(n207), .A2(n208), .ZN(n68) );
  AOI22_X1 U210 ( .A1(A[13]), .A2(n254), .B1(A[14]), .B2(n253), .ZN(n208) );
  AOI22_X1 U211 ( .A1(A[12]), .A2(n252), .B1(A[11]), .B2(n251), .ZN(n207) );
  NAND2_X1 U212 ( .A1(n209), .A2(n210), .ZN(B[10]) );
  AOI21_X1 U213 ( .B1(n248), .B2(n79), .A(n211), .ZN(n210) );
  OAI21_X1 U214 ( .B1(n282), .B2(n61), .A(n212), .ZN(n211) );
  NAND2_X1 U215 ( .A1(n287), .A2(n141), .ZN(n212) );
  NAND2_X1 U216 ( .A1(n213), .A2(n214), .ZN(n141) );
  AOI22_X1 U217 ( .A1(A[24]), .A2(n102), .B1(A[25]), .B2(n253), .ZN(n214) );
  AOI22_X1 U218 ( .A1(A[23]), .A2(n252), .B1(A[22]), .B2(n251), .ZN(n213) );
  NAND2_X1 U219 ( .A1(n215), .A2(n216), .ZN(n166) );
  AOI22_X1 U220 ( .A1(A[20]), .A2(n102), .B1(A[21]), .B2(n253), .ZN(n216) );
  AOI22_X1 U221 ( .A1(n104), .A2(A[19]), .B1(n251), .B2(A[18]), .ZN(n215) );
  NAND2_X1 U222 ( .A1(n217), .A2(n218), .ZN(n79) );
  AOI22_X1 U223 ( .A1(A[16]), .A2(n254), .B1(A[17]), .B2(n253), .ZN(n218) );
  AOI22_X1 U224 ( .A1(A[15]), .A2(n252), .B1(A[14]), .B2(n251), .ZN(n217) );
  AOI22_X1 U225 ( .A1(n250), .A2(n76), .B1(n255), .B2(n124), .ZN(n209) );
  OAI21_X1 U226 ( .B1(n281), .B2(n291), .A(n219), .ZN(n124) );
  AOI21_X1 U227 ( .B1(n126), .B2(n138), .A(n286), .ZN(n219) );
  NAND2_X1 U228 ( .A1(\A[31] ), .A2(SH[3]), .ZN(n131) );
  MUX2_X2 U229 ( .A(\A[31] ), .B(A[30]), .S(n251), .Z(n138) );
  NAND2_X1 U230 ( .A1(n220), .A2(n221), .ZN(n140) );
  AOI22_X1 U231 ( .A1(A[28]), .A2(n102), .B1(A[29]), .B2(n253), .ZN(n221) );
  AOI22_X1 U232 ( .A1(A[27]), .A2(n252), .B1(A[26]), .B2(n251), .ZN(n220) );
  NAND2_X1 U233 ( .A1(n222), .A2(n223), .ZN(n76) );
  AOI22_X1 U234 ( .A1(A[12]), .A2(n254), .B1(A[13]), .B2(n253), .ZN(n223) );
  AOI22_X1 U235 ( .A1(A[11]), .A2(n252), .B1(A[10]), .B2(n251), .ZN(n222) );
  NAND2_X1 U236 ( .A1(n224), .A2(n225), .ZN(B[0]) );
  NOR3_X1 U237 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n225) );
  NAND2_X1 U239 ( .A1(n229), .A2(n257), .ZN(n61) );
  NAND2_X1 U240 ( .A1(n230), .A2(n231), .ZN(n64) );
  AOI22_X1 U241 ( .A1(A[10]), .A2(n102), .B1(A[11]), .B2(n253), .ZN(n231) );
  AOI22_X1 U242 ( .A1(A[9]), .A2(n104), .B1(A[8]), .B2(n251), .ZN(n230) );
  AOI21_X1 U243 ( .B1(n232), .B2(n233), .A(n290), .ZN(n227) );
  NOR2_X1 U244 ( .A1(n291), .A2(n255), .ZN(n54) );
  AOI22_X1 U245 ( .A1(A[2]), .A2(n254), .B1(A[3]), .B2(n253), .ZN(n233) );
  AOI22_X1 U246 ( .A1(A[1]), .A2(n104), .B1(A[0]), .B2(n251), .ZN(n232) );
  NAND2_X1 U247 ( .A1(SH[2]), .A2(n229), .ZN(n50) );
  NOR2_X1 U248 ( .A1(n256), .A2(n255), .ZN(n229) );
  NAND2_X1 U249 ( .A1(n234), .A2(n235), .ZN(n59) );
  AOI22_X1 U250 ( .A1(A[14]), .A2(n102), .B1(A[15]), .B2(n253), .ZN(n235) );
  AOI22_X1 U251 ( .A1(A[13]), .A2(n104), .B1(A[12]), .B2(n251), .ZN(n234) );
  AOI22_X1 U252 ( .A1(n248), .A2(n93), .B1(n255), .B2(n169), .ZN(n224) );
  NAND2_X1 U253 ( .A1(n236), .A2(n237), .ZN(n169) );
  AOI22_X1 U254 ( .A1(n165), .A2(n132), .B1(n137), .B2(n128), .ZN(n237) );
  NAND2_X1 U255 ( .A1(n238), .A2(n239), .ZN(n128) );
  AOI22_X1 U256 ( .A1(A[26]), .A2(n254), .B1(A[27]), .B2(n253), .ZN(n239) );
  AOI22_X1 U257 ( .A1(A[25]), .A2(n252), .B1(A[24]), .B2(n251), .ZN(n238) );
  NOR2_X1 U258 ( .A1(n256), .A2(SH[2]), .ZN(n137) );
  NAND2_X1 U259 ( .A1(n240), .A2(n241), .ZN(n132) );
  AOI22_X1 U260 ( .A1(A[30]), .A2(n102), .B1(\A[31] ), .B2(n253), .ZN(n241) );
  AOI22_X1 U261 ( .A1(A[29]), .A2(n252), .B1(A[28]), .B2(n251), .ZN(n240) );
  NOR2_X1 U262 ( .A1(n257), .A2(n256), .ZN(n165) );
  AOI22_X1 U263 ( .A1(n126), .A2(n63), .B1(n249), .B2(n92), .ZN(n236) );
  NAND2_X1 U264 ( .A1(n242), .A2(n243), .ZN(n92) );
  AOI22_X1 U265 ( .A1(A[18]), .A2(n102), .B1(n103), .B2(A[19]), .ZN(n243) );
  AOI22_X1 U266 ( .A1(A[17]), .A2(n252), .B1(A[16]), .B2(n251), .ZN(n242) );
  NOR2_X1 U267 ( .A1(SH[2]), .A2(SH[3]), .ZN(n129) );
  NAND2_X1 U268 ( .A1(n244), .A2(n245), .ZN(n63) );
  AOI22_X1 U269 ( .A1(A[22]), .A2(n102), .B1(A[23]), .B2(n253), .ZN(n245) );
  AOI22_X1 U270 ( .A1(A[21]), .A2(n252), .B1(n251), .B2(A[20]), .ZN(n244) );
  NAND2_X1 U271 ( .A1(n246), .A2(n247), .ZN(n93) );
  AOI22_X1 U272 ( .A1(A[6]), .A2(n102), .B1(A[7]), .B2(n253), .ZN(n247) );
  NOR2_X1 U273 ( .A1(n259), .A2(n258), .ZN(n103) );
  NOR2_X1 U274 ( .A1(n258), .A2(SH[0]), .ZN(n102) );
  AOI22_X1 U275 ( .A1(A[5]), .A2(n104), .B1(A[4]), .B2(n251), .ZN(n246) );
  NOR2_X1 U276 ( .A1(SH[0]), .A2(SH[1]), .ZN(n105) );
  NOR2_X1 U277 ( .A1(n259), .A2(SH[1]), .ZN(n104) );
  NOR2_X1 U278 ( .A1(n289), .A2(n255), .ZN(n47) );
  NOR2_X1 U279 ( .A1(n257), .A2(SH[3]), .ZN(n126) );
  AOI21_X1 U6 ( .B1(n222), .B2(n223), .A(n61), .ZN(n115) );
  AOI21_X1 U7 ( .B1(n152), .B2(n153), .A(n61), .ZN(n151) );
  AOI21_X1 U8 ( .B1(n207), .B2(n208), .A(n61), .ZN(n99) );
  AOI21_X1 U9 ( .B1(n230), .B2(n231), .A(n61), .ZN(n228) );
  INV_X1 U10 ( .A(n250), .ZN(n290) );
  INV_X1 U11 ( .A(n61), .ZN(n288) );
  CLKBUF_X1 U12 ( .A(n103), .Z(n253) );
  CLKBUF_X1 U13 ( .A(n47), .Z(n248) );
  CLKBUF_X1 U14 ( .A(n54), .Z(n250) );
  INV_X1 U15 ( .A(n129), .ZN(n291) );
  INV_X1 U16 ( .A(n122), .ZN(n279) );
  INV_X1 U17 ( .A(n65), .ZN(n277) );
  INV_X1 U18 ( .A(n73), .ZN(n266) );
  INV_X1 U19 ( .A(n56), .ZN(n263) );
  INV_X1 U20 ( .A(n124), .ZN(n280) );
  INV_X1 U21 ( .A(n126), .ZN(n289) );
  INV_X1 U22 ( .A(n156), .ZN(n261) );
  INV_X1 U23 ( .A(n87), .ZN(n262) );
  INV_X1 U24 ( .A(n118), .ZN(n271) );
  INV_X1 U25 ( .A(n81), .ZN(n272) );
  INV_X1 U26 ( .A(n106), .ZN(n268) );
  INV_X1 U27 ( .A(n132), .ZN(n278) );
  CLKBUF_X1 U28 ( .A(n105), .Z(n251) );
  INV_X1 U29 ( .A(n121), .ZN(n283) );
  INV_X1 U30 ( .A(n109), .ZN(n284) );
  INV_X1 U31 ( .A(n123), .ZN(n270) );
  CLKBUF_X1 U32 ( .A(n102), .Z(n254) );
  CLKBUF_X1 U33 ( .A(n104), .Z(n252) );
  INV_X1 U34 ( .A(n53), .ZN(n260) );
  INV_X1 U35 ( .A(n52), .ZN(n265) );
  INV_X1 U36 ( .A(n94), .ZN(n275) );
  INV_X1 U37 ( .A(n169), .ZN(n274) );
  CLKBUF_X1 U38 ( .A(n129), .Z(n249) );
  INV_X1 U39 ( .A(n50), .ZN(n287) );
  INV_X1 U40 ( .A(n131), .ZN(n286) );
  INV_X1 U41 ( .A(n161), .ZN(n267) );
  INV_X1 U42 ( .A(n140), .ZN(n281) );
  INV_X1 U43 ( .A(n144), .ZN(n264) );
  INV_X1 U44 ( .A(n92), .ZN(n276) );
  INV_X1 U45 ( .A(n162), .ZN(n269) );
  INV_X1 U46 ( .A(n166), .ZN(n282) );
  INV_X1 U47 ( .A(n63), .ZN(n273) );
  CLKBUF_X1 U48 ( .A(SH[4]), .Z(n255) );
  INV_X1 U49 ( .A(\A[31] ), .ZN(n285) );
  INV_X1 U82 ( .A(SH[3]), .ZN(n256) );
  INV_X1 U93 ( .A(SH[2]), .ZN(n257) );
  INV_X1 U128 ( .A(SH[1]), .ZN(n258) );
  INV_X1 U238 ( .A(SH[0]), .ZN(n259) );
endmodule



    module DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW_rash_0 ( 
        A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n249, n251, n253, n254, n255, n256, n259, n260, n261,
         n262, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275;

  AOI21_X1 U3 ( .B1(n211), .B2(n212), .A(n45), .ZN(n110) );
  AOI21_X1 U4 ( .B1(n137), .B2(n138), .A(n45), .ZN(n136) );
  AOI21_X1 U5 ( .B1(n193), .B2(n194), .A(n45), .ZN(n93) );
  AOI21_X1 U6 ( .B1(n219), .B2(n220), .A(n45), .ZN(n217) );
  NAND2_X1 U7 ( .A1(n242), .A2(n88), .ZN(n1) );
  NAND2_X1 U9 ( .A1(n242), .A2(n82), .ZN(n2) );
  NAND2_X1 U11 ( .A1(n242), .A2(n76), .ZN(n3) );
  NAND2_X1 U13 ( .A1(n242), .A2(n68), .ZN(n4) );
  AOI21_X1 U15 ( .B1(n225), .B2(n226), .A(SH[4]), .ZN(B[16]) );
  AOI21_X1 U16 ( .B1(n152), .B2(n153), .A(SH[4]), .ZN(B[17]) );
  AOI21_X1 U17 ( .B1(n147), .B2(n148), .A(SH[4]), .ZN(B[18]) );
  NAND2_X1 U18 ( .A1(n242), .A2(n101), .ZN(n5) );
  NAND2_X1 U20 ( .A1(n242), .A2(n59), .ZN(n6) );
  NAND2_X1 U22 ( .A1(n242), .A2(n50), .ZN(n7) );
  NAND2_X1 U56 ( .A1(n40), .A2(n41), .ZN(B[9]) );
  AOI21_X1 U57 ( .B1(n42), .B2(n43), .A(n44), .ZN(n41) );
  OAI21_X1 U58 ( .B1(n261), .B2(n45), .A(n46), .ZN(n44) );
  NAND2_X1 U59 ( .A1(n270), .A2(n47), .ZN(n46) );
  AOI22_X1 U60 ( .A1(n273), .A2(n49), .B1(SH[4]), .B2(n50), .ZN(n40) );
  NAND2_X1 U61 ( .A1(n51), .A2(n52), .ZN(B[8]) );
  AOI21_X1 U62 ( .B1(n42), .B2(n53), .A(n54), .ZN(n52) );
  OAI21_X1 U63 ( .B1(n260), .B2(n55), .A(n56), .ZN(n54) );
  NAND2_X1 U64 ( .A1(n271), .A2(n57), .ZN(n56) );
  AOI22_X1 U65 ( .A1(n273), .A2(n58), .B1(SH[4]), .B2(n59), .ZN(n51) );
  NAND2_X1 U66 ( .A1(n60), .A2(n61), .ZN(B[7]) );
  AOI21_X1 U67 ( .B1(n237), .B2(n62), .A(n63), .ZN(n61) );
  OAI21_X1 U68 ( .B1(n247), .B2(n55), .A(n64), .ZN(n63) );
  NAND2_X1 U69 ( .A1(n271), .A2(n65), .ZN(n64) );
  AOI22_X1 U70 ( .A1(n273), .A2(n67), .B1(SH[4]), .B2(n68), .ZN(n60) );
  NAND2_X1 U71 ( .A1(n69), .A2(n70), .ZN(B[6]) );
  AOI21_X1 U72 ( .B1(n42), .B2(n71), .A(n72), .ZN(n70) );
  OAI21_X1 U73 ( .B1(n254), .B2(n55), .A(n73), .ZN(n72) );
  NAND2_X1 U74 ( .A1(n271), .A2(n74), .ZN(n73) );
  AOI22_X1 U75 ( .A1(n273), .A2(n75), .B1(SH[4]), .B2(n76), .ZN(n69) );
  NAND2_X1 U76 ( .A1(n77), .A2(n78), .ZN(B[5]) );
  AOI21_X1 U77 ( .B1(n237), .B2(n49), .A(n79), .ZN(n78) );
  OAI21_X1 U78 ( .B1(n262), .B2(n45), .A(n80), .ZN(n79) );
  NAND2_X1 U79 ( .A1(n270), .A2(n48), .ZN(n80) );
  AOI22_X1 U80 ( .A1(n273), .A2(n81), .B1(SH[4]), .B2(n82), .ZN(n77) );
  NAND2_X1 U81 ( .A1(n83), .A2(n84), .ZN(B[4]) );
  AOI21_X1 U82 ( .B1(n237), .B2(n58), .A(n85), .ZN(n84) );
  OAI21_X1 U83 ( .B1(n256), .B2(n45), .A(n86), .ZN(n85) );
  NAND2_X1 U84 ( .A1(n270), .A2(n57), .ZN(n86) );
  AOI22_X1 U85 ( .A1(n273), .A2(n87), .B1(SH[4]), .B2(n88), .ZN(n83) );
  NAND2_X1 U86 ( .A1(n89), .A2(n90), .ZN(B[3]) );
  NOR3_X1 U87 ( .A1(n91), .A2(n92), .A3(n93), .ZN(n90) );
  AOI21_X1 U88 ( .B1(n94), .B2(n95), .A(n96), .ZN(n92) );
  AOI22_X1 U89 ( .A1(A[6]), .A2(n241), .B1(A[5]), .B2(n240), .ZN(n95) );
  AOI22_X1 U90 ( .A1(A[4]), .A2(n239), .B1(A[3]), .B2(n238), .ZN(n94) );
  AOI22_X1 U92 ( .A1(n237), .A2(n67), .B1(SH[4]), .B2(n101), .ZN(n89) );
  NAND2_X1 U93 ( .A1(n102), .A2(n103), .ZN(n67) );
  AOI22_X1 U94 ( .A1(A[10]), .A2(n241), .B1(A[9]), .B2(n98), .ZN(n103) );
  AOI22_X1 U95 ( .A1(A[8]), .A2(n239), .B1(A[7]), .B2(n100), .ZN(n102) );
  NOR2_X1 U96 ( .A1(n96), .A2(n104), .ZN(B[31]) );
  NOR2_X1 U97 ( .A1(n105), .A2(n96), .ZN(B[30]) );
  NAND2_X1 U98 ( .A1(n106), .A2(n107), .ZN(B[2]) );
  NOR3_X1 U99 ( .A1(n108), .A2(n109), .A3(n110), .ZN(n107) );
  AOI21_X1 U100 ( .B1(n111), .B2(n112), .A(n96), .ZN(n109) );
  AOI22_X1 U101 ( .A1(A[5]), .A2(n241), .B1(A[4]), .B2(n98), .ZN(n112) );
  AOI22_X1 U102 ( .A1(A[3]), .A2(n239), .B1(A[2]), .B2(n100), .ZN(n111) );
  AOI22_X1 U104 ( .A1(n42), .A2(n75), .B1(SH[4]), .B2(n113), .ZN(n106) );
  NAND2_X1 U105 ( .A1(n114), .A2(n115), .ZN(n75) );
  AOI22_X1 U106 ( .A1(A[9]), .A2(n241), .B1(A[8]), .B2(n98), .ZN(n115) );
  AOI22_X1 U107 ( .A1(A[7]), .A2(n239), .B1(A[6]), .B2(n100), .ZN(n114) );
  NOR2_X1 U108 ( .A1(n116), .A2(n96), .ZN(B[29]) );
  NOR2_X1 U109 ( .A1(n259), .A2(n96), .ZN(B[28]) );
  NOR3_X1 U110 ( .A1(n249), .A2(SH[4]), .A3(SH[3]), .ZN(B[27]) );
  NOR2_X1 U111 ( .A1(SH[4]), .A2(n117), .ZN(B[26]) );
  OAI21_X1 U112 ( .B1(n116), .B2(n118), .A(n119), .ZN(n50) );
  NAND2_X1 U113 ( .A1(n274), .A2(n120), .ZN(n119) );
  OAI21_X1 U114 ( .B1(n259), .B2(n118), .A(n121), .ZN(n59) );
  NAND2_X1 U115 ( .A1(n274), .A2(n122), .ZN(n121) );
  OAI21_X1 U116 ( .B1(n251), .B2(n124), .A(n125), .ZN(n68) );
  AOI22_X1 U117 ( .A1(n126), .A2(n269), .B1(n275), .B2(n127), .ZN(n125) );
  OAI21_X1 U118 ( .B1(n253), .B2(n124), .A(n128), .ZN(n76) );
  AOI22_X1 U119 ( .A1(n126), .A2(n266), .B1(n275), .B2(n129), .ZN(n128) );
  OAI21_X1 U120 ( .B1(n265), .B2(n124), .A(n130), .ZN(n82) );
  AOI22_X1 U121 ( .A1(n126), .A2(n267), .B1(n275), .B2(n120), .ZN(n130) );
  OAI21_X1 U122 ( .B1(n260), .B2(n124), .A(n131), .ZN(n88) );
  AOI22_X1 U123 ( .A1(n126), .A2(n123), .B1(n275), .B2(n122), .ZN(n131) );
  NAND2_X1 U124 ( .A1(n132), .A2(n133), .ZN(B[1]) );
  NOR3_X1 U125 ( .A1(n134), .A2(n135), .A3(n136), .ZN(n133) );
  NAND2_X1 U126 ( .A1(n137), .A2(n138), .ZN(n49) );
  AOI22_X1 U127 ( .A1(A[12]), .A2(n241), .B1(A[11]), .B2(n98), .ZN(n138) );
  AOI22_X1 U128 ( .A1(A[10]), .A2(n99), .B1(A[9]), .B2(n100), .ZN(n137) );
  AOI21_X1 U129 ( .B1(n139), .B2(n140), .A(n96), .ZN(n135) );
  AOI22_X1 U130 ( .A1(A[4]), .A2(n97), .B1(A[3]), .B2(n98), .ZN(n140) );
  AOI22_X1 U131 ( .A1(A[2]), .A2(n99), .B1(A[1]), .B2(n100), .ZN(n139) );
  NOR2_X1 U132 ( .A1(n262), .A2(n55), .ZN(n134) );
  AOI22_X1 U133 ( .A1(n237), .A2(n81), .B1(SH[4]), .B2(n141), .ZN(n132) );
  NAND2_X1 U134 ( .A1(n142), .A2(n143), .ZN(n81) );
  AOI22_X1 U135 ( .A1(A[8]), .A2(n97), .B1(A[7]), .B2(n98), .ZN(n143) );
  AOI22_X1 U136 ( .A1(A[6]), .A2(n99), .B1(A[5]), .B2(n100), .ZN(n142) );
  OAI21_X1 U137 ( .B1(n249), .B2(n243), .A(n144), .ZN(n101) );
  AOI22_X1 U138 ( .A1(n275), .A2(n145), .B1(n274), .B2(n66), .ZN(n144) );
  NAND2_X1 U139 ( .A1(n147), .A2(n148), .ZN(n113) );
  AOI22_X1 U140 ( .A1(n149), .A2(n266), .B1(n126), .B2(n129), .ZN(n148) );
  AOI22_X1 U141 ( .A1(n275), .A2(n150), .B1(n274), .B2(n151), .ZN(n147) );
  NAND2_X1 U142 ( .A1(n152), .A2(n153), .ZN(n141) );
  AOI22_X1 U143 ( .A1(n149), .A2(n267), .B1(n126), .B2(n120), .ZN(n153) );
  AOI22_X1 U144 ( .A1(n275), .A2(n47), .B1(n274), .B2(n48), .ZN(n152) );
  NAND2_X1 U145 ( .A1(n155), .A2(n156), .ZN(B[15]) );
  AOI21_X1 U146 ( .B1(n270), .B2(n127), .A(n157), .ZN(n156) );
  OAI21_X1 U147 ( .B1(n251), .B2(n45), .A(n158), .ZN(n157) );
  NAND2_X1 U148 ( .A1(n272), .A2(n269), .ZN(n158) );
  AOI22_X1 U149 ( .A1(n42), .A2(n66), .B1(n273), .B2(n65), .ZN(n155) );
  NAND2_X1 U150 ( .A1(n159), .A2(n160), .ZN(B[14]) );
  AOI21_X1 U151 ( .B1(n270), .B2(n129), .A(n161), .ZN(n160) );
  OAI21_X1 U152 ( .B1(n253), .B2(n45), .A(n162), .ZN(n161) );
  NAND2_X1 U153 ( .A1(n272), .A2(n266), .ZN(n162) );
  AOI22_X1 U154 ( .A1(n237), .A2(n151), .B1(n273), .B2(n74), .ZN(n159) );
  NAND2_X1 U155 ( .A1(n163), .A2(n164), .ZN(B[13]) );
  AOI21_X1 U156 ( .B1(n270), .B2(n120), .A(n165), .ZN(n164) );
  OAI21_X1 U157 ( .B1(n116), .B2(n166), .A(n167), .ZN(n165) );
  NAND2_X1 U158 ( .A1(n271), .A2(n47), .ZN(n167) );
  NAND2_X1 U159 ( .A1(n168), .A2(n169), .ZN(n47) );
  AOI22_X1 U160 ( .A1(A[24]), .A2(n97), .B1(A[23]), .B2(n98), .ZN(n169) );
  AOI22_X1 U161 ( .A1(A[22]), .A2(n99), .B1(A[21]), .B2(n100), .ZN(n168) );
  AOI21_X1 U162 ( .B1(n238), .B2(A[29]), .A(n268), .ZN(n116) );
  AOI22_X1 U163 ( .A1(A[31]), .A2(n240), .B1(A[30]), .B2(n239), .ZN(n170) );
  NAND2_X1 U164 ( .A1(n171), .A2(n172), .ZN(n120) );
  AOI22_X1 U165 ( .A1(A[28]), .A2(n97), .B1(A[27]), .B2(n98), .ZN(n172) );
  AOI22_X1 U166 ( .A1(A[26]), .A2(n99), .B1(A[25]), .B2(n100), .ZN(n171) );
  AOI22_X1 U167 ( .A1(n42), .A2(n48), .B1(n273), .B2(n43), .ZN(n163) );
  NAND2_X1 U168 ( .A1(n173), .A2(n174), .ZN(n43) );
  AOI22_X1 U169 ( .A1(A[16]), .A2(n97), .B1(A[15]), .B2(n98), .ZN(n174) );
  AOI22_X1 U170 ( .A1(A[14]), .A2(n99), .B1(A[13]), .B2(n238), .ZN(n173) );
  NAND2_X1 U171 ( .A1(n175), .A2(n176), .ZN(n48) );
  AOI22_X1 U172 ( .A1(A[20]), .A2(n97), .B1(A[19]), .B2(n98), .ZN(n176) );
  AOI22_X1 U173 ( .A1(A[18]), .A2(n239), .B1(A[17]), .B2(n238), .ZN(n175) );
  NAND2_X1 U174 ( .A1(n177), .A2(n178), .ZN(B[12]) );
  AOI21_X1 U175 ( .B1(n270), .B2(n122), .A(n179), .ZN(n178) );
  OAI21_X1 U176 ( .B1(n260), .B2(n45), .A(n180), .ZN(n179) );
  NAND2_X1 U177 ( .A1(n272), .A2(n123), .ZN(n180) );
  NAND2_X1 U178 ( .A1(SH[4]), .A2(n274), .ZN(n166) );
  AOI22_X1 U179 ( .A1(n42), .A2(n57), .B1(n273), .B2(n53), .ZN(n177) );
  NAND2_X1 U180 ( .A1(n182), .A2(n183), .ZN(B[11]) );
  AOI21_X1 U181 ( .B1(n270), .B2(n145), .A(n184), .ZN(n183) );
  OAI21_X1 U182 ( .B1(n242), .B2(n185), .A(n186), .ZN(n184) );
  NAND2_X1 U183 ( .A1(n271), .A2(n66), .ZN(n186) );
  NAND2_X1 U184 ( .A1(n187), .A2(n188), .ZN(n66) );
  AOI22_X1 U185 ( .A1(A[22]), .A2(n241), .B1(A[21]), .B2(n240), .ZN(n188) );
  AOI22_X1 U186 ( .A1(n239), .A2(A[20]), .B1(n100), .B2(A[19]), .ZN(n187) );
  NAND2_X1 U187 ( .A1(n146), .A2(n243), .ZN(n185) );
  MUX2_X2 U188 ( .A(n127), .B(n269), .S(SH[2]), .Z(n146) );
  NAND2_X1 U189 ( .A1(A[31]), .A2(n238), .ZN(n104) );
  NAND2_X1 U190 ( .A1(n189), .A2(n190), .ZN(n127) );
  AOI22_X1 U191 ( .A1(A[30]), .A2(n241), .B1(A[29]), .B2(n240), .ZN(n190) );
  AOI22_X1 U192 ( .A1(A[28]), .A2(n99), .B1(A[27]), .B2(n238), .ZN(n189) );
  NAND2_X1 U193 ( .A1(n191), .A2(n192), .ZN(n145) );
  AOI22_X1 U194 ( .A1(A[26]), .A2(n241), .B1(A[25]), .B2(n240), .ZN(n192) );
  AOI22_X1 U195 ( .A1(A[24]), .A2(n239), .B1(A[23]), .B2(n238), .ZN(n191) );
  AOI22_X1 U196 ( .A1(n237), .A2(n65), .B1(n273), .B2(n62), .ZN(n182) );
  NAND2_X1 U197 ( .A1(n193), .A2(n194), .ZN(n62) );
  AOI22_X1 U198 ( .A1(A[14]), .A2(n241), .B1(A[13]), .B2(n240), .ZN(n194) );
  AOI22_X1 U199 ( .A1(A[12]), .A2(n99), .B1(A[11]), .B2(n238), .ZN(n193) );
  NAND2_X1 U200 ( .A1(n195), .A2(n196), .ZN(n65) );
  AOI22_X1 U201 ( .A1(A[18]), .A2(n241), .B1(A[17]), .B2(n240), .ZN(n196) );
  AOI22_X1 U202 ( .A1(A[16]), .A2(n99), .B1(A[15]), .B2(n238), .ZN(n195) );
  NAND2_X1 U203 ( .A1(n197), .A2(n198), .ZN(B[10]) );
  AOI21_X1 U204 ( .B1(n237), .B2(n74), .A(n199), .ZN(n198) );
  OAI21_X1 U205 ( .B1(n254), .B2(n45), .A(n200), .ZN(n199) );
  NAND2_X1 U206 ( .A1(n270), .A2(n150), .ZN(n200) );
  NAND2_X1 U207 ( .A1(n201), .A2(n202), .ZN(n150) );
  AOI22_X1 U208 ( .A1(A[25]), .A2(n241), .B1(A[24]), .B2(n240), .ZN(n202) );
  AOI22_X1 U209 ( .A1(A[23]), .A2(n99), .B1(A[22]), .B2(n238), .ZN(n201) );
  NAND2_X1 U210 ( .A1(n203), .A2(n204), .ZN(n151) );
  AOI22_X1 U211 ( .A1(A[21]), .A2(n241), .B1(n98), .B2(A[20]), .ZN(n204) );
  AOI22_X1 U212 ( .A1(n239), .A2(A[19]), .B1(n100), .B2(A[18]), .ZN(n203) );
  NAND2_X1 U213 ( .A1(n205), .A2(n206), .ZN(n74) );
  AOI22_X1 U214 ( .A1(A[17]), .A2(n241), .B1(A[16]), .B2(n240), .ZN(n206) );
  AOI22_X1 U215 ( .A1(A[15]), .A2(n239), .B1(A[14]), .B2(n238), .ZN(n205) );
  AOI22_X1 U216 ( .A1(n273), .A2(n71), .B1(SH[4]), .B2(n255), .ZN(n197) );
  AOI21_X1 U217 ( .B1(n129), .B2(n274), .A(n207), .ZN(n117) );
  NOR2_X1 U218 ( .A1(n118), .A2(n105), .ZN(n207) );
  AOI21_X1 U219 ( .B1(n239), .B2(A[31]), .A(n208), .ZN(n105) );
  AND2_X2 U220 ( .A1(A[30]), .A2(n238), .ZN(n208) );
  NAND2_X1 U221 ( .A1(n209), .A2(n210), .ZN(n129) );
  AOI22_X1 U222 ( .A1(A[29]), .A2(n241), .B1(A[28]), .B2(n240), .ZN(n210) );
  AOI22_X1 U223 ( .A1(A[27]), .A2(n99), .B1(A[26]), .B2(n238), .ZN(n209) );
  NAND2_X1 U224 ( .A1(n211), .A2(n212), .ZN(n71) );
  AOI22_X1 U225 ( .A1(A[13]), .A2(n241), .B1(A[12]), .B2(n240), .ZN(n212) );
  AOI22_X1 U226 ( .A1(A[11]), .A2(n239), .B1(A[10]), .B2(n238), .ZN(n211) );
  NAND2_X1 U227 ( .A1(n213), .A2(n214), .ZN(B[0]) );
  NOR3_X1 U228 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n214) );
  NAND2_X1 U229 ( .A1(n218), .A2(n244), .ZN(n45) );
  NAND2_X1 U230 ( .A1(n219), .A2(n220), .ZN(n58) );
  AOI22_X1 U231 ( .A1(A[11]), .A2(n241), .B1(A[10]), .B2(n240), .ZN(n220) );
  AOI22_X1 U232 ( .A1(A[9]), .A2(n239), .B1(A[8]), .B2(n238), .ZN(n219) );
  AOI21_X1 U233 ( .B1(n221), .B2(n222), .A(n96), .ZN(n216) );
  NAND2_X1 U234 ( .A1(n274), .A2(n242), .ZN(n96) );
  AOI22_X1 U235 ( .A1(A[3]), .A2(n241), .B1(A[2]), .B2(n240), .ZN(n222) );
  AOI22_X1 U236 ( .A1(A[1]), .A2(n239), .B1(A[0]), .B2(n238), .ZN(n221) );
  NOR2_X1 U237 ( .A1(n256), .A2(n55), .ZN(n215) );
  NAND2_X1 U238 ( .A1(SH[2]), .A2(n218), .ZN(n55) );
  NOR2_X1 U239 ( .A1(n243), .A2(SH[4]), .ZN(n218) );
  NAND2_X1 U240 ( .A1(n223), .A2(n224), .ZN(n53) );
  AOI22_X1 U241 ( .A1(A[15]), .A2(n97), .B1(A[14]), .B2(n240), .ZN(n224) );
  AOI22_X1 U242 ( .A1(A[13]), .A2(n239), .B1(A[12]), .B2(n238), .ZN(n223) );
  AOI22_X1 U243 ( .A1(n42), .A2(n87), .B1(SH[4]), .B2(n154), .ZN(n213) );
  NAND2_X1 U244 ( .A1(n225), .A2(n226), .ZN(n154) );
  AOI22_X1 U245 ( .A1(n149), .A2(n123), .B1(n126), .B2(n122), .ZN(n226) );
  NAND2_X1 U246 ( .A1(n227), .A2(n228), .ZN(n122) );
  AOI22_X1 U247 ( .A1(A[27]), .A2(n241), .B1(A[26]), .B2(n240), .ZN(n228) );
  AOI22_X1 U248 ( .A1(A[25]), .A2(n239), .B1(A[24]), .B2(n238), .ZN(n227) );
  NOR2_X1 U249 ( .A1(n243), .A2(SH[2]), .ZN(n126) );
  NAND2_X1 U250 ( .A1(n229), .A2(n230), .ZN(n123) );
  AOI22_X1 U251 ( .A1(A[31]), .A2(n97), .B1(A[30]), .B2(n240), .ZN(n230) );
  AOI22_X1 U252 ( .A1(A[29]), .A2(n239), .B1(A[28]), .B2(n238), .ZN(n229) );
  NOR2_X1 U253 ( .A1(n244), .A2(n243), .ZN(n149) );
  AOI22_X1 U254 ( .A1(n275), .A2(n181), .B1(n274), .B2(n57), .ZN(n225) );
  NAND2_X1 U255 ( .A1(n231), .A2(n232), .ZN(n57) );
  AOI22_X1 U256 ( .A1(A[19]), .A2(n97), .B1(A[18]), .B2(n240), .ZN(n232) );
  AOI22_X1 U257 ( .A1(A[17]), .A2(n239), .B1(A[16]), .B2(n238), .ZN(n231) );
  NAND2_X1 U258 ( .A1(n244), .A2(n243), .ZN(n124) );
  NAND2_X1 U259 ( .A1(n233), .A2(n234), .ZN(n181) );
  AOI22_X1 U260 ( .A1(A[23]), .A2(n97), .B1(A[22]), .B2(n240), .ZN(n234) );
  AOI22_X1 U261 ( .A1(A[21]), .A2(n239), .B1(n100), .B2(A[20]), .ZN(n233) );
  NAND2_X1 U262 ( .A1(n235), .A2(n236), .ZN(n87) );
  AOI22_X1 U263 ( .A1(A[7]), .A2(n97), .B1(A[6]), .B2(n240), .ZN(n236) );
  NOR2_X1 U264 ( .A1(n245), .A2(SH[0]), .ZN(n98) );
  NOR2_X1 U265 ( .A1(n245), .A2(n246), .ZN(n97) );
  AOI22_X1 U266 ( .A1(A[5]), .A2(n239), .B1(A[4]), .B2(n238), .ZN(n235) );
  NOR2_X1 U267 ( .A1(SH[0]), .A2(SH[1]), .ZN(n100) );
  NOR2_X1 U268 ( .A1(n246), .A2(SH[1]), .ZN(n99) );
  NOR2_X1 U269 ( .A1(n118), .A2(SH[4]), .ZN(n42) );
  NAND2_X1 U270 ( .A1(SH[2]), .A2(n243), .ZN(n118) );
  AOI21_X1 U8 ( .B1(n205), .B2(n206), .A(n55), .ZN(n108) );
  AOI21_X1 U10 ( .B1(n195), .B2(n196), .A(n55), .ZN(n91) );
  INV_X1 U12 ( .A(n55), .ZN(n270) );
  CLKBUF_X1 U14 ( .A(n42), .Z(n237) );
  INV_X1 U19 ( .A(n166), .ZN(n272) );
  INV_X1 U21 ( .A(n96), .ZN(n273) );
  INV_X1 U23 ( .A(n117), .ZN(n255) );
  INV_X1 U24 ( .A(n124), .ZN(n274) );
  INV_X1 U25 ( .A(n118), .ZN(n275) );
  CLKBUF_X1 U26 ( .A(n97), .Z(n241) );
  INV_X1 U27 ( .A(n45), .ZN(n271) );
  INV_X1 U28 ( .A(n146), .ZN(n249) );
  INV_X1 U29 ( .A(n47), .ZN(n265) );
  INV_X1 U30 ( .A(n48), .ZN(n261) );
  CLKBUF_X1 U31 ( .A(n100), .Z(n238) );
  CLKBUF_X1 U32 ( .A(n98), .Z(n240) );
  INV_X1 U33 ( .A(n66), .ZN(n247) );
  INV_X1 U34 ( .A(n5), .ZN(B[19]) );
  INV_X1 U35 ( .A(n2), .ZN(B[21]) );
  INV_X1 U36 ( .A(n3), .ZN(B[22]) );
  INV_X1 U37 ( .A(n4), .ZN(B[23]) );
  INV_X1 U38 ( .A(n7), .ZN(B[25]) );
  CLKBUF_X1 U39 ( .A(n99), .Z(n239) );
  INV_X1 U40 ( .A(n116), .ZN(n267) );
  INV_X1 U41 ( .A(n105), .ZN(n266) );
  INV_X1 U42 ( .A(n104), .ZN(n269) );
  INV_X1 U43 ( .A(n181), .ZN(n260) );
  INV_X1 U44 ( .A(n123), .ZN(n259) );
  INV_X1 U45 ( .A(n43), .ZN(n262) );
  INV_X1 U46 ( .A(n53), .ZN(n256) );
  INV_X1 U47 ( .A(n145), .ZN(n251) );
  INV_X1 U48 ( .A(n150), .ZN(n253) );
  INV_X1 U49 ( .A(n151), .ZN(n254) );
  INV_X1 U50 ( .A(n6), .ZN(B[24]) );
  INV_X1 U51 ( .A(n1), .ZN(B[20]) );
  INV_X1 U52 ( .A(n170), .ZN(n268) );
  INV_X1 U53 ( .A(SH[2]), .ZN(n244) );
  INV_X1 U54 ( .A(SH[4]), .ZN(n242) );
  INV_X1 U55 ( .A(SH[3]), .ZN(n243) );
  INV_X1 U91 ( .A(SH[1]), .ZN(n245) );
  INV_X1 U103 ( .A(SH[0]), .ZN(n246) );
endmodule



    module DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW01_ash_0 ( 
        A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[3][31] , \ML_int[3][30] ,
         \ML_int[3][29] , \ML_int[3][28] , \ML_int[3][27] , \ML_int[3][26] ,
         \ML_int[3][25] , \ML_int[3][24] , \ML_int[3][23] , \ML_int[3][22] ,
         \ML_int[3][21] , \ML_int[3][20] , \ML_int[3][19] , \ML_int[3][18] ,
         \ML_int[3][17] , \ML_int[3][16] , \ML_int[3][15] , \ML_int[3][14] ,
         \ML_int[3][13] , \ML_int[3][12] , \ML_int[3][11] , \ML_int[3][10] ,
         \ML_int[3][9] , \ML_int[3][8] , \ML_int[3][7] , \ML_int[3][6] ,
         \ML_int[3][5] , \ML_int[3][4] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[5][31] , \ML_int[5][30] , \ML_int[5][29] , \ML_int[5][28] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] , \ML_int[5][16] ,
         \ML_int[5][7] , \ML_int[5][6] , \ML_int[5][5] , \ML_int[5][4] ,
         \ML_int[5][3] , \ML_int[5][2] , \ML_int[5][1] , \ML_int[5][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n49,
         n50, n53, n54, n55, n61, n62, n63, n64, n65, n66;
  assign B[31] = \ML_int[5][31] ;
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;
  assign B[22] = \ML_int[5][22] ;
  assign B[21] = \ML_int[5][21] ;
  assign B[20] = \ML_int[5][20] ;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[7] = \ML_int[5][7] ;
  assign B[6] = \ML_int[5][6] ;
  assign B[5] = \ML_int[5][5] ;
  assign B[4] = \ML_int[5][4] ;
  assign B[3] = \ML_int[5][3] ;
  assign B[2] = \ML_int[5][2] ;
  assign B[1] = \ML_int[5][1] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2_X2 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n39), .Z(
        \ML_int[5][31] ) );
  MUX2_X2 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n39), .Z(
        \ML_int[5][30] ) );
  MUX2_X2 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n39), .Z(
        \ML_int[5][29] ) );
  MUX2_X2 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n39), .Z(
        \ML_int[5][28] ) );
  MUX2_X2 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n39), .Z(
        \ML_int[5][27] ) );
  MUX2_X2 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n39), .Z(
        \ML_int[5][26] ) );
  MUX2_X2 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n39), .Z(
        \ML_int[5][25] ) );
  MUX2_X2 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n39), .Z(
        \ML_int[5][24] ) );
  MUX2_X2 M1_4_23 ( .A(\ML_int[4][23] ), .B(n61), .S(n39), .Z(\ML_int[5][23] )
         );
  MUX2_X2 M1_4_22 ( .A(\ML_int[4][22] ), .B(n55), .S(n39), .Z(\ML_int[5][22] )
         );
  MUX2_X2 M1_4_21 ( .A(\ML_int[4][21] ), .B(n62), .S(n39), .Z(\ML_int[5][21] )
         );
  MUX2_X2 M1_4_20 ( .A(\ML_int[4][20] ), .B(n47), .S(n39), .Z(\ML_int[5][20] )
         );
  MUX2_X2 M1_4_19 ( .A(\ML_int[4][19] ), .B(n63), .S(n39), .Z(\ML_int[5][19] )
         );
  MUX2_X2 M1_4_18 ( .A(\ML_int[4][18] ), .B(n53), .S(n39), .Z(\ML_int[5][18] )
         );
  MUX2_X2 M1_4_17 ( .A(\ML_int[4][17] ), .B(n66), .S(n39), .Z(\ML_int[5][17] )
         );
  MUX2_X2 M1_4_16 ( .A(\ML_int[4][16] ), .B(n50), .S(n39), .Z(\ML_int[5][16] )
         );
  MUX2_X2 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(SH[3]), .Z(
        \ML_int[4][31] ) );
  MUX2_X2 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(SH[3]), .Z(
        \ML_int[4][30] ) );
  MUX2_X2 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(SH[3]), .Z(
        \ML_int[4][29] ) );
  MUX2_X2 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(SH[3]), .Z(
        \ML_int[4][28] ) );
  MUX2_X2 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(SH[3]), .Z(
        \ML_int[4][27] ) );
  MUX2_X2 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(SH[3]), .Z(
        \ML_int[4][26] ) );
  MUX2_X2 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(SH[3]), .Z(
        \ML_int[4][25] ) );
  MUX2_X2 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(SH[3]), .Z(
        \ML_int[4][24] ) );
  MUX2_X2 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(SH[3]), .Z(
        \ML_int[4][23] ) );
  MUX2_X2 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(SH[3]), .Z(
        \ML_int[4][22] ) );
  MUX2_X2 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(SH[3]), .Z(
        \ML_int[4][21] ) );
  MUX2_X2 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(SH[3]), .Z(
        \ML_int[4][20] ) );
  MUX2_X2 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2_X2 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2_X2 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2_X2 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(SH[3]), .Z(
        \ML_int[4][16] ) );
  MUX2_X2 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(SH[3]), .Z(
        \ML_int[4][15] ) );
  MUX2_X2 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(SH[3]), .Z(
        \ML_int[4][14] ) );
  MUX2_X2 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(SH[3]), .Z(
        \ML_int[4][13] ) );
  MUX2_X2 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(SH[3]), .Z(
        \ML_int[4][12] ) );
  MUX2_X2 M1_3_11 ( .A(\ML_int[3][11] ), .B(n64), .S(SH[3]), .Z(
        \ML_int[4][11] ) );
  MUX2_X2 M1_3_10 ( .A(\ML_int[3][10] ), .B(n54), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2_X2 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2_X2 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2_X2 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n42), .Z(
        \ML_int[3][31] ) );
  MUX2_X2 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(SH[2]), .Z(
        \ML_int[3][30] ) );
  MUX2_X2 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(SH[2]), .Z(
        \ML_int[3][29] ) );
  MUX2_X2 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n42), .Z(
        \ML_int[3][28] ) );
  MUX2_X2 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n42), .Z(
        \ML_int[3][27] ) );
  MUX2_X2 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(SH[2]), .Z(
        \ML_int[3][26] ) );
  MUX2_X2 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(SH[2]), .Z(
        \ML_int[3][25] ) );
  MUX2_X2 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n42), .Z(
        \ML_int[3][24] ) );
  MUX2_X2 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(SH[2]), .Z(
        \ML_int[3][23] ) );
  MUX2_X2 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(SH[2]), .Z(
        \ML_int[3][22] ) );
  MUX2_X2 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(SH[2]), .Z(
        \ML_int[3][21] ) );
  MUX2_X2 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n42), .Z(
        \ML_int[3][20] ) );
  MUX2_X2 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2_X2 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n42), .Z(
        \ML_int[3][18] ) );
  MUX2_X2 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n42), .Z(
        \ML_int[3][17] ) );
  MUX2_X2 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n42), .Z(
        \ML_int[3][16] ) );
  MUX2_X2 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n42), .Z(
        \ML_int[3][15] ) );
  MUX2_X2 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n42), .Z(
        \ML_int[3][14] ) );
  MUX2_X2 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n42), .Z(
        \ML_int[3][13] ) );
  MUX2_X2 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n42), .Z(
        \ML_int[3][12] ) );
  MUX2_X2 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n42), .Z(
        \ML_int[3][11] ) );
  MUX2_X2 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n42), .Z(
        \ML_int[3][10] ) );
  MUX2_X2 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n42), .Z(
        \ML_int[3][9] ) );
  MUX2_X2 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2_X2 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2_X2 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n42), .Z(
        \ML_int[3][6] ) );
  MUX2_X2 M1_2_5 ( .A(\ML_int[2][5] ), .B(n65), .S(SH[2]), .Z(\ML_int[3][5] )
         );
  MUX2_X2 M1_2_4 ( .A(\ML_int[2][4] ), .B(n49), .S(n42), .Z(\ML_int[3][4] ) );
  MUX2_X2 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(SH[1]), .Z(
        \ML_int[2][31] ) );
  MUX2_X2 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(SH[1]), .Z(
        \ML_int[2][30] ) );
  MUX2_X2 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(SH[1]), .Z(
        \ML_int[2][29] ) );
  MUX2_X2 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(SH[1]), .Z(
        \ML_int[2][28] ) );
  MUX2_X2 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(SH[1]), .Z(
        \ML_int[2][27] ) );
  MUX2_X2 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(SH[1]), .Z(
        \ML_int[2][26] ) );
  MUX2_X2 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(SH[1]), .Z(
        \ML_int[2][25] ) );
  MUX2_X2 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(SH[1]), .Z(
        \ML_int[2][24] ) );
  MUX2_X2 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(SH[1]), .Z(
        \ML_int[2][23] ) );
  MUX2_X2 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(SH[1]), .Z(
        \ML_int[2][22] ) );
  MUX2_X2 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(SH[1]), .Z(
        \ML_int[2][21] ) );
  MUX2_X2 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(SH[1]), .Z(
        \ML_int[2][20] ) );
  MUX2_X2 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2_X2 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2_X2 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2_X2 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2_X2 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2_X2 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2_X2 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2_X2 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2_X2 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2_X2 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2_X2 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2_X2 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2_X2 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2_X2 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2_X2 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2_X2 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2_X2 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2_X2 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2_X2 M1_0_31 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Z(\ML_int[1][31] ) );
  MUX2_X2 M1_0_30 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Z(\ML_int[1][30] ) );
  MUX2_X2 M1_0_29 ( .A(A[29]), .B(A[28]), .S(SH[0]), .Z(\ML_int[1][29] ) );
  MUX2_X2 M1_0_28 ( .A(A[28]), .B(A[27]), .S(SH[0]), .Z(\ML_int[1][28] ) );
  MUX2_X2 M1_0_27 ( .A(A[27]), .B(A[26]), .S(SH[0]), .Z(\ML_int[1][27] ) );
  MUX2_X2 M1_0_26 ( .A(A[26]), .B(A[25]), .S(SH[0]), .Z(\ML_int[1][26] ) );
  MUX2_X2 M1_0_25 ( .A(A[25]), .B(A[24]), .S(SH[0]), .Z(\ML_int[1][25] ) );
  MUX2_X2 M1_0_24 ( .A(A[24]), .B(A[23]), .S(SH[0]), .Z(\ML_int[1][24] ) );
  MUX2_X2 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n45), .Z(\ML_int[1][23] ) );
  MUX2_X2 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n45), .Z(\ML_int[1][22] ) );
  MUX2_X2 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n45), .Z(\ML_int[1][21] ) );
  MUX2_X2 M1_0_20 ( .A(A[20]), .B(A[19]), .S(SH[0]), .Z(\ML_int[1][20] ) );
  MUX2_X2 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n45), .Z(\ML_int[1][19] ) );
  MUX2_X2 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n45), .Z(\ML_int[1][18] ) );
  MUX2_X2 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n45), .Z(\ML_int[1][17] ) );
  MUX2_X2 M1_0_16 ( .A(A[16]), .B(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2_X2 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n45), .Z(\ML_int[1][15] ) );
  MUX2_X2 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n45), .Z(\ML_int[1][14] ) );
  MUX2_X2 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n45), .Z(\ML_int[1][13] ) );
  MUX2_X2 M1_0_12 ( .A(A[12]), .B(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2_X2 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n45), .Z(\ML_int[1][11] ) );
  MUX2_X2 M1_0_10 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2_X2 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n45), .Z(\ML_int[1][9] ) );
  MUX2_X2 M1_0_8 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2_X2 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n45), .Z(\ML_int[1][7] ) );
  MUX2_X2 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n45), .Z(\ML_int[1][6] ) );
  MUX2_X2 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n45), .Z(\ML_int[1][5] ) );
  MUX2_X2 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n45), .Z(\ML_int[1][4] ) );
  MUX2_X2 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n45), .Z(\ML_int[1][3] ) );
  MUX2_X2 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n45), .Z(\ML_int[1][2] ) );
  MUX2_X2 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n45), .Z(\ML_int[1][1] ) );
  NAND2_X1 U3 ( .A1(\ML_int[4][8] ), .A2(n40), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\ML_int[4][9] ), .A2(n40), .ZN(n2) );
  NAND2_X1 U7 ( .A1(\ML_int[4][10] ), .A2(n40), .ZN(n3) );
  NAND2_X1 U9 ( .A1(\ML_int[4][11] ), .A2(n40), .ZN(n4) );
  NAND2_X1 U11 ( .A1(\ML_int[4][13] ), .A2(n40), .ZN(n5) );
  NAND2_X1 U13 ( .A1(\ML_int[4][14] ), .A2(n40), .ZN(n6) );
  NAND2_X1 U15 ( .A1(\ML_int[2][2] ), .A2(n43), .ZN(n7) );
  NAND2_X1 U17 ( .A1(\ML_int[4][15] ), .A2(n40), .ZN(n8) );
  NAND2_X1 U19 ( .A1(\ML_int[2][3] ), .A2(n43), .ZN(n9) );
  NAND2_X1 U21 ( .A1(\ML_int[4][12] ), .A2(n40), .ZN(n10) );
  NOR2_X1 U41 ( .A1(SH[4]), .A2(n29), .ZN(\ML_int[5][7] ) );
  NOR2_X1 U42 ( .A1(SH[4]), .A2(n30), .ZN(\ML_int[5][6] ) );
  NOR2_X1 U43 ( .A1(SH[4]), .A2(n31), .ZN(\ML_int[5][5] ) );
  NOR2_X1 U44 ( .A1(n39), .A2(n32), .ZN(\ML_int[5][4] ) );
  NOR2_X1 U45 ( .A1(n39), .A2(n33), .ZN(\ML_int[5][3] ) );
  NOR2_X1 U46 ( .A1(SH[4]), .A2(n34), .ZN(\ML_int[5][2] ) );
  NOR2_X1 U47 ( .A1(SH[4]), .A2(n35), .ZN(\ML_int[5][1] ) );
  NOR2_X1 U48 ( .A1(n39), .A2(n36), .ZN(\ML_int[5][0] ) );
  NAND2_X1 U49 ( .A1(\ML_int[3][7] ), .A2(n41), .ZN(n29) );
  NAND2_X1 U50 ( .A1(\ML_int[3][6] ), .A2(n41), .ZN(n30) );
  NAND2_X1 U51 ( .A1(\ML_int[3][5] ), .A2(n41), .ZN(n31) );
  NAND2_X1 U52 ( .A1(\ML_int[3][4] ), .A2(n41), .ZN(n32) );
  NAND2_X1 U53 ( .A1(n64), .A2(n41), .ZN(n33) );
  NAND2_X1 U54 ( .A1(n54), .A2(n41), .ZN(n34) );
  NAND2_X1 U55 ( .A1(\ML_int[3][1] ), .A2(n41), .ZN(n35) );
  NAND2_X1 U56 ( .A1(\ML_int[3][0] ), .A2(n41), .ZN(n36) );
  NOR2_X1 U57 ( .A1(n37), .A2(n42), .ZN(\ML_int[3][1] ) );
  NOR2_X1 U58 ( .A1(n38), .A2(SH[2]), .ZN(\ML_int[3][0] ) );
  NAND2_X1 U59 ( .A1(\ML_int[1][1] ), .A2(n44), .ZN(n37) );
  NAND2_X1 U60 ( .A1(\ML_int[1][0] ), .A2(n44), .ZN(n38) );
  AND2_X2 U61 ( .A1(A[0]), .A2(n46), .ZN(\ML_int[1][0] ) );
  INV_X1 U4 ( .A(n31), .ZN(n62) );
  INV_X1 U6 ( .A(n30), .ZN(n55) );
  INV_X1 U8 ( .A(n29), .ZN(n61) );
  INV_X1 U10 ( .A(n34), .ZN(n53) );
  INV_X1 U12 ( .A(n33), .ZN(n63) );
  INV_X1 U14 ( .A(n35), .ZN(n66) );
  INV_X1 U16 ( .A(n37), .ZN(n65) );
  INV_X1 U18 ( .A(n38), .ZN(n49) );
  INV_X1 U20 ( .A(n46), .ZN(n45) );
  INV_X1 U22 ( .A(n43), .ZN(n42) );
  INV_X1 U23 ( .A(n40), .ZN(n39) );
  INV_X1 U24 ( .A(n32), .ZN(n47) );
  INV_X1 U25 ( .A(n36), .ZN(n50) );
  INV_X1 U26 ( .A(n1), .ZN(B[8]) );
  INV_X1 U27 ( .A(n10), .ZN(B[12]) );
  INV_X1 U28 ( .A(n2), .ZN(B[9]) );
  INV_X1 U29 ( .A(n3), .ZN(B[10]) );
  INV_X1 U30 ( .A(n4), .ZN(B[11]) );
  INV_X1 U31 ( .A(n5), .ZN(B[13]) );
  INV_X1 U32 ( .A(n6), .ZN(B[14]) );
  INV_X1 U33 ( .A(n8), .ZN(B[15]) );
  INV_X1 U34 ( .A(n7), .ZN(n54) );
  INV_X1 U35 ( .A(n9), .ZN(n64) );
  INV_X1 U36 ( .A(SH[4]), .ZN(n40) );
  INV_X1 U37 ( .A(SH[3]), .ZN(n41) );
  INV_X1 U38 ( .A(SH[1]), .ZN(n44) );
  INV_X1 U39 ( .A(SH[2]), .ZN(n43) );
  INV_X1 U40 ( .A(SH[0]), .ZN(n46) );
endmodule



    module DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW01_inc_0 ( 
        A, SUM );
  input [17:0] A;
  output [17:0] SUM;

  wire   [17:2] carry;
  assign carry[2] = A[1];

  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2_X1 U2 ( .A(carry[17]), .B(A[17]), .Z(SUM[17]) );
  INV_X1 U1 ( .A(carry[2]), .ZN(SUM[1]) );
endmodule



    module DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW01_inc_1 ( 
        A, SUM );
  input [17:0] A;
  output [17:0] SUM;

  wire   [17:2] carry;

  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U2 ( .A(carry[17]), .B(A[17]), .Z(SUM[17]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
endmodule



    module DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4 ( 
        Clk, Rst, PC_out, IR_in, DataAddr, DataOut, DataIn_w, DataIn_hw, 
        DataIn_b, DRAM_WE, DRAM_RE, DRAMOP_SEL, SPILL, FILL, stackBus_In, 
        stackBus_Out );
  output [31:0] PC_out;
  input [31:0] IR_in;
  output [31:0] DataAddr;
  output [31:0] DataOut;
  input [31:0] DataIn_w;
  input [15:0] DataIn_hw;
  input [7:0] DataIn_b;
  input [127:0] stackBus_In;
  output [127:0] stackBus_Out;
  input Clk, Rst;
  output DRAM_WE, DRAM_RE, DRAMOP_SEL, SPILL, FILL;
  wire   n74605, \DLX_Datapath/N358 , \DLX_Datapath/N357 , \DLX_Datapath/N356 ,
         \DLX_Datapath/N355 , \DLX_Datapath/N354 , \DLX_Datapath/N353 ,
         \DLX_Datapath/N352 , \DLX_Datapath/N351 , \DLX_Datapath/N350 ,
         \DLX_Datapath/N349 , \DLX_Datapath/N348 , \DLX_Datapath/N347 ,
         \DLX_Datapath/N346 , \DLX_Datapath/N345 , \DLX_Datapath/N344 ,
         \DLX_Datapath/N343 , \DLX_Datapath/next_A_IDEX[0] ,
         \DLX_Datapath/next_A_IDEX[1] , \DLX_Datapath/next_A_IDEX[2] ,
         \DLX_Datapath/next_A_IDEX[3] , \DLX_Datapath/next_A_IDEX[4] ,
         \DLX_Datapath/next_A_IDEX[5] , \DLX_Datapath/next_A_IDEX[6] ,
         \DLX_Datapath/next_A_IDEX[7] , \DLX_Datapath/next_A_IDEX[8] ,
         \DLX_Datapath/next_A_IDEX[9] , \DLX_Datapath/next_A_IDEX[10] ,
         \DLX_Datapath/next_A_IDEX[11] , \DLX_Datapath/next_A_IDEX[12] ,
         \DLX_Datapath/next_A_IDEX[13] , \DLX_Datapath/next_A_IDEX[14] ,
         \DLX_Datapath/next_A_IDEX[15] , \DLX_Datapath/next_A_IDEX[16] ,
         \DLX_Datapath/next_A_IDEX[17] , \DLX_Datapath/next_A_IDEX[18] ,
         \DLX_Datapath/next_A_IDEX[19] , \DLX_Datapath/next_A_IDEX[20] ,
         \DLX_Datapath/next_A_IDEX[21] , \DLX_Datapath/next_A_IDEX[22] ,
         \DLX_Datapath/next_A_IDEX[23] , \DLX_Datapath/next_A_IDEX[24] ,
         \DLX_Datapath/next_A_IDEX[25] , \DLX_Datapath/next_A_IDEX[26] ,
         \DLX_Datapath/next_A_IDEX[27] , \DLX_Datapath/next_A_IDEX[28] ,
         \DLX_Datapath/next_A_IDEX[29] , \DLX_Datapath/next_A_IDEX[30] ,
         \DLX_Datapath/next_A_IDEX[31] , \DLX_Datapath/CWP_IDEX[1] ,
         \DLX_Datapath/CWP_IDEX[2] , \DLX_Datapath/IR_EXMEM[15] ,
         \DLX_Datapath/IR_EXMEM[20] , \DLX_Datapath/IR_EXMEM[27] ,
         \DLX_Datapath/IR_EXMEM[29] , \DLX_Datapath/IR_EXMEM[31] ,
         \DLX_Datapath/IR_IDEX[15] , \DLX_Datapath/IR_IDEX[20] ,
         \DLX_Datapath/IR_IDEX[27] , \DLX_Datapath/IR_IDEX[29] ,
         \DLX_Datapath/IR_IDEX[31] , \DLX_Datapath/IR_IFID[11] ,
         \DLX_Datapath/IR_IFID[12] , \DLX_Datapath/IR_IFID[13] ,
         \DLX_Datapath/HazardDetUnit/N140 , \DLX_Datapath/HazardDetUnit/N139 ,
         \DLX_Datapath/HazardDetUnit/N138 , \DLX_Datapath/HazardDetUnit/N137 ,
         \DLX_Datapath/HazardDetUnit/N126 , \DLX_Datapath/HazardDetUnit/N125 ,
         \DLX_Datapath/HazardDetUnit/N124 , \DLX_Datapath/HazardDetUnit/N123 ,
         \DLX_Datapath/HazardDetUnit/N112 , \DLX_Datapath/HazardDetUnit/N111 ,
         \DLX_Datapath/HazardDetUnit/N110 , \DLX_Datapath/HazardDetUnit/N109 ,
         \DLX_Datapath/HazardDetUnit/N98 , \DLX_Datapath/HazardDetUnit/N97 ,
         \DLX_Datapath/HazardDetUnit/N96 , \DLX_Datapath/HazardDetUnit/N95 ,
         \DLX_Datapath/RegisterFile/N46899 ,
         \DLX_Datapath/RegisterFile/N46898 ,
         \DLX_Datapath/RegisterFile/N46866 ,
         \DLX_Datapath/RegisterFile/N46424 ,
         \DLX_Datapath/RegisterFile/N46178 ,
         \DLX_Datapath/RegisterFile/N46177 ,
         \DLX_Datapath/RegisterFile/N27074 ,
         \DLX_Datapath/RegisterFile/N26858 ,
         \DLX_Datapath/RegisterFile/N26857 ,
         \DLX_Datapath/RegisterFile/N26856 ,
         \DLX_Datapath/RegisterFile/N26855 ,
         \DLX_Datapath/RegisterFile/N26854 ,
         \DLX_Datapath/RegisterFile/N26853 ,
         \DLX_Datapath/RegisterFile/N26852 ,
         \DLX_Datapath/RegisterFile/N26851 ,
         \DLX_Datapath/RegisterFile/N26850 ,
         \DLX_Datapath/RegisterFile/N26849 ,
         \DLX_Datapath/RegisterFile/N26848 ,
         \DLX_Datapath/RegisterFile/N26847 ,
         \DLX_Datapath/RegisterFile/N26846 ,
         \DLX_Datapath/RegisterFile/N26845 ,
         \DLX_Datapath/RegisterFile/N26844 ,
         \DLX_Datapath/RegisterFile/N26843 ,
         \DLX_Datapath/RegisterFile/N26842 ,
         \DLX_Datapath/RegisterFile/N26841 ,
         \DLX_Datapath/RegisterFile/N26840 ,
         \DLX_Datapath/RegisterFile/N26839 ,
         \DLX_Datapath/RegisterFile/N26838 ,
         \DLX_Datapath/RegisterFile/N26837 ,
         \DLX_Datapath/RegisterFile/N26836 ,
         \DLX_Datapath/RegisterFile/N26835 ,
         \DLX_Datapath/RegisterFile/N26834 ,
         \DLX_Datapath/RegisterFile/N26833 ,
         \DLX_Datapath/RegisterFile/N26832 ,
         \DLX_Datapath/RegisterFile/N26831 ,
         \DLX_Datapath/RegisterFile/N26830 ,
         \DLX_Datapath/RegisterFile/N26829 ,
         \DLX_Datapath/RegisterFile/N26828 ,
         \DLX_Datapath/RegisterFile/N26827 ,
         \DLX_Datapath/RegisterFile/N26826 ,
         \DLX_Datapath/RegisterFile/N26825 ,
         \DLX_Datapath/RegisterFile/N26824 ,
         \DLX_Datapath/RegisterFile/N26823 ,
         \DLX_Datapath/RegisterFile/N26822 ,
         \DLX_Datapath/RegisterFile/N26821 ,
         \DLX_Datapath/RegisterFile/N26820 ,
         \DLX_Datapath/RegisterFile/N26819 ,
         \DLX_Datapath/RegisterFile/N26818 ,
         \DLX_Datapath/RegisterFile/N26817 ,
         \DLX_Datapath/RegisterFile/N26816 ,
         \DLX_Datapath/RegisterFile/N26815 ,
         \DLX_Datapath/RegisterFile/N26814 ,
         \DLX_Datapath/RegisterFile/N26813 ,
         \DLX_Datapath/RegisterFile/N26812 ,
         \DLX_Datapath/RegisterFile/N26811 ,
         \DLX_Datapath/RegisterFile/N26810 ,
         \DLX_Datapath/RegisterFile/N26809 ,
         \DLX_Datapath/RegisterFile/N26808 ,
         \DLX_Datapath/RegisterFile/N26807 ,
         \DLX_Datapath/RegisterFile/N26806 ,
         \DLX_Datapath/RegisterFile/N26805 ,
         \DLX_Datapath/RegisterFile/N26804 ,
         \DLX_Datapath/RegisterFile/N26803 ,
         \DLX_Datapath/RegisterFile/N26802 ,
         \DLX_Datapath/RegisterFile/N26801 ,
         \DLX_Datapath/RegisterFile/N26800 ,
         \DLX_Datapath/RegisterFile/N26799 ,
         \DLX_Datapath/RegisterFile/N26798 ,
         \DLX_Datapath/RegisterFile/N26797 ,
         \DLX_Datapath/RegisterFile/N26796 ,
         \DLX_Datapath/RegisterFile/N26795 ,
         \DLX_Datapath/RegisterFile/N26762 ,
         \DLX_Datapath/RegisterFile/N26761 ,
         \DLX_Datapath/RegisterFile/N26760 ,
         \DLX_Datapath/RegisterFile/N26759 ,
         \DLX_Datapath/RegisterFile/N26758 ,
         \DLX_Datapath/RegisterFile/N26757 ,
         \DLX_Datapath/RegisterFile/N26756 ,
         \DLX_Datapath/RegisterFile/N26755 ,
         \DLX_Datapath/RegisterFile/N26754 ,
         \DLX_Datapath/RegisterFile/N26753 ,
         \DLX_Datapath/RegisterFile/N26752 ,
         \DLX_Datapath/RegisterFile/N26751 ,
         \DLX_Datapath/RegisterFile/N26750 ,
         \DLX_Datapath/RegisterFile/N26749 ,
         \DLX_Datapath/RegisterFile/N26748 ,
         \DLX_Datapath/RegisterFile/N26747 ,
         \DLX_Datapath/RegisterFile/N26746 ,
         \DLX_Datapath/RegisterFile/N26745 ,
         \DLX_Datapath/RegisterFile/N26744 ,
         \DLX_Datapath/RegisterFile/N26743 ,
         \DLX_Datapath/RegisterFile/N26742 ,
         \DLX_Datapath/RegisterFile/N26741 ,
         \DLX_Datapath/RegisterFile/N26739 ,
         \DLX_Datapath/RegisterFile/N26738 ,
         \DLX_Datapath/RegisterFile/N26736 ,
         \DLX_Datapath/RegisterFile/N26735 ,
         \DLX_Datapath/RegisterFile/N26734 ,
         \DLX_Datapath/RegisterFile/N26732 ,
         \DLX_Datapath/RegisterFile/N26731 ,
         \DLX_Datapath/RegisterFile/N26730 ,
         \DLX_Datapath/RegisterFile/N26729 ,
         \DLX_Datapath/RegisterFile/N26728 ,
         \DLX_Datapath/RegisterFile/N26727 ,
         \DLX_Datapath/RegisterFile/N26726 ,
         \DLX_Datapath/RegisterFile/N26725 ,
         \DLX_Datapath/RegisterFile/N26724 ,
         \DLX_Datapath/RegisterFile/N26723 ,
         \DLX_Datapath/RegisterFile/N26722 ,
         \DLX_Datapath/RegisterFile/N26721 ,
         \DLX_Datapath/RegisterFile/N26720 ,
         \DLX_Datapath/RegisterFile/N26719 ,
         \DLX_Datapath/RegisterFile/N26718 ,
         \DLX_Datapath/RegisterFile/N26717 ,
         \DLX_Datapath/RegisterFile/N26716 ,
         \DLX_Datapath/RegisterFile/N26715 ,
         \DLX_Datapath/RegisterFile/N26714 ,
         \DLX_Datapath/RegisterFile/N26713 ,
         \DLX_Datapath/RegisterFile/N26712 ,
         \DLX_Datapath/RegisterFile/N26711 ,
         \DLX_Datapath/RegisterFile/N26710 ,
         \DLX_Datapath/RegisterFile/N26709 ,
         \DLX_Datapath/RegisterFile/N26708 ,
         \DLX_Datapath/RegisterFile/N26707 ,
         \DLX_Datapath/RegisterFile/N26706 ,
         \DLX_Datapath/RegisterFile/N26705 ,
         \DLX_Datapath/RegisterFile/N26704 ,
         \DLX_Datapath/RegisterFile/N26703 ,
         \DLX_Datapath/RegisterFile/N26702 ,
         \DLX_Datapath/RegisterFile/N26701 ,
         \DLX_Datapath/RegisterFile/N26700 ,
         \DLX_Datapath/RegisterFile/N26699 ,
         \DLX_Datapath/RegisterFile/N26698 ,
         \DLX_Datapath/RegisterFile/N26697 ,
         \DLX_Datapath/RegisterFile/N26696 ,
         \DLX_Datapath/RegisterFile/N26695 ,
         \DLX_Datapath/RegisterFile/N26694 ,
         \DLX_Datapath/RegisterFile/N26693 ,
         \DLX_Datapath/RegisterFile/N26692 ,
         \DLX_Datapath/RegisterFile/N26691 ,
         \DLX_Datapath/RegisterFile/N26690 ,
         \DLX_Datapath/RegisterFile/N26689 ,
         \DLX_Datapath/RegisterFile/N26688 ,
         \DLX_Datapath/RegisterFile/N26687 ,
         \DLX_Datapath/RegisterFile/N26686 ,
         \DLX_Datapath/RegisterFile/N26685 ,
         \DLX_Datapath/RegisterFile/N26684 ,
         \DLX_Datapath/RegisterFile/N26683 ,
         \DLX_Datapath/RegisterFile/N26682 ,
         \DLX_Datapath/RegisterFile/N26681 ,
         \DLX_Datapath/RegisterFile/N26680 ,
         \DLX_Datapath/RegisterFile/N26679 ,
         \DLX_Datapath/RegisterFile/N26678 ,
         \DLX_Datapath/RegisterFile/N26677 ,
         \DLX_Datapath/RegisterFile/N26676 ,
         \DLX_Datapath/RegisterFile/N26675 ,
         \DLX_Datapath/RegisterFile/N26674 ,
         \DLX_Datapath/RegisterFile/N26673 ,
         \DLX_Datapath/RegisterFile/N26672 ,
         \DLX_Datapath/RegisterFile/N26671 ,
         \DLX_Datapath/RegisterFile/N26670 ,
         \DLX_Datapath/RegisterFile/N26669 ,
         \DLX_Datapath/RegisterFile/N26668 ,
         \DLX_Datapath/RegisterFile/N26667 ,
         \DLX_Datapath/RegisterFile/N26634 ,
         \DLX_Datapath/RegisterFile/N26633 ,
         \DLX_Datapath/RegisterFile/N26632 ,
         \DLX_Datapath/RegisterFile/N26631 ,
         \DLX_Datapath/RegisterFile/N26630 ,
         \DLX_Datapath/RegisterFile/N26629 ,
         \DLX_Datapath/RegisterFile/N26628 ,
         \DLX_Datapath/RegisterFile/N26627 ,
         \DLX_Datapath/RegisterFile/N26626 ,
         \DLX_Datapath/RegisterFile/N26625 ,
         \DLX_Datapath/RegisterFile/N26624 ,
         \DLX_Datapath/RegisterFile/N26623 ,
         \DLX_Datapath/RegisterFile/N26622 ,
         \DLX_Datapath/RegisterFile/N26621 ,
         \DLX_Datapath/RegisterFile/N26620 ,
         \DLX_Datapath/RegisterFile/N26619 ,
         \DLX_Datapath/RegisterFile/N26618 ,
         \DLX_Datapath/RegisterFile/N26617 ,
         \DLX_Datapath/RegisterFile/N26616 ,
         \DLX_Datapath/RegisterFile/N26615 ,
         \DLX_Datapath/RegisterFile/N26614 ,
         \DLX_Datapath/RegisterFile/N26613 ,
         \DLX_Datapath/RegisterFile/N26612 ,
         \DLX_Datapath/RegisterFile/N26611 ,
         \DLX_Datapath/RegisterFile/N26610 ,
         \DLX_Datapath/RegisterFile/N26609 ,
         \DLX_Datapath/RegisterFile/N26608 ,
         \DLX_Datapath/RegisterFile/N26607 ,
         \DLX_Datapath/RegisterFile/N26606 ,
         \DLX_Datapath/RegisterFile/N26605 ,
         \DLX_Datapath/RegisterFile/N26604 ,
         \DLX_Datapath/RegisterFile/N26603 ,
         \DLX_Datapath/RegisterFile/N26602 ,
         \DLX_Datapath/RegisterFile/N26601 ,
         \DLX_Datapath/RegisterFile/N26600 ,
         \DLX_Datapath/RegisterFile/N26599 ,
         \DLX_Datapath/RegisterFile/N26598 ,
         \DLX_Datapath/RegisterFile/N26597 ,
         \DLX_Datapath/RegisterFile/N26596 ,
         \DLX_Datapath/RegisterFile/N26595 ,
         \DLX_Datapath/RegisterFile/N26594 ,
         \DLX_Datapath/RegisterFile/N26593 ,
         \DLX_Datapath/RegisterFile/N26592 ,
         \DLX_Datapath/RegisterFile/N26591 ,
         \DLX_Datapath/RegisterFile/N26590 ,
         \DLX_Datapath/RegisterFile/N26589 ,
         \DLX_Datapath/RegisterFile/N26588 ,
         \DLX_Datapath/RegisterFile/N26587 ,
         \DLX_Datapath/RegisterFile/N26586 ,
         \DLX_Datapath/RegisterFile/N26585 ,
         \DLX_Datapath/RegisterFile/N26584 ,
         \DLX_Datapath/RegisterFile/N26583 ,
         \DLX_Datapath/RegisterFile/N26582 ,
         \DLX_Datapath/RegisterFile/N26581 ,
         \DLX_Datapath/RegisterFile/N26580 ,
         \DLX_Datapath/RegisterFile/N26579 ,
         \DLX_Datapath/RegisterFile/N26578 ,
         \DLX_Datapath/RegisterFile/N26577 ,
         \DLX_Datapath/RegisterFile/N26576 ,
         \DLX_Datapath/RegisterFile/N26575 ,
         \DLX_Datapath/RegisterFile/N26574 ,
         \DLX_Datapath/RegisterFile/N26573 ,
         \DLX_Datapath/RegisterFile/N26572 ,
         \DLX_Datapath/RegisterFile/N26571 ,
         \DLX_Datapath/RegisterFile/N26570 ,
         \DLX_Datapath/RegisterFile/N26569 ,
         \DLX_Datapath/RegisterFile/N26568 ,
         \DLX_Datapath/RegisterFile/N26567 ,
         \DLX_Datapath/RegisterFile/N26566 ,
         \DLX_Datapath/RegisterFile/N26565 ,
         \DLX_Datapath/RegisterFile/N26564 ,
         \DLX_Datapath/RegisterFile/N26563 ,
         \DLX_Datapath/RegisterFile/N26562 ,
         \DLX_Datapath/RegisterFile/N26561 ,
         \DLX_Datapath/RegisterFile/N26560 ,
         \DLX_Datapath/RegisterFile/N26559 ,
         \DLX_Datapath/RegisterFile/N26558 ,
         \DLX_Datapath/RegisterFile/N26557 ,
         \DLX_Datapath/RegisterFile/N26556 ,
         \DLX_Datapath/RegisterFile/N26555 ,
         \DLX_Datapath/RegisterFile/N26554 ,
         \DLX_Datapath/RegisterFile/N26553 ,
         \DLX_Datapath/RegisterFile/N26552 ,
         \DLX_Datapath/RegisterFile/N26551 ,
         \DLX_Datapath/RegisterFile/N26550 ,
         \DLX_Datapath/RegisterFile/N26549 ,
         \DLX_Datapath/RegisterFile/N26548 ,
         \DLX_Datapath/RegisterFile/N26547 ,
         \DLX_Datapath/RegisterFile/N26546 ,
         \DLX_Datapath/RegisterFile/N26545 ,
         \DLX_Datapath/RegisterFile/N26544 ,
         \DLX_Datapath/RegisterFile/N26543 ,
         \DLX_Datapath/RegisterFile/N26542 ,
         \DLX_Datapath/RegisterFile/N26541 ,
         \DLX_Datapath/RegisterFile/N26540 ,
         \DLX_Datapath/RegisterFile/N26539 ,
         \DLX_Datapath/RegisterFile/N26538 ,
         \DLX_Datapath/RegisterFile/N26537 ,
         \DLX_Datapath/RegisterFile/N26536 ,
         \DLX_Datapath/RegisterFile/N26535 ,
         \DLX_Datapath/RegisterFile/N26534 ,
         \DLX_Datapath/RegisterFile/N26533 ,
         \DLX_Datapath/RegisterFile/N26532 ,
         \DLX_Datapath/RegisterFile/N26531 ,
         \DLX_Datapath/RegisterFile/N26530 ,
         \DLX_Datapath/RegisterFile/N26529 ,
         \DLX_Datapath/RegisterFile/N26528 ,
         \DLX_Datapath/RegisterFile/N26527 ,
         \DLX_Datapath/RegisterFile/N26526 ,
         \DLX_Datapath/RegisterFile/N26525 ,
         \DLX_Datapath/RegisterFile/N26524 ,
         \DLX_Datapath/RegisterFile/N26523 ,
         \DLX_Datapath/RegisterFile/N26522 ,
         \DLX_Datapath/RegisterFile/N26521 ,
         \DLX_Datapath/RegisterFile/N26520 ,
         \DLX_Datapath/RegisterFile/N26519 ,
         \DLX_Datapath/RegisterFile/N26518 ,
         \DLX_Datapath/RegisterFile/N26517 ,
         \DLX_Datapath/RegisterFile/N26516 ,
         \DLX_Datapath/RegisterFile/N26515 ,
         \DLX_Datapath/RegisterFile/N26514 ,
         \DLX_Datapath/RegisterFile/N26513 ,
         \DLX_Datapath/RegisterFile/N26512 ,
         \DLX_Datapath/RegisterFile/N26511 ,
         \DLX_Datapath/RegisterFile/N26510 ,
         \DLX_Datapath/RegisterFile/N26509 ,
         \DLX_Datapath/RegisterFile/N26508 ,
         \DLX_Datapath/RegisterFile/N26507 ,
         \DLX_Datapath/RegisterFile/N26506 ,
         \DLX_Datapath/RegisterFile/N26505 ,
         \DLX_Datapath/RegisterFile/N26504 ,
         \DLX_Datapath/RegisterFile/N26503 ,
         \DLX_Datapath/RegisterFile/N26502 ,
         \DLX_Datapath/RegisterFile/N26501 ,
         \DLX_Datapath/RegisterFile/N26500 ,
         \DLX_Datapath/RegisterFile/N26499 ,
         \DLX_Datapath/RegisterFile/N26498 ,
         \DLX_Datapath/RegisterFile/N26497 ,
         \DLX_Datapath/RegisterFile/N26496 ,
         \DLX_Datapath/RegisterFile/N26495 ,
         \DLX_Datapath/RegisterFile/N26494 ,
         \DLX_Datapath/RegisterFile/N26493 ,
         \DLX_Datapath/RegisterFile/N26492 ,
         \DLX_Datapath/RegisterFile/N26491 ,
         \DLX_Datapath/RegisterFile/N26490 ,
         \DLX_Datapath/RegisterFile/N26489 ,
         \DLX_Datapath/RegisterFile/N26488 ,
         \DLX_Datapath/RegisterFile/N26487 ,
         \DLX_Datapath/RegisterFile/N26486 ,
         \DLX_Datapath/RegisterFile/N26485 ,
         \DLX_Datapath/RegisterFile/N26484 ,
         \DLX_Datapath/RegisterFile/N26483 ,
         \DLX_Datapath/RegisterFile/N26482 ,
         \DLX_Datapath/RegisterFile/N26481 ,
         \DLX_Datapath/RegisterFile/N26480 ,
         \DLX_Datapath/RegisterFile/N26479 ,
         \DLX_Datapath/RegisterFile/N26478 ,
         \DLX_Datapath/RegisterFile/N26477 ,
         \DLX_Datapath/RegisterFile/N26476 ,
         \DLX_Datapath/RegisterFile/N26475 ,
         \DLX_Datapath/RegisterFile/N26474 ,
         \DLX_Datapath/RegisterFile/N26473 ,
         \DLX_Datapath/RegisterFile/N26472 ,
         \DLX_Datapath/RegisterFile/N26471 ,
         \DLX_Datapath/RegisterFile/N26470 ,
         \DLX_Datapath/RegisterFile/N26469 ,
         \DLX_Datapath/RegisterFile/N26468 ,
         \DLX_Datapath/RegisterFile/N26467 ,
         \DLX_Datapath/RegisterFile/N26466 ,
         \DLX_Datapath/RegisterFile/N26465 ,
         \DLX_Datapath/RegisterFile/N26464 ,
         \DLX_Datapath/RegisterFile/N26463 ,
         \DLX_Datapath/RegisterFile/N26462 ,
         \DLX_Datapath/RegisterFile/N26461 ,
         \DLX_Datapath/RegisterFile/N26460 ,
         \DLX_Datapath/RegisterFile/N26459 ,
         \DLX_Datapath/RegisterFile/N26458 ,
         \DLX_Datapath/RegisterFile/N26457 ,
         \DLX_Datapath/RegisterFile/N26456 ,
         \DLX_Datapath/RegisterFile/N26455 ,
         \DLX_Datapath/RegisterFile/N26454 ,
         \DLX_Datapath/RegisterFile/N26453 ,
         \DLX_Datapath/RegisterFile/N26452 ,
         \DLX_Datapath/RegisterFile/N26451 ,
         \DLX_Datapath/RegisterFile/N26450 ,
         \DLX_Datapath/RegisterFile/N26449 ,
         \DLX_Datapath/RegisterFile/N26448 ,
         \DLX_Datapath/RegisterFile/N26447 ,
         \DLX_Datapath/RegisterFile/N26446 ,
         \DLX_Datapath/RegisterFile/N26445 ,
         \DLX_Datapath/RegisterFile/N26444 ,
         \DLX_Datapath/RegisterFile/N26443 ,
         \DLX_Datapath/RegisterFile/N26442 ,
         \DLX_Datapath/RegisterFile/N26441 ,
         \DLX_Datapath/RegisterFile/N26440 ,
         \DLX_Datapath/RegisterFile/N26439 ,
         \DLX_Datapath/RegisterFile/N26438 ,
         \DLX_Datapath/RegisterFile/N26437 ,
         \DLX_Datapath/RegisterFile/N26436 ,
         \DLX_Datapath/RegisterFile/N26435 ,
         \DLX_Datapath/RegisterFile/N26434 ,
         \DLX_Datapath/RegisterFile/N26433 ,
         \DLX_Datapath/RegisterFile/N26432 ,
         \DLX_Datapath/RegisterFile/N26431 ,
         \DLX_Datapath/RegisterFile/N26430 ,
         \DLX_Datapath/RegisterFile/N26429 ,
         \DLX_Datapath/RegisterFile/N26428 ,
         \DLX_Datapath/RegisterFile/N26427 ,
         \DLX_Datapath/RegisterFile/N26426 ,
         \DLX_Datapath/RegisterFile/N26425 ,
         \DLX_Datapath/RegisterFile/N26424 ,
         \DLX_Datapath/RegisterFile/N26423 ,
         \DLX_Datapath/RegisterFile/N26422 ,
         \DLX_Datapath/RegisterFile/N26421 ,
         \DLX_Datapath/RegisterFile/N26420 ,
         \DLX_Datapath/RegisterFile/N26419 ,
         \DLX_Datapath/RegisterFile/N26418 ,
         \DLX_Datapath/RegisterFile/N26417 ,
         \DLX_Datapath/RegisterFile/N26416 ,
         \DLX_Datapath/RegisterFile/N26415 ,
         \DLX_Datapath/RegisterFile/N26414 ,
         \DLX_Datapath/RegisterFile/N26413 ,
         \DLX_Datapath/RegisterFile/N26412 ,
         \DLX_Datapath/RegisterFile/N26411 ,
         \DLX_Datapath/RegisterFile/N26410 ,
         \DLX_Datapath/RegisterFile/N26409 ,
         \DLX_Datapath/RegisterFile/N26408 ,
         \DLX_Datapath/RegisterFile/N26407 ,
         \DLX_Datapath/RegisterFile/N26406 ,
         \DLX_Datapath/RegisterFile/N26405 ,
         \DLX_Datapath/RegisterFile/N26404 ,
         \DLX_Datapath/RegisterFile/N26403 ,
         \DLX_Datapath/RegisterFile/N26402 ,
         \DLX_Datapath/RegisterFile/N26401 ,
         \DLX_Datapath/RegisterFile/N26400 ,
         \DLX_Datapath/RegisterFile/N26399 ,
         \DLX_Datapath/RegisterFile/N26398 ,
         \DLX_Datapath/RegisterFile/N26397 ,
         \DLX_Datapath/RegisterFile/N26396 ,
         \DLX_Datapath/RegisterFile/N26395 ,
         \DLX_Datapath/RegisterFile/N26394 ,
         \DLX_Datapath/RegisterFile/N26393 ,
         \DLX_Datapath/RegisterFile/N26392 ,
         \DLX_Datapath/RegisterFile/N26391 ,
         \DLX_Datapath/RegisterFile/N26390 ,
         \DLX_Datapath/RegisterFile/N26389 ,
         \DLX_Datapath/RegisterFile/N26388 ,
         \DLX_Datapath/RegisterFile/N26387 ,
         \DLX_Datapath/RegisterFile/N26386 ,
         \DLX_Datapath/RegisterFile/N26385 ,
         \DLX_Datapath/RegisterFile/N26384 ,
         \DLX_Datapath/RegisterFile/N26383 ,
         \DLX_Datapath/RegisterFile/N26382 ,
         \DLX_Datapath/RegisterFile/N26381 ,
         \DLX_Datapath/RegisterFile/N26380 ,
         \DLX_Datapath/RegisterFile/N26379 ,
         \DLX_Datapath/RegisterFile/N26378 ,
         \DLX_Datapath/RegisterFile/N26377 ,
         \DLX_Datapath/RegisterFile/N26376 ,
         \DLX_Datapath/RegisterFile/N26375 ,
         \DLX_Datapath/RegisterFile/N26374 ,
         \DLX_Datapath/RegisterFile/N26373 ,
         \DLX_Datapath/RegisterFile/N26372 ,
         \DLX_Datapath/RegisterFile/N26371 ,
         \DLX_Datapath/RegisterFile/N26370 ,
         \DLX_Datapath/RegisterFile/N26369 ,
         \DLX_Datapath/RegisterFile/N26368 ,
         \DLX_Datapath/RegisterFile/N26367 ,
         \DLX_Datapath/RegisterFile/N26366 ,
         \DLX_Datapath/RegisterFile/N26365 ,
         \DLX_Datapath/RegisterFile/N26364 ,
         \DLX_Datapath/RegisterFile/N26363 ,
         \DLX_Datapath/RegisterFile/N26362 ,
         \DLX_Datapath/RegisterFile/N26361 ,
         \DLX_Datapath/RegisterFile/N26360 ,
         \DLX_Datapath/RegisterFile/N26359 ,
         \DLX_Datapath/RegisterFile/N26358 ,
         \DLX_Datapath/RegisterFile/N26357 ,
         \DLX_Datapath/RegisterFile/N26356 ,
         \DLX_Datapath/RegisterFile/N26355 ,
         \DLX_Datapath/RegisterFile/N26354 ,
         \DLX_Datapath/RegisterFile/N26353 ,
         \DLX_Datapath/RegisterFile/N26352 ,
         \DLX_Datapath/RegisterFile/N26351 ,
         \DLX_Datapath/RegisterFile/N26350 ,
         \DLX_Datapath/RegisterFile/N26349 ,
         \DLX_Datapath/RegisterFile/N26348 ,
         \DLX_Datapath/RegisterFile/N26347 ,
         \DLX_Datapath/RegisterFile/N26346 ,
         \DLX_Datapath/RegisterFile/N26345 ,
         \DLX_Datapath/RegisterFile/N26344 ,
         \DLX_Datapath/RegisterFile/N26343 ,
         \DLX_Datapath/RegisterFile/N26342 ,
         \DLX_Datapath/RegisterFile/N26341 ,
         \DLX_Datapath/RegisterFile/N26340 ,
         \DLX_Datapath/RegisterFile/N26339 ,
         \DLX_Datapath/RegisterFile/N26338 ,
         \DLX_Datapath/RegisterFile/N26337 ,
         \DLX_Datapath/RegisterFile/N26336 ,
         \DLX_Datapath/RegisterFile/N26335 ,
         \DLX_Datapath/RegisterFile/N26334 ,
         \DLX_Datapath/RegisterFile/N26333 ,
         \DLX_Datapath/RegisterFile/N26332 ,
         \DLX_Datapath/RegisterFile/N26331 ,
         \DLX_Datapath/RegisterFile/N26330 ,
         \DLX_Datapath/RegisterFile/N26329 ,
         \DLX_Datapath/RegisterFile/N26328 ,
         \DLX_Datapath/RegisterFile/N26327 ,
         \DLX_Datapath/RegisterFile/N26326 ,
         \DLX_Datapath/RegisterFile/N26325 ,
         \DLX_Datapath/RegisterFile/N26324 ,
         \DLX_Datapath/RegisterFile/N26323 ,
         \DLX_Datapath/RegisterFile/N26322 ,
         \DLX_Datapath/RegisterFile/N26321 ,
         \DLX_Datapath/RegisterFile/N26320 ,
         \DLX_Datapath/RegisterFile/N26319 ,
         \DLX_Datapath/RegisterFile/N26318 ,
         \DLX_Datapath/RegisterFile/N26317 ,
         \DLX_Datapath/RegisterFile/N26316 ,
         \DLX_Datapath/RegisterFile/N26315 ,
         \DLX_Datapath/RegisterFile/N26314 ,
         \DLX_Datapath/RegisterFile/N26313 ,
         \DLX_Datapath/RegisterFile/N26312 ,
         \DLX_Datapath/RegisterFile/N26311 ,
         \DLX_Datapath/RegisterFile/N26310 ,
         \DLX_Datapath/RegisterFile/N26309 ,
         \DLX_Datapath/RegisterFile/N26308 ,
         \DLX_Datapath/RegisterFile/N26307 ,
         \DLX_Datapath/RegisterFile/N26306 ,
         \DLX_Datapath/RegisterFile/N26305 ,
         \DLX_Datapath/RegisterFile/N26304 ,
         \DLX_Datapath/RegisterFile/N26303 ,
         \DLX_Datapath/RegisterFile/N26302 ,
         \DLX_Datapath/RegisterFile/N26301 ,
         \DLX_Datapath/RegisterFile/N26300 ,
         \DLX_Datapath/RegisterFile/N26299 ,
         \DLX_Datapath/RegisterFile/N26294 ,
         \DLX_Datapath/RegisterFile/N26292 ,
         \DLX_Datapath/RegisterFile/N26291 ,
         \DLX_Datapath/RegisterFile/N26290 ,
         \DLX_Datapath/RegisterFile/N26289 ,
         \DLX_Datapath/RegisterFile/N26288 ,
         \DLX_Datapath/RegisterFile/N26287 ,
         \DLX_Datapath/RegisterFile/N26286 ,
         \DLX_Datapath/RegisterFile/N26285 ,
         \DLX_Datapath/RegisterFile/N26284 ,
         \DLX_Datapath/RegisterFile/N26283 ,
         \DLX_Datapath/RegisterFile/N26282 ,
         \DLX_Datapath/RegisterFile/N26281 ,
         \DLX_Datapath/RegisterFile/N26280 ,
         \DLX_Datapath/RegisterFile/N26279 ,
         \DLX_Datapath/RegisterFile/N26278 ,
         \DLX_Datapath/RegisterFile/N26277 ,
         \DLX_Datapath/RegisterFile/N26276 ,
         \DLX_Datapath/RegisterFile/N26275 ,
         \DLX_Datapath/RegisterFile/N26274 ,
         \DLX_Datapath/RegisterFile/N26273 ,
         \DLX_Datapath/RegisterFile/N26272 ,
         \DLX_Datapath/RegisterFile/N26271 ,
         \DLX_Datapath/RegisterFile/N26270 ,
         \DLX_Datapath/RegisterFile/N26269 ,
         \DLX_Datapath/RegisterFile/N26268 ,
         \DLX_Datapath/RegisterFile/N26267 ,
         \DLX_Datapath/RegisterFile/N26266 ,
         \DLX_Datapath/RegisterFile/N26265 ,
         \DLX_Datapath/RegisterFile/N26264 ,
         \DLX_Datapath/RegisterFile/N26263 ,
         \DLX_Datapath/RegisterFile/N26262 ,
         \DLX_Datapath/RegisterFile/N26261 ,
         \DLX_Datapath/RegisterFile/N26260 ,
         \DLX_Datapath/RegisterFile/N26259 ,
         \DLX_Datapath/RegisterFile/N26258 ,
         \DLX_Datapath/RegisterFile/N26257 ,
         \DLX_Datapath/RegisterFile/N26256 ,
         \DLX_Datapath/RegisterFile/N26255 ,
         \DLX_Datapath/RegisterFile/N26254 ,
         \DLX_Datapath/RegisterFile/N26253 ,
         \DLX_Datapath/RegisterFile/N26252 ,
         \DLX_Datapath/RegisterFile/N26251 ,
         \DLX_Datapath/RegisterFile/N26250 ,
         \DLX_Datapath/RegisterFile/N26249 ,
         \DLX_Datapath/RegisterFile/N26248 ,
         \DLX_Datapath/RegisterFile/N26247 ,
         \DLX_Datapath/RegisterFile/N26246 ,
         \DLX_Datapath/RegisterFile/N26245 ,
         \DLX_Datapath/RegisterFile/N26244 ,
         \DLX_Datapath/RegisterFile/N26243 ,
         \DLX_Datapath/RegisterFile/N26242 ,
         \DLX_Datapath/RegisterFile/N26241 ,
         \DLX_Datapath/RegisterFile/N26240 ,
         \DLX_Datapath/RegisterFile/N26239 ,
         \DLX_Datapath/RegisterFile/N26238 ,
         \DLX_Datapath/RegisterFile/N26237 ,
         \DLX_Datapath/RegisterFile/N26236 ,
         \DLX_Datapath/RegisterFile/N26235 ,
         \DLX_Datapath/RegisterFile/N26234 ,
         \DLX_Datapath/RegisterFile/N26233 ,
         \DLX_Datapath/RegisterFile/N26232 ,
         \DLX_Datapath/RegisterFile/N26231 ,
         \DLX_Datapath/RegisterFile/N26230 ,
         \DLX_Datapath/RegisterFile/N26229 ,
         \DLX_Datapath/RegisterFile/N26228 ,
         \DLX_Datapath/RegisterFile/N26227 ,
         \DLX_Datapath/RegisterFile/N26226 ,
         \DLX_Datapath/RegisterFile/N26225 ,
         \DLX_Datapath/RegisterFile/N26224 ,
         \DLX_Datapath/RegisterFile/N26223 ,
         \DLX_Datapath/RegisterFile/N26222 ,
         \DLX_Datapath/RegisterFile/N26221 ,
         \DLX_Datapath/RegisterFile/N26220 ,
         \DLX_Datapath/RegisterFile/N26219 ,
         \DLX_Datapath/RegisterFile/N26218 ,
         \DLX_Datapath/RegisterFile/N26217 ,
         \DLX_Datapath/RegisterFile/N26216 ,
         \DLX_Datapath/RegisterFile/N26215 ,
         \DLX_Datapath/RegisterFile/N26214 ,
         \DLX_Datapath/RegisterFile/N26213 ,
         \DLX_Datapath/RegisterFile/N26212 ,
         \DLX_Datapath/RegisterFile/N26211 ,
         \DLX_Datapath/RegisterFile/N26210 ,
         \DLX_Datapath/RegisterFile/N26209 ,
         \DLX_Datapath/RegisterFile/N26208 ,
         \DLX_Datapath/RegisterFile/N26207 ,
         \DLX_Datapath/RegisterFile/N26206 ,
         \DLX_Datapath/RegisterFile/N26205 ,
         \DLX_Datapath/RegisterFile/N26204 ,
         \DLX_Datapath/RegisterFile/N26203 ,
         \DLX_Datapath/RegisterFile/N26202 ,
         \DLX_Datapath/RegisterFile/N26201 ,
         \DLX_Datapath/RegisterFile/N26200 ,
         \DLX_Datapath/RegisterFile/N26199 ,
         \DLX_Datapath/RegisterFile/N26198 ,
         \DLX_Datapath/RegisterFile/N26197 ,
         \DLX_Datapath/RegisterFile/N26196 ,
         \DLX_Datapath/RegisterFile/N26195 ,
         \DLX_Datapath/RegisterFile/N26194 ,
         \DLX_Datapath/RegisterFile/N26193 ,
         \DLX_Datapath/RegisterFile/N26192 ,
         \DLX_Datapath/RegisterFile/N26191 ,
         \DLX_Datapath/RegisterFile/N26190 ,
         \DLX_Datapath/RegisterFile/N26189 ,
         \DLX_Datapath/RegisterFile/N26188 ,
         \DLX_Datapath/RegisterFile/N26187 ,
         \DLX_Datapath/RegisterFile/N26179 ,
         \DLX_Datapath/RegisterFile/N26178 ,
         \DLX_Datapath/RegisterFile/N26176 ,
         \DLX_Datapath/RegisterFile/N26172 ,
         \DLX_Datapath/RegisterFile/N26171 ,
         \DLX_Datapath/RegisterFile/N26170 ,
         \DLX_Datapath/RegisterFile/N26169 ,
         \DLX_Datapath/RegisterFile/N26168 ,
         \DLX_Datapath/RegisterFile/N26167 ,
         \DLX_Datapath/RegisterFile/N26166 ,
         \DLX_Datapath/RegisterFile/N26165 ,
         \DLX_Datapath/RegisterFile/N26164 ,
         \DLX_Datapath/RegisterFile/N26163 ,
         \DLX_Datapath/RegisterFile/N26162 ,
         \DLX_Datapath/RegisterFile/N26161 ,
         \DLX_Datapath/RegisterFile/N26160 ,
         \DLX_Datapath/RegisterFile/N26159 ,
         \DLX_Datapath/RegisterFile/N26158 ,
         \DLX_Datapath/RegisterFile/N26157 ,
         \DLX_Datapath/RegisterFile/N26156 ,
         \DLX_Datapath/RegisterFile/N26155 ,
         \DLX_Datapath/RegisterFile/N26154 ,
         \DLX_Datapath/RegisterFile/N26153 ,
         \DLX_Datapath/RegisterFile/N26152 ,
         \DLX_Datapath/RegisterFile/N26151 ,
         \DLX_Datapath/RegisterFile/N26150 ,
         \DLX_Datapath/RegisterFile/N26149 ,
         \DLX_Datapath/RegisterFile/N26148 ,
         \DLX_Datapath/RegisterFile/N26147 ,
         \DLX_Datapath/RegisterFile/N26146 ,
         \DLX_Datapath/RegisterFile/N26145 ,
         \DLX_Datapath/RegisterFile/N26144 ,
         \DLX_Datapath/RegisterFile/N26143 ,
         \DLX_Datapath/RegisterFile/N26142 ,
         \DLX_Datapath/RegisterFile/N26141 ,
         \DLX_Datapath/RegisterFile/N26140 ,
         \DLX_Datapath/RegisterFile/N26139 ,
         \DLX_Datapath/RegisterFile/N26138 ,
         \DLX_Datapath/RegisterFile/N26137 ,
         \DLX_Datapath/RegisterFile/N26136 ,
         \DLX_Datapath/RegisterFile/N26135 ,
         \DLX_Datapath/RegisterFile/N26134 ,
         \DLX_Datapath/RegisterFile/N26133 ,
         \DLX_Datapath/RegisterFile/N26132 ,
         \DLX_Datapath/RegisterFile/N26131 ,
         \DLX_Datapath/RegisterFile/N26130 ,
         \DLX_Datapath/RegisterFile/N26129 ,
         \DLX_Datapath/RegisterFile/N26128 ,
         \DLX_Datapath/RegisterFile/N26127 ,
         \DLX_Datapath/RegisterFile/N26126 ,
         \DLX_Datapath/RegisterFile/N26125 ,
         \DLX_Datapath/RegisterFile/N26124 ,
         \DLX_Datapath/RegisterFile/N26123 ,
         \DLX_Datapath/RegisterFile/N26122 ,
         \DLX_Datapath/RegisterFile/N26121 ,
         \DLX_Datapath/RegisterFile/N26120 ,
         \DLX_Datapath/RegisterFile/N26119 ,
         \DLX_Datapath/RegisterFile/N26118 ,
         \DLX_Datapath/RegisterFile/N26117 ,
         \DLX_Datapath/RegisterFile/N26116 ,
         \DLX_Datapath/RegisterFile/N26115 ,
         \DLX_Datapath/RegisterFile/N26114 ,
         \DLX_Datapath/RegisterFile/N26113 ,
         \DLX_Datapath/RegisterFile/N26112 ,
         \DLX_Datapath/RegisterFile/N26111 ,
         \DLX_Datapath/RegisterFile/N26110 ,
         \DLX_Datapath/RegisterFile/N26109 ,
         \DLX_Datapath/RegisterFile/N26108 ,
         \DLX_Datapath/RegisterFile/N26107 ,
         \DLX_Datapath/RegisterFile/N26106 ,
         \DLX_Datapath/RegisterFile/N26105 ,
         \DLX_Datapath/RegisterFile/N26104 ,
         \DLX_Datapath/RegisterFile/N26103 ,
         \DLX_Datapath/RegisterFile/N26102 ,
         \DLX_Datapath/RegisterFile/N26101 ,
         \DLX_Datapath/RegisterFile/N26100 ,
         \DLX_Datapath/RegisterFile/N26099 ,
         \DLX_Datapath/RegisterFile/N26098 ,
         \DLX_Datapath/RegisterFile/N26097 ,
         \DLX_Datapath/RegisterFile/N26096 ,
         \DLX_Datapath/RegisterFile/N26095 ,
         \DLX_Datapath/RegisterFile/N26094 ,
         \DLX_Datapath/RegisterFile/N26093 ,
         \DLX_Datapath/RegisterFile/N26092 ,
         \DLX_Datapath/RegisterFile/N26091 ,
         \DLX_Datapath/RegisterFile/N26090 ,
         \DLX_Datapath/RegisterFile/N26089 ,
         \DLX_Datapath/RegisterFile/N26088 ,
         \DLX_Datapath/RegisterFile/N26087 ,
         \DLX_Datapath/RegisterFile/N26086 ,
         \DLX_Datapath/RegisterFile/N26085 ,
         \DLX_Datapath/RegisterFile/N26084 ,
         \DLX_Datapath/RegisterFile/N26083 ,
         \DLX_Datapath/RegisterFile/N26082 ,
         \DLX_Datapath/RegisterFile/N26081 ,
         \DLX_Datapath/RegisterFile/N26080 ,
         \DLX_Datapath/RegisterFile/N26079 ,
         \DLX_Datapath/RegisterFile/N26078 ,
         \DLX_Datapath/RegisterFile/N26077 ,
         \DLX_Datapath/RegisterFile/N26076 ,
         \DLX_Datapath/RegisterFile/N26075 ,
         \DLX_Datapath/RegisterFile/N26074 ,
         \DLX_Datapath/RegisterFile/N26073 ,
         \DLX_Datapath/RegisterFile/N26072 ,
         \DLX_Datapath/RegisterFile/N26071 ,
         \DLX_Datapath/RegisterFile/N26070 ,
         \DLX_Datapath/RegisterFile/N26069 ,
         \DLX_Datapath/RegisterFile/N26068 ,
         \DLX_Datapath/RegisterFile/N26067 ,
         \DLX_Datapath/RegisterFile/N26066 ,
         \DLX_Datapath/RegisterFile/N26065 ,
         \DLX_Datapath/RegisterFile/N26064 ,
         \DLX_Datapath/RegisterFile/N26063 ,
         \DLX_Datapath/RegisterFile/N26062 ,
         \DLX_Datapath/RegisterFile/N26061 ,
         \DLX_Datapath/RegisterFile/N26060 ,
         \DLX_Datapath/RegisterFile/N26059 ,
         \DLX_Datapath/RegisterFile/N26058 ,
         \DLX_Datapath/RegisterFile/N26057 ,
         \DLX_Datapath/RegisterFile/N26056 ,
         \DLX_Datapath/RegisterFile/N26055 ,
         \DLX_Datapath/RegisterFile/N26054 ,
         \DLX_Datapath/RegisterFile/N26053 ,
         \DLX_Datapath/RegisterFile/N26052 ,
         \DLX_Datapath/RegisterFile/N26051 ,
         \DLX_Datapath/RegisterFile/N26050 ,
         \DLX_Datapath/RegisterFile/N26049 ,
         \DLX_Datapath/RegisterFile/N26048 ,
         \DLX_Datapath/RegisterFile/N26047 ,
         \DLX_Datapath/RegisterFile/N26046 ,
         \DLX_Datapath/RegisterFile/N26045 ,
         \DLX_Datapath/RegisterFile/N26044 ,
         \DLX_Datapath/RegisterFile/N26043 ,
         \DLX_Datapath/RegisterFile/N26038 ,
         \DLX_Datapath/RegisterFile/N26036 ,
         \DLX_Datapath/RegisterFile/N26034 ,
         \DLX_Datapath/RegisterFile/N26033 ,
         \DLX_Datapath/RegisterFile/N26031 ,
         \DLX_Datapath/RegisterFile/N26026 ,
         \DLX_Datapath/RegisterFile/N26025 ,
         \DLX_Datapath/RegisterFile/N26024 ,
         \DLX_Datapath/RegisterFile/N26023 ,
         \DLX_Datapath/RegisterFile/N26022 ,
         \DLX_Datapath/RegisterFile/N26021 ,
         \DLX_Datapath/RegisterFile/N26020 ,
         \DLX_Datapath/RegisterFile/N26019 ,
         \DLX_Datapath/RegisterFile/N26018 ,
         \DLX_Datapath/RegisterFile/N26017 ,
         \DLX_Datapath/RegisterFile/N26016 ,
         \DLX_Datapath/RegisterFile/N26015 ,
         \DLX_Datapath/RegisterFile/N26014 ,
         \DLX_Datapath/RegisterFile/N26013 ,
         \DLX_Datapath/RegisterFile/N26012 ,
         \DLX_Datapath/RegisterFile/N26011 ,
         \DLX_Datapath/RegisterFile/N26010 ,
         \DLX_Datapath/RegisterFile/N26009 ,
         \DLX_Datapath/RegisterFile/N26008 ,
         \DLX_Datapath/RegisterFile/N26007 ,
         \DLX_Datapath/RegisterFile/N26006 ,
         \DLX_Datapath/RegisterFile/N26005 ,
         \DLX_Datapath/RegisterFile/N26004 ,
         \DLX_Datapath/RegisterFile/N26003 ,
         \DLX_Datapath/RegisterFile/N26002 ,
         \DLX_Datapath/RegisterFile/N26001 ,
         \DLX_Datapath/RegisterFile/N26000 ,
         \DLX_Datapath/RegisterFile/N25999 ,
         \DLX_Datapath/RegisterFile/N25998 ,
         \DLX_Datapath/RegisterFile/N25997 ,
         \DLX_Datapath/RegisterFile/N25996 ,
         \DLX_Datapath/RegisterFile/N25995 ,
         \DLX_Datapath/RegisterFile/N25994 ,
         \DLX_Datapath/RegisterFile/N25993 ,
         \DLX_Datapath/RegisterFile/N25992 ,
         \DLX_Datapath/RegisterFile/N25991 ,
         \DLX_Datapath/RegisterFile/N25990 ,
         \DLX_Datapath/RegisterFile/N25989 ,
         \DLX_Datapath/RegisterFile/N25988 ,
         \DLX_Datapath/RegisterFile/N25987 ,
         \DLX_Datapath/RegisterFile/N25986 ,
         \DLX_Datapath/RegisterFile/N25985 ,
         \DLX_Datapath/RegisterFile/N25984 ,
         \DLX_Datapath/RegisterFile/N25983 ,
         \DLX_Datapath/RegisterFile/N25982 ,
         \DLX_Datapath/RegisterFile/N25981 ,
         \DLX_Datapath/RegisterFile/N25980 ,
         \DLX_Datapath/RegisterFile/N25979 ,
         \DLX_Datapath/RegisterFile/N25978 ,
         \DLX_Datapath/RegisterFile/N25977 ,
         \DLX_Datapath/RegisterFile/N25976 ,
         \DLX_Datapath/RegisterFile/N25975 ,
         \DLX_Datapath/RegisterFile/N25974 ,
         \DLX_Datapath/RegisterFile/N25973 ,
         \DLX_Datapath/RegisterFile/N25972 ,
         \DLX_Datapath/RegisterFile/N25971 ,
         \DLX_Datapath/RegisterFile/N25970 ,
         \DLX_Datapath/RegisterFile/N25968 ,
         \DLX_Datapath/RegisterFile/N25967 ,
         \DLX_Datapath/RegisterFile/N25966 ,
         \DLX_Datapath/RegisterFile/N25964 ,
         \DLX_Datapath/RegisterFile/N25963 ,
         \DLX_Datapath/RegisterFile/N25962 ,
         \DLX_Datapath/RegisterFile/N25961 ,
         \DLX_Datapath/RegisterFile/N25960 ,
         \DLX_Datapath/RegisterFile/N25959 ,
         \DLX_Datapath/RegisterFile/N25958 ,
         \DLX_Datapath/RegisterFile/N25957 ,
         \DLX_Datapath/RegisterFile/N25956 ,
         \DLX_Datapath/RegisterFile/N25955 ,
         \DLX_Datapath/RegisterFile/N25954 ,
         \DLX_Datapath/RegisterFile/N25953 ,
         \DLX_Datapath/RegisterFile/N25952 ,
         \DLX_Datapath/RegisterFile/N25951 ,
         \DLX_Datapath/RegisterFile/N25950 ,
         \DLX_Datapath/RegisterFile/N25949 ,
         \DLX_Datapath/RegisterFile/N25948 ,
         \DLX_Datapath/RegisterFile/N25947 ,
         \DLX_Datapath/RegisterFile/N25946 ,
         \DLX_Datapath/RegisterFile/N25945 ,
         \DLX_Datapath/RegisterFile/N25944 ,
         \DLX_Datapath/RegisterFile/N25943 ,
         \DLX_Datapath/RegisterFile/N25942 ,
         \DLX_Datapath/RegisterFile/N25941 ,
         \DLX_Datapath/RegisterFile/N25940 ,
         \DLX_Datapath/RegisterFile/N25939 ,
         \DLX_Datapath/RegisterFile/N25938 ,
         \DLX_Datapath/RegisterFile/N25937 ,
         \DLX_Datapath/RegisterFile/N25936 ,
         \DLX_Datapath/RegisterFile/N25935 ,
         \DLX_Datapath/RegisterFile/N25934 ,
         \DLX_Datapath/RegisterFile/N25933 ,
         \DLX_Datapath/RegisterFile/N25932 ,
         \DLX_Datapath/RegisterFile/N25931 ,
         \DLX_Datapath/RegisterFile/N25926 ,
         \DLX_Datapath/RegisterFile/N25924 ,
         \DLX_Datapath/RegisterFile/N25922 ,
         \DLX_Datapath/RegisterFile/N25920 ,
         \DLX_Datapath/RegisterFile/N25919 ,
         \DLX_Datapath/RegisterFile/N25898 ,
         \DLX_Datapath/RegisterFile/N25897 ,
         \DLX_Datapath/RegisterFile/N25896 ,
         \DLX_Datapath/RegisterFile/N25895 ,
         \DLX_Datapath/RegisterFile/N25894 ,
         \DLX_Datapath/RegisterFile/N25893 ,
         \DLX_Datapath/RegisterFile/N25892 ,
         \DLX_Datapath/RegisterFile/N25891 ,
         \DLX_Datapath/RegisterFile/N25890 ,
         \DLX_Datapath/RegisterFile/N25889 ,
         \DLX_Datapath/RegisterFile/N25888 ,
         \DLX_Datapath/RegisterFile/N25887 ,
         \DLX_Datapath/RegisterFile/N25886 ,
         \DLX_Datapath/RegisterFile/N25885 ,
         \DLX_Datapath/RegisterFile/N25884 ,
         \DLX_Datapath/RegisterFile/N25883 ,
         \DLX_Datapath/RegisterFile/N25882 ,
         \DLX_Datapath/RegisterFile/N25881 ,
         \DLX_Datapath/RegisterFile/N25880 ,
         \DLX_Datapath/RegisterFile/N25879 ,
         \DLX_Datapath/RegisterFile/N25878 ,
         \DLX_Datapath/RegisterFile/N25877 ,
         \DLX_Datapath/RegisterFile/N25876 ,
         \DLX_Datapath/RegisterFile/N25875 ,
         \DLX_Datapath/RegisterFile/N25874 ,
         \DLX_Datapath/RegisterFile/N25873 ,
         \DLX_Datapath/RegisterFile/N25872 ,
         \DLX_Datapath/RegisterFile/N25871 ,
         \DLX_Datapath/RegisterFile/N25870 ,
         \DLX_Datapath/RegisterFile/N25869 ,
         \DLX_Datapath/RegisterFile/N25868 ,
         \DLX_Datapath/RegisterFile/N25867 ,
         \DLX_Datapath/RegisterFile/N25866 ,
         \DLX_Datapath/RegisterFile/N25865 ,
         \DLX_Datapath/RegisterFile/N25864 ,
         \DLX_Datapath/RegisterFile/N25863 ,
         \DLX_Datapath/RegisterFile/N25862 ,
         \DLX_Datapath/RegisterFile/N25861 ,
         \DLX_Datapath/RegisterFile/N25860 ,
         \DLX_Datapath/RegisterFile/N25859 ,
         \DLX_Datapath/RegisterFile/N25858 ,
         \DLX_Datapath/RegisterFile/N25857 ,
         \DLX_Datapath/RegisterFile/N25856 ,
         \DLX_Datapath/RegisterFile/N25855 ,
         \DLX_Datapath/RegisterFile/N25854 ,
         \DLX_Datapath/RegisterFile/N25853 ,
         \DLX_Datapath/RegisterFile/N25852 ,
         \DLX_Datapath/RegisterFile/N25851 ,
         \DLX_Datapath/RegisterFile/N25850 ,
         \DLX_Datapath/RegisterFile/N25849 ,
         \DLX_Datapath/RegisterFile/N25848 ,
         \DLX_Datapath/RegisterFile/N25847 ,
         \DLX_Datapath/RegisterFile/N25846 ,
         \DLX_Datapath/RegisterFile/N25845 ,
         \DLX_Datapath/RegisterFile/N25844 ,
         \DLX_Datapath/RegisterFile/N25843 ,
         \DLX_Datapath/RegisterFile/N25842 ,
         \DLX_Datapath/RegisterFile/N25841 ,
         \DLX_Datapath/RegisterFile/N25840 ,
         \DLX_Datapath/RegisterFile/N25839 ,
         \DLX_Datapath/RegisterFile/N25838 ,
         \DLX_Datapath/RegisterFile/N25837 ,
         \DLX_Datapath/RegisterFile/N25836 ,
         \DLX_Datapath/RegisterFile/N25835 ,
         \DLX_Datapath/RegisterFile/N25834 ,
         \DLX_Datapath/RegisterFile/N25833 ,
         \DLX_Datapath/RegisterFile/N25832 ,
         \DLX_Datapath/RegisterFile/N25831 ,
         \DLX_Datapath/RegisterFile/N25830 ,
         \DLX_Datapath/RegisterFile/N25829 ,
         \DLX_Datapath/RegisterFile/N25828 ,
         \DLX_Datapath/RegisterFile/N25827 ,
         \DLX_Datapath/RegisterFile/N25826 ,
         \DLX_Datapath/RegisterFile/N25825 ,
         \DLX_Datapath/RegisterFile/N25824 ,
         \DLX_Datapath/RegisterFile/N25823 ,
         \DLX_Datapath/RegisterFile/N25822 ,
         \DLX_Datapath/RegisterFile/N25821 ,
         \DLX_Datapath/RegisterFile/N25820 ,
         \DLX_Datapath/RegisterFile/N25819 ,
         \DLX_Datapath/RegisterFile/N25818 ,
         \DLX_Datapath/RegisterFile/N25817 ,
         \DLX_Datapath/RegisterFile/N25816 ,
         \DLX_Datapath/RegisterFile/N25815 ,
         \DLX_Datapath/RegisterFile/N25814 ,
         \DLX_Datapath/RegisterFile/N25813 ,
         \DLX_Datapath/RegisterFile/N25812 ,
         \DLX_Datapath/RegisterFile/N25811 ,
         \DLX_Datapath/RegisterFile/N25810 ,
         \DLX_Datapath/RegisterFile/N25809 ,
         \DLX_Datapath/RegisterFile/N25808 ,
         \DLX_Datapath/RegisterFile/N25807 ,
         \DLX_Datapath/RegisterFile/N25806 ,
         \DLX_Datapath/RegisterFile/N25805 ,
         \DLX_Datapath/RegisterFile/N25804 ,
         \DLX_Datapath/RegisterFile/N25803 ,
         \DLX_Datapath/RegisterFile/N25802 ,
         \DLX_Datapath/RegisterFile/N25800 ,
         \DLX_Datapath/RegisterFile/N25799 ,
         \DLX_Datapath/RegisterFile/N25798 ,
         \DLX_Datapath/RegisterFile/N25797 ,
         \DLX_Datapath/RegisterFile/N25796 ,
         \DLX_Datapath/RegisterFile/N25795 ,
         \DLX_Datapath/RegisterFile/N25794 ,
         \DLX_Datapath/RegisterFile/N25793 ,
         \DLX_Datapath/RegisterFile/N25792 ,
         \DLX_Datapath/RegisterFile/N25791 ,
         \DLX_Datapath/RegisterFile/N25790 ,
         \DLX_Datapath/RegisterFile/N25789 ,
         \DLX_Datapath/RegisterFile/N25788 ,
         \DLX_Datapath/RegisterFile/N25787 ,
         \DLX_Datapath/RegisterFile/N25785 ,
         \DLX_Datapath/RegisterFile/N25784 ,
         \DLX_Datapath/RegisterFile/N25783 ,
         \DLX_Datapath/RegisterFile/N25782 ,
         \DLX_Datapath/RegisterFile/N25780 ,
         \DLX_Datapath/RegisterFile/N25779 ,
         \DLX_Datapath/RegisterFile/N25778 ,
         \DLX_Datapath/RegisterFile/N25777 ,
         \DLX_Datapath/RegisterFile/N25776 ,
         \DLX_Datapath/RegisterFile/N25775 ,
         \DLX_Datapath/RegisterFile/N25771 ,
         \DLX_Datapath/RegisterFile/N25770 ,
         \DLX_Datapath/RegisterFile/N25769 ,
         \DLX_Datapath/RegisterFile/N25768 ,
         \DLX_Datapath/RegisterFile/N25767 ,
         \DLX_Datapath/RegisterFile/N25766 ,
         \DLX_Datapath/RegisterFile/N25765 ,
         \DLX_Datapath/RegisterFile/N25764 ,
         \DLX_Datapath/RegisterFile/N25763 ,
         \DLX_Datapath/RegisterFile/N25762 ,
         \DLX_Datapath/RegisterFile/N25761 ,
         \DLX_Datapath/RegisterFile/N25760 ,
         \DLX_Datapath/RegisterFile/N25759 ,
         \DLX_Datapath/RegisterFile/N25758 ,
         \DLX_Datapath/RegisterFile/N25757 ,
         \DLX_Datapath/RegisterFile/N25756 ,
         \DLX_Datapath/RegisterFile/N25755 ,
         \DLX_Datapath/RegisterFile/N25754 ,
         \DLX_Datapath/RegisterFile/N25753 ,
         \DLX_Datapath/RegisterFile/N25752 ,
         \DLX_Datapath/RegisterFile/N25751 ,
         \DLX_Datapath/RegisterFile/N25750 ,
         \DLX_Datapath/RegisterFile/N25749 ,
         \DLX_Datapath/RegisterFile/N25748 ,
         \DLX_Datapath/RegisterFile/N25747 ,
         \DLX_Datapath/RegisterFile/N25746 ,
         \DLX_Datapath/RegisterFile/N25745 ,
         \DLX_Datapath/RegisterFile/N25744 ,
         \DLX_Datapath/RegisterFile/N25743 ,
         \DLX_Datapath/RegisterFile/N25742 ,
         \DLX_Datapath/RegisterFile/N25741 ,
         \DLX_Datapath/RegisterFile/N25740 ,
         \DLX_Datapath/RegisterFile/N25739 ,
         \DLX_Datapath/RegisterFile/N25738 ,
         \DLX_Datapath/RegisterFile/N25737 ,
         \DLX_Datapath/RegisterFile/N25735 ,
         \DLX_Datapath/RegisterFile/N25734 ,
         \DLX_Datapath/RegisterFile/N25733 ,
         \DLX_Datapath/RegisterFile/N25731 ,
         \DLX_Datapath/RegisterFile/N25730 ,
         \DLX_Datapath/RegisterFile/N25729 ,
         \DLX_Datapath/RegisterFile/N25728 ,
         \DLX_Datapath/RegisterFile/N25727 ,
         \DLX_Datapath/RegisterFile/N25726 ,
         \DLX_Datapath/RegisterFile/N25725 ,
         \DLX_Datapath/RegisterFile/N25724 ,
         \DLX_Datapath/RegisterFile/N25723 ,
         \DLX_Datapath/RegisterFile/N25722 ,
         \DLX_Datapath/RegisterFile/N25721 ,
         \DLX_Datapath/RegisterFile/N25720 ,
         \DLX_Datapath/RegisterFile/N25719 ,
         \DLX_Datapath/RegisterFile/N25718 ,
         \DLX_Datapath/RegisterFile/N25716 ,
         \DLX_Datapath/RegisterFile/N25715 ,
         \DLX_Datapath/RegisterFile/N25714 ,
         \DLX_Datapath/RegisterFile/N25712 ,
         \DLX_Datapath/RegisterFile/N25711 ,
         \DLX_Datapath/RegisterFile/N25710 ,
         \DLX_Datapath/RegisterFile/N25709 ,
         \DLX_Datapath/RegisterFile/N25708 ,
         \DLX_Datapath/RegisterFile/N25707 ,
         \DLX_Datapath/RegisterFile/N25706 ,
         \DLX_Datapath/RegisterFile/N25705 ,
         \DLX_Datapath/RegisterFile/N25704 ,
         \DLX_Datapath/RegisterFile/N25703 ,
         \DLX_Datapath/RegisterFile/N25702 ,
         \DLX_Datapath/RegisterFile/N25701 ,
         \DLX_Datapath/RegisterFile/N25700 ,
         \DLX_Datapath/RegisterFile/N25699 ,
         \DLX_Datapath/RegisterFile/N25698 ,
         \DLX_Datapath/RegisterFile/N25697 ,
         \DLX_Datapath/RegisterFile/N25696 ,
         \DLX_Datapath/RegisterFile/N25695 ,
         \DLX_Datapath/RegisterFile/N25694 ,
         \DLX_Datapath/RegisterFile/N25693 ,
         \DLX_Datapath/RegisterFile/N25692 ,
         \DLX_Datapath/RegisterFile/N25691 ,
         \DLX_Datapath/RegisterFile/N25690 ,
         \DLX_Datapath/RegisterFile/N25689 ,
         \DLX_Datapath/RegisterFile/N25688 ,
         \DLX_Datapath/RegisterFile/N25687 ,
         \DLX_Datapath/RegisterFile/N25686 ,
         \DLX_Datapath/RegisterFile/N25685 ,
         \DLX_Datapath/RegisterFile/N25684 ,
         \DLX_Datapath/RegisterFile/N25683 ,
         \DLX_Datapath/RegisterFile/N25682 ,
         \DLX_Datapath/RegisterFile/N25681 ,
         \DLX_Datapath/RegisterFile/N25680 ,
         \DLX_Datapath/RegisterFile/N25679 ,
         \DLX_Datapath/RegisterFile/N25678 ,
         \DLX_Datapath/RegisterFile/N25677 ,
         \DLX_Datapath/RegisterFile/N25676 ,
         \DLX_Datapath/RegisterFile/N25675 ,
         \DLX_Datapath/RegisterFile/N25671 ,
         \DLX_Datapath/RegisterFile/N25670 ,
         \DLX_Datapath/RegisterFile/N25669 ,
         \DLX_Datapath/RegisterFile/N25668 ,
         \DLX_Datapath/RegisterFile/N25667 ,
         \DLX_Datapath/RegisterFile/N25666 ,
         \DLX_Datapath/RegisterFile/N25665 ,
         \DLX_Datapath/RegisterFile/N25664 ,
         \DLX_Datapath/RegisterFile/N25663 ,
         \DLX_Datapath/RegisterFile/N25662 ,
         \DLX_Datapath/RegisterFile/N25661 ,
         \DLX_Datapath/RegisterFile/N25660 ,
         \DLX_Datapath/RegisterFile/N25659 ,
         \DLX_Datapath/RegisterFile/N25657 ,
         \DLX_Datapath/RegisterFile/N25656 ,
         \DLX_Datapath/RegisterFile/N25655 ,
         \DLX_Datapath/RegisterFile/N25654 ,
         \DLX_Datapath/RegisterFile/N25653 ,
         \DLX_Datapath/RegisterFile/N25652 ,
         \DLX_Datapath/RegisterFile/N25651 ,
         \DLX_Datapath/RegisterFile/N25650 ,
         \DLX_Datapath/RegisterFile/N25649 ,
         \DLX_Datapath/RegisterFile/N25648 ,
         \DLX_Datapath/RegisterFile/N25647 ,
         \DLX_Datapath/RegisterFile/N25646 ,
         \DLX_Datapath/RegisterFile/N25644 ,
         \DLX_Datapath/RegisterFile/N25643 ,
         \DLX_Datapath/RegisterFile/N25642 ,
         \DLX_Datapath/RegisterFile/N25641 ,
         \DLX_Datapath/RegisterFile/N25640 ,
         \DLX_Datapath/RegisterFile/N25639 ,
         \DLX_Datapath/RegisterFile/N25638 ,
         \DLX_Datapath/RegisterFile/N25637 ,
         \DLX_Datapath/RegisterFile/N25636 ,
         \DLX_Datapath/RegisterFile/N25635 ,
         \DLX_Datapath/RegisterFile/N25634 ,
         \DLX_Datapath/RegisterFile/N25633 ,
         \DLX_Datapath/RegisterFile/N25632 ,
         \DLX_Datapath/RegisterFile/N25631 ,
         \DLX_Datapath/RegisterFile/N25630 ,
         \DLX_Datapath/RegisterFile/N25629 ,
         \DLX_Datapath/RegisterFile/N25628 ,
         \DLX_Datapath/RegisterFile/N25627 ,
         \DLX_Datapath/RegisterFile/N25626 ,
         \DLX_Datapath/RegisterFile/N25625 ,
         \DLX_Datapath/RegisterFile/N25624 ,
         \DLX_Datapath/RegisterFile/N25623 ,
         \DLX_Datapath/RegisterFile/N25622 ,
         \DLX_Datapath/RegisterFile/N25621 ,
         \DLX_Datapath/RegisterFile/N25620 ,
         \DLX_Datapath/RegisterFile/N25619 ,
         \DLX_Datapath/RegisterFile/N25618 ,
         \DLX_Datapath/RegisterFile/N25617 ,
         \DLX_Datapath/RegisterFile/N25616 ,
         \DLX_Datapath/RegisterFile/N25615 ,
         \DLX_Datapath/RegisterFile/N25614 ,
         \DLX_Datapath/RegisterFile/N25613 ,
         \DLX_Datapath/RegisterFile/N25612 ,
         \DLX_Datapath/RegisterFile/N25611 ,
         \DLX_Datapath/RegisterFile/N25610 ,
         \DLX_Datapath/RegisterFile/N25609 ,
         \DLX_Datapath/RegisterFile/N25608 ,
         \DLX_Datapath/RegisterFile/N25607 ,
         \DLX_Datapath/RegisterFile/N25606 ,
         \DLX_Datapath/RegisterFile/N25605 ,
         \DLX_Datapath/RegisterFile/N25604 ,
         \DLX_Datapath/RegisterFile/N25603 ,
         \DLX_Datapath/RegisterFile/N25602 ,
         \DLX_Datapath/RegisterFile/N25601 ,
         \DLX_Datapath/RegisterFile/N25600 ,
         \DLX_Datapath/RegisterFile/N25599 ,
         \DLX_Datapath/RegisterFile/N25598 ,
         \DLX_Datapath/RegisterFile/N25597 ,
         \DLX_Datapath/RegisterFile/N25596 ,
         \DLX_Datapath/RegisterFile/N25595 ,
         \DLX_Datapath/RegisterFile/N25594 ,
         \DLX_Datapath/RegisterFile/N25593 ,
         \DLX_Datapath/RegisterFile/N25592 ,
         \DLX_Datapath/RegisterFile/N25591 ,
         \DLX_Datapath/RegisterFile/N25590 ,
         \DLX_Datapath/RegisterFile/N25589 ,
         \DLX_Datapath/RegisterFile/N25588 ,
         \DLX_Datapath/RegisterFile/N25587 ,
         \DLX_Datapath/RegisterFile/N25586 ,
         \DLX_Datapath/RegisterFile/N25585 ,
         \DLX_Datapath/RegisterFile/N25584 ,
         \DLX_Datapath/RegisterFile/N25583 ,
         \DLX_Datapath/RegisterFile/N25582 ,
         \DLX_Datapath/RegisterFile/N25581 ,
         \DLX_Datapath/RegisterFile/N25580 ,
         \DLX_Datapath/RegisterFile/N25579 ,
         \DLX_Datapath/RegisterFile/N25578 ,
         \DLX_Datapath/RegisterFile/N25577 ,
         \DLX_Datapath/RegisterFile/N25576 ,
         \DLX_Datapath/RegisterFile/N25575 ,
         \DLX_Datapath/RegisterFile/N25574 ,
         \DLX_Datapath/RegisterFile/N25573 ,
         \DLX_Datapath/RegisterFile/N25572 ,
         \DLX_Datapath/RegisterFile/N25571 ,
         \DLX_Datapath/RegisterFile/N25570 ,
         \DLX_Datapath/RegisterFile/N25569 ,
         \DLX_Datapath/RegisterFile/N25568 ,
         \DLX_Datapath/RegisterFile/N25567 ,
         \DLX_Datapath/RegisterFile/N25566 ,
         \DLX_Datapath/RegisterFile/N25565 ,
         \DLX_Datapath/RegisterFile/N25564 ,
         \DLX_Datapath/RegisterFile/N25563 ,
         \DLX_Datapath/RegisterFile/N25562 ,
         \DLX_Datapath/RegisterFile/N25561 ,
         \DLX_Datapath/RegisterFile/N25560 ,
         \DLX_Datapath/RegisterFile/N25559 ,
         \DLX_Datapath/RegisterFile/N25558 ,
         \DLX_Datapath/RegisterFile/N25557 ,
         \DLX_Datapath/RegisterFile/N25556 ,
         \DLX_Datapath/RegisterFile/N25555 ,
         \DLX_Datapath/RegisterFile/N25554 ,
         \DLX_Datapath/RegisterFile/N25553 ,
         \DLX_Datapath/RegisterFile/N25552 ,
         \DLX_Datapath/RegisterFile/N25551 ,
         \DLX_Datapath/RegisterFile/N25550 ,
         \DLX_Datapath/RegisterFile/N25549 ,
         \DLX_Datapath/RegisterFile/N25548 ,
         \DLX_Datapath/RegisterFile/N25547 ,
         \DLX_Datapath/RegisterFile/N25546 ,
         \DLX_Datapath/RegisterFile/N25545 ,
         \DLX_Datapath/RegisterFile/N25544 ,
         \DLX_Datapath/RegisterFile/N25543 ,
         \DLX_Datapath/RegisterFile/N25542 ,
         \DLX_Datapath/RegisterFile/N25541 ,
         \DLX_Datapath/RegisterFile/N25540 ,
         \DLX_Datapath/RegisterFile/N25539 ,
         \DLX_Datapath/RegisterFile/N25538 ,
         \DLX_Datapath/RegisterFile/N25537 ,
         \DLX_Datapath/RegisterFile/N25536 ,
         \DLX_Datapath/RegisterFile/N25535 ,
         \DLX_Datapath/RegisterFile/N25534 ,
         \DLX_Datapath/RegisterFile/N25533 ,
         \DLX_Datapath/RegisterFile/N25532 ,
         \DLX_Datapath/RegisterFile/N25531 ,
         \DLX_Datapath/RegisterFile/N25530 ,
         \DLX_Datapath/RegisterFile/N25529 ,
         \DLX_Datapath/RegisterFile/N25528 ,
         \DLX_Datapath/RegisterFile/N25527 ,
         \DLX_Datapath/RegisterFile/N25526 ,
         \DLX_Datapath/RegisterFile/N25525 ,
         \DLX_Datapath/RegisterFile/N25524 ,
         \DLX_Datapath/RegisterFile/N25523 ,
         \DLX_Datapath/RegisterFile/N25522 ,
         \DLX_Datapath/RegisterFile/N25521 ,
         \DLX_Datapath/RegisterFile/N25520 ,
         \DLX_Datapath/RegisterFile/N25519 ,
         \DLX_Datapath/RegisterFile/N25518 ,
         \DLX_Datapath/RegisterFile/N25517 ,
         \DLX_Datapath/RegisterFile/N25516 ,
         \DLX_Datapath/RegisterFile/N25515 ,
         \DLX_Datapath/RegisterFile/N25514 ,
         \DLX_Datapath/RegisterFile/N25513 ,
         \DLX_Datapath/RegisterFile/N25512 ,
         \DLX_Datapath/RegisterFile/N25511 ,
         \DLX_Datapath/RegisterFile/N25510 ,
         \DLX_Datapath/RegisterFile/N25509 ,
         \DLX_Datapath/RegisterFile/N25508 ,
         \DLX_Datapath/RegisterFile/N25507 ,
         \DLX_Datapath/RegisterFile/N25506 ,
         \DLX_Datapath/RegisterFile/N25505 ,
         \DLX_Datapath/RegisterFile/N25504 ,
         \DLX_Datapath/RegisterFile/N25503 ,
         \DLX_Datapath/RegisterFile/N25502 ,
         \DLX_Datapath/RegisterFile/N25501 ,
         \DLX_Datapath/RegisterFile/N25500 ,
         \DLX_Datapath/RegisterFile/N25499 ,
         \DLX_Datapath/RegisterFile/N25498 ,
         \DLX_Datapath/RegisterFile/N25497 ,
         \DLX_Datapath/RegisterFile/N25496 ,
         \DLX_Datapath/RegisterFile/N25495 ,
         \DLX_Datapath/RegisterFile/N25494 ,
         \DLX_Datapath/RegisterFile/N25493 ,
         \DLX_Datapath/RegisterFile/N25492 ,
         \DLX_Datapath/RegisterFile/N25491 ,
         \DLX_Datapath/RegisterFile/N25490 ,
         \DLX_Datapath/RegisterFile/N25489 ,
         \DLX_Datapath/RegisterFile/N25488 ,
         \DLX_Datapath/RegisterFile/N25487 ,
         \DLX_Datapath/RegisterFile/N25486 ,
         \DLX_Datapath/RegisterFile/N25485 ,
         \DLX_Datapath/RegisterFile/N25484 ,
         \DLX_Datapath/RegisterFile/N25483 ,
         \DLX_Datapath/RegisterFile/N25482 ,
         \DLX_Datapath/RegisterFile/N25481 ,
         \DLX_Datapath/RegisterFile/N25480 ,
         \DLX_Datapath/RegisterFile/N25479 ,
         \DLX_Datapath/RegisterFile/N25478 ,
         \DLX_Datapath/RegisterFile/N25477 ,
         \DLX_Datapath/RegisterFile/N25476 ,
         \DLX_Datapath/RegisterFile/N25475 ,
         \DLX_Datapath/RegisterFile/N25474 ,
         \DLX_Datapath/RegisterFile/N25473 ,
         \DLX_Datapath/RegisterFile/N25472 ,
         \DLX_Datapath/RegisterFile/N25471 ,
         \DLX_Datapath/RegisterFile/N25470 ,
         \DLX_Datapath/RegisterFile/N25469 ,
         \DLX_Datapath/RegisterFile/N25468 ,
         \DLX_Datapath/RegisterFile/N25467 ,
         \DLX_Datapath/RegisterFile/N25466 ,
         \DLX_Datapath/RegisterFile/N25465 ,
         \DLX_Datapath/RegisterFile/N25464 ,
         \DLX_Datapath/RegisterFile/N25463 ,
         \DLX_Datapath/RegisterFile/N25462 ,
         \DLX_Datapath/RegisterFile/N25461 ,
         \DLX_Datapath/RegisterFile/N25460 ,
         \DLX_Datapath/RegisterFile/N25459 ,
         \DLX_Datapath/RegisterFile/N25458 ,
         \DLX_Datapath/RegisterFile/N25457 ,
         \DLX_Datapath/RegisterFile/N25456 ,
         \DLX_Datapath/RegisterFile/N25455 ,
         \DLX_Datapath/RegisterFile/N25454 ,
         \DLX_Datapath/RegisterFile/N25453 ,
         \DLX_Datapath/RegisterFile/N25452 ,
         \DLX_Datapath/RegisterFile/N25451 ,
         \DLX_Datapath/RegisterFile/N25450 ,
         \DLX_Datapath/RegisterFile/N25449 ,
         \DLX_Datapath/RegisterFile/N25448 ,
         \DLX_Datapath/RegisterFile/N25447 ,
         \DLX_Datapath/RegisterFile/N25446 ,
         \DLX_Datapath/RegisterFile/N25445 ,
         \DLX_Datapath/RegisterFile/N25444 ,
         \DLX_Datapath/RegisterFile/N25443 ,
         \DLX_Datapath/RegisterFile/N25442 ,
         \DLX_Datapath/RegisterFile/N25441 ,
         \DLX_Datapath/RegisterFile/N25440 ,
         \DLX_Datapath/RegisterFile/N25439 ,
         \DLX_Datapath/RegisterFile/N25438 ,
         \DLX_Datapath/RegisterFile/N25437 ,
         \DLX_Datapath/RegisterFile/N25436 ,
         \DLX_Datapath/RegisterFile/N25435 ,
         \DLX_Datapath/RegisterFile/N25434 ,
         \DLX_Datapath/RegisterFile/N25433 ,
         \DLX_Datapath/RegisterFile/N25432 ,
         \DLX_Datapath/RegisterFile/N25431 ,
         \DLX_Datapath/RegisterFile/N25430 ,
         \DLX_Datapath/RegisterFile/N25429 ,
         \DLX_Datapath/RegisterFile/N25428 ,
         \DLX_Datapath/RegisterFile/N25427 ,
         \DLX_Datapath/RegisterFile/N25426 ,
         \DLX_Datapath/RegisterFile/N25425 ,
         \DLX_Datapath/RegisterFile/N25424 ,
         \DLX_Datapath/RegisterFile/N25423 ,
         \DLX_Datapath/RegisterFile/N25422 ,
         \DLX_Datapath/RegisterFile/N25421 ,
         \DLX_Datapath/RegisterFile/N25420 ,
         \DLX_Datapath/RegisterFile/N25419 ,
         \DLX_Datapath/RegisterFile/N25418 ,
         \DLX_Datapath/RegisterFile/N25417 ,
         \DLX_Datapath/RegisterFile/N25416 ,
         \DLX_Datapath/RegisterFile/N25415 ,
         \DLX_Datapath/RegisterFile/N25414 ,
         \DLX_Datapath/RegisterFile/N25413 ,
         \DLX_Datapath/RegisterFile/N25412 ,
         \DLX_Datapath/RegisterFile/N25411 ,
         \DLX_Datapath/RegisterFile/N25410 ,
         \DLX_Datapath/RegisterFile/N25409 ,
         \DLX_Datapath/RegisterFile/N25408 ,
         \DLX_Datapath/RegisterFile/N25407 ,
         \DLX_Datapath/RegisterFile/N25406 ,
         \DLX_Datapath/RegisterFile/N25405 ,
         \DLX_Datapath/RegisterFile/N25404 ,
         \DLX_Datapath/RegisterFile/N25403 ,
         \DLX_Datapath/RegisterFile/N25402 ,
         \DLX_Datapath/RegisterFile/N25401 ,
         \DLX_Datapath/RegisterFile/N25400 ,
         \DLX_Datapath/RegisterFile/N25399 ,
         \DLX_Datapath/RegisterFile/N25398 ,
         \DLX_Datapath/RegisterFile/N25397 ,
         \DLX_Datapath/RegisterFile/N25396 ,
         \DLX_Datapath/RegisterFile/N25395 ,
         \DLX_Datapath/RegisterFile/N25394 ,
         \DLX_Datapath/RegisterFile/N25393 ,
         \DLX_Datapath/RegisterFile/N25392 ,
         \DLX_Datapath/RegisterFile/N25391 ,
         \DLX_Datapath/RegisterFile/N25390 ,
         \DLX_Datapath/RegisterFile/N25389 ,
         \DLX_Datapath/RegisterFile/N25388 ,
         \DLX_Datapath/RegisterFile/N25387 ,
         \DLX_Datapath/RegisterFile/N25386 ,
         \DLX_Datapath/RegisterFile/N25385 ,
         \DLX_Datapath/RegisterFile/N25384 ,
         \DLX_Datapath/RegisterFile/N25383 ,
         \DLX_Datapath/RegisterFile/N25382 ,
         \DLX_Datapath/RegisterFile/N25381 ,
         \DLX_Datapath/RegisterFile/N25380 ,
         \DLX_Datapath/RegisterFile/N25379 ,
         \DLX_Datapath/RegisterFile/N25378 ,
         \DLX_Datapath/RegisterFile/N25377 ,
         \DLX_Datapath/RegisterFile/N25376 ,
         \DLX_Datapath/RegisterFile/N25375 ,
         \DLX_Datapath/RegisterFile/N25374 ,
         \DLX_Datapath/RegisterFile/N25373 ,
         \DLX_Datapath/RegisterFile/N25372 ,
         \DLX_Datapath/RegisterFile/N25371 ,
         \DLX_Datapath/RegisterFile/N25370 ,
         \DLX_Datapath/RegisterFile/N25369 ,
         \DLX_Datapath/RegisterFile/N25368 ,
         \DLX_Datapath/RegisterFile/N25367 ,
         \DLX_Datapath/RegisterFile/N25366 ,
         \DLX_Datapath/RegisterFile/N25365 ,
         \DLX_Datapath/RegisterFile/N25364 ,
         \DLX_Datapath/RegisterFile/N25363 ,
         \DLX_Datapath/RegisterFile/N25362 ,
         \DLX_Datapath/RegisterFile/N25361 ,
         \DLX_Datapath/RegisterFile/N25360 ,
         \DLX_Datapath/RegisterFile/N25359 ,
         \DLX_Datapath/RegisterFile/N25358 ,
         \DLX_Datapath/RegisterFile/N25357 ,
         \DLX_Datapath/RegisterFile/N25356 ,
         \DLX_Datapath/RegisterFile/N25355 ,
         \DLX_Datapath/RegisterFile/N25353 ,
         \DLX_Datapath/RegisterFile/N25349 ,
         \DLX_Datapath/RegisterFile/N25348 ,
         \DLX_Datapath/RegisterFile/N25347 ,
         \DLX_Datapath/RegisterFile/N25346 ,
         \DLX_Datapath/RegisterFile/N25344 ,
         \DLX_Datapath/RegisterFile/N25341 ,
         \DLX_Datapath/RegisterFile/N25340 ,
         \DLX_Datapath/RegisterFile/N25339 ,
         \DLX_Datapath/RegisterFile/N25337 ,
         \DLX_Datapath/RegisterFile/N25335 ,
         \DLX_Datapath/RegisterFile/N25334 ,
         \DLX_Datapath/RegisterFile/N25330 ,
         \DLX_Datapath/RegisterFile/N25328 ,
         \DLX_Datapath/RegisterFile/N25327 ,
         \DLX_Datapath/RegisterFile/N25326 ,
         \DLX_Datapath/RegisterFile/N25325 ,
         \DLX_Datapath/RegisterFile/N25323 ,
         \DLX_Datapath/RegisterFile/N25322 ,
         \DLX_Datapath/RegisterFile/N25321 ,
         \DLX_Datapath/RegisterFile/N25320 ,
         \DLX_Datapath/RegisterFile/N25319 ,
         \DLX_Datapath/RegisterFile/N25318 ,
         \DLX_Datapath/RegisterFile/N25317 ,
         \DLX_Datapath/RegisterFile/N25316 ,
         \DLX_Datapath/RegisterFile/N25315 ,
         \DLX_Datapath/RegisterFile/N25314 ,
         \DLX_Datapath/RegisterFile/N25313 ,
         \DLX_Datapath/RegisterFile/N25312 ,
         \DLX_Datapath/RegisterFile/N25311 ,
         \DLX_Datapath/RegisterFile/N25310 ,
         \DLX_Datapath/RegisterFile/N25309 ,
         \DLX_Datapath/RegisterFile/N25308 ,
         \DLX_Datapath/RegisterFile/N25307 ,
         \DLX_Datapath/RegisterFile/N25306 ,
         \DLX_Datapath/RegisterFile/N25305 ,
         \DLX_Datapath/RegisterFile/N25304 ,
         \DLX_Datapath/RegisterFile/N25303 ,
         \DLX_Datapath/RegisterFile/N25302 ,
         \DLX_Datapath/RegisterFile/N25301 ,
         \DLX_Datapath/RegisterFile/N25300 ,
         \DLX_Datapath/RegisterFile/N25299 ,
         \DLX_Datapath/RegisterFile/N25298 ,
         \DLX_Datapath/RegisterFile/N25297 ,
         \DLX_Datapath/RegisterFile/N25296 ,
         \DLX_Datapath/RegisterFile/N25295 ,
         \DLX_Datapath/RegisterFile/N25294 ,
         \DLX_Datapath/RegisterFile/N25293 ,
         \DLX_Datapath/RegisterFile/N25292 ,
         \DLX_Datapath/RegisterFile/N25291 ,
         \DLX_Datapath/RegisterFile/N25290 ,
         \DLX_Datapath/RegisterFile/N25289 ,
         \DLX_Datapath/RegisterFile/N25288 ,
         \DLX_Datapath/RegisterFile/N25287 ,
         \DLX_Datapath/RegisterFile/N25286 ,
         \DLX_Datapath/RegisterFile/N25285 ,
         \DLX_Datapath/RegisterFile/N25284 ,
         \DLX_Datapath/RegisterFile/N25283 ,
         \DLX_Datapath/RegisterFile/N25282 ,
         \DLX_Datapath/RegisterFile/N25281 ,
         \DLX_Datapath/RegisterFile/N25280 ,
         \DLX_Datapath/RegisterFile/N25279 ,
         \DLX_Datapath/RegisterFile/N25278 ,
         \DLX_Datapath/RegisterFile/N25277 ,
         \DLX_Datapath/RegisterFile/N25276 ,
         \DLX_Datapath/RegisterFile/N25275 ,
         \DLX_Datapath/RegisterFile/N25274 ,
         \DLX_Datapath/RegisterFile/N25273 ,
         \DLX_Datapath/RegisterFile/N25272 ,
         \DLX_Datapath/RegisterFile/N25271 ,
         \DLX_Datapath/RegisterFile/N25270 ,
         \DLX_Datapath/RegisterFile/N25269 ,
         \DLX_Datapath/RegisterFile/N25268 ,
         \DLX_Datapath/RegisterFile/N25267 ,
         \DLX_Datapath/RegisterFile/N25266 ,
         \DLX_Datapath/RegisterFile/N25265 ,
         \DLX_Datapath/RegisterFile/N25264 ,
         \DLX_Datapath/RegisterFile/N25263 ,
         \DLX_Datapath/RegisterFile/N25262 ,
         \DLX_Datapath/RegisterFile/N25261 ,
         \DLX_Datapath/RegisterFile/N25260 ,
         \DLX_Datapath/RegisterFile/N25259 ,
         \DLX_Datapath/RegisterFile/N25258 ,
         \DLX_Datapath/RegisterFile/N25257 ,
         \DLX_Datapath/RegisterFile/N25256 ,
         \DLX_Datapath/RegisterFile/N25255 ,
         \DLX_Datapath/RegisterFile/N25254 ,
         \DLX_Datapath/RegisterFile/N25253 ,
         \DLX_Datapath/RegisterFile/N25252 ,
         \DLX_Datapath/RegisterFile/N25251 ,
         \DLX_Datapath/RegisterFile/N25250 ,
         \DLX_Datapath/RegisterFile/N25249 ,
         \DLX_Datapath/RegisterFile/N25248 ,
         \DLX_Datapath/RegisterFile/N25247 ,
         \DLX_Datapath/RegisterFile/N25246 ,
         \DLX_Datapath/RegisterFile/N25245 ,
         \DLX_Datapath/RegisterFile/N25244 ,
         \DLX_Datapath/RegisterFile/N25243 ,
         \DLX_Datapath/RegisterFile/N25242 ,
         \DLX_Datapath/RegisterFile/N25241 ,
         \DLX_Datapath/RegisterFile/N25240 ,
         \DLX_Datapath/RegisterFile/N25239 ,
         \DLX_Datapath/RegisterFile/N25238 ,
         \DLX_Datapath/RegisterFile/N25237 ,
         \DLX_Datapath/RegisterFile/N25236 ,
         \DLX_Datapath/RegisterFile/N25235 ,
         \DLX_Datapath/RegisterFile/N25234 ,
         \DLX_Datapath/RegisterFile/N25233 ,
         \DLX_Datapath/RegisterFile/N25232 ,
         \DLX_Datapath/RegisterFile/N25231 ,
         \DLX_Datapath/RegisterFile/N25230 ,
         \DLX_Datapath/RegisterFile/N25229 ,
         \DLX_Datapath/RegisterFile/N25228 ,
         \DLX_Datapath/RegisterFile/N25227 ,
         \DLX_Datapath/RegisterFile/N25226 ,
         \DLX_Datapath/RegisterFile/N25225 ,
         \DLX_Datapath/RegisterFile/N25224 ,
         \DLX_Datapath/RegisterFile/N25223 ,
         \DLX_Datapath/RegisterFile/N25222 ,
         \DLX_Datapath/RegisterFile/N25221 ,
         \DLX_Datapath/RegisterFile/N25220 ,
         \DLX_Datapath/RegisterFile/N25219 ,
         \DLX_Datapath/RegisterFile/N25218 ,
         \DLX_Datapath/RegisterFile/N25217 ,
         \DLX_Datapath/RegisterFile/N25216 ,
         \DLX_Datapath/RegisterFile/N25215 ,
         \DLX_Datapath/RegisterFile/N25214 ,
         \DLX_Datapath/RegisterFile/N25213 ,
         \DLX_Datapath/RegisterFile/N25212 ,
         \DLX_Datapath/RegisterFile/N25211 ,
         \DLX_Datapath/RegisterFile/N25210 ,
         \DLX_Datapath/RegisterFile/N25209 ,
         \DLX_Datapath/RegisterFile/N25208 ,
         \DLX_Datapath/RegisterFile/N25207 ,
         \DLX_Datapath/RegisterFile/N25206 ,
         \DLX_Datapath/RegisterFile/N25205 ,
         \DLX_Datapath/RegisterFile/N25204 ,
         \DLX_Datapath/RegisterFile/N25203 ,
         \DLX_Datapath/RegisterFile/N25202 ,
         \DLX_Datapath/RegisterFile/N25201 ,
         \DLX_Datapath/RegisterFile/N25200 ,
         \DLX_Datapath/RegisterFile/N25199 ,
         \DLX_Datapath/RegisterFile/N25198 ,
         \DLX_Datapath/RegisterFile/N25197 ,
         \DLX_Datapath/RegisterFile/N25196 ,
         \DLX_Datapath/RegisterFile/N25195 ,
         \DLX_Datapath/RegisterFile/N25194 ,
         \DLX_Datapath/RegisterFile/N25193 ,
         \DLX_Datapath/RegisterFile/N25192 ,
         \DLX_Datapath/RegisterFile/N25191 ,
         \DLX_Datapath/RegisterFile/N25190 ,
         \DLX_Datapath/RegisterFile/N25189 ,
         \DLX_Datapath/RegisterFile/N25188 ,
         \DLX_Datapath/RegisterFile/N25187 ,
         \DLX_Datapath/RegisterFile/N25186 ,
         \DLX_Datapath/RegisterFile/N25185 ,
         \DLX_Datapath/RegisterFile/N25184 ,
         \DLX_Datapath/RegisterFile/N25183 ,
         \DLX_Datapath/RegisterFile/N25182 ,
         \DLX_Datapath/RegisterFile/N25181 ,
         \DLX_Datapath/RegisterFile/N25180 ,
         \DLX_Datapath/RegisterFile/N25179 ,
         \DLX_Datapath/RegisterFile/N25178 ,
         \DLX_Datapath/RegisterFile/N25177 ,
         \DLX_Datapath/RegisterFile/N25176 ,
         \DLX_Datapath/RegisterFile/N25175 ,
         \DLX_Datapath/RegisterFile/N25174 ,
         \DLX_Datapath/RegisterFile/N25173 ,
         \DLX_Datapath/RegisterFile/N25172 ,
         \DLX_Datapath/RegisterFile/N25171 ,
         \DLX_Datapath/RegisterFile/N25170 ,
         \DLX_Datapath/RegisterFile/N25169 ,
         \DLX_Datapath/RegisterFile/N25168 ,
         \DLX_Datapath/RegisterFile/N25167 ,
         \DLX_Datapath/RegisterFile/N25166 ,
         \DLX_Datapath/RegisterFile/N25165 ,
         \DLX_Datapath/RegisterFile/N25164 ,
         \DLX_Datapath/RegisterFile/N25163 ,
         \DLX_Datapath/RegisterFile/N25162 ,
         \DLX_Datapath/RegisterFile/N25161 ,
         \DLX_Datapath/RegisterFile/N25160 ,
         \DLX_Datapath/RegisterFile/N25159 ,
         \DLX_Datapath/RegisterFile/N25158 ,
         \DLX_Datapath/RegisterFile/N25157 ,
         \DLX_Datapath/RegisterFile/N25156 ,
         \DLX_Datapath/RegisterFile/N25155 ,
         \DLX_Datapath/RegisterFile/N25154 ,
         \DLX_Datapath/RegisterFile/N25153 ,
         \DLX_Datapath/RegisterFile/N25152 ,
         \DLX_Datapath/RegisterFile/N25151 ,
         \DLX_Datapath/RegisterFile/N25148 ,
         \DLX_Datapath/RegisterFile/N25147 ,
         \DLX_Datapath/RegisterFile/N25144 ,
         \DLX_Datapath/RegisterFile/N25143 ,
         \DLX_Datapath/RegisterFile/N25142 ,
         \DLX_Datapath/RegisterFile/N25139 ,
         \DLX_Datapath/RegisterFile/N25138 ,
         \DLX_Datapath/RegisterFile/N25137 ,
         \DLX_Datapath/RegisterFile/N25136 ,
         \DLX_Datapath/RegisterFile/N25135 ,
         \DLX_Datapath/RegisterFile/N25134 ,
         \DLX_Datapath/RegisterFile/N25133 ,
         \DLX_Datapath/RegisterFile/N25132 ,
         \DLX_Datapath/RegisterFile/N25131 ,
         \DLX_Datapath/RegisterFile/N25130 ,
         \DLX_Datapath/RegisterFile/N25129 ,
         \DLX_Datapath/RegisterFile/N25128 ,
         \DLX_Datapath/RegisterFile/N25127 ,
         \DLX_Datapath/RegisterFile/N25126 ,
         \DLX_Datapath/RegisterFile/N25125 ,
         \DLX_Datapath/RegisterFile/N25124 ,
         \DLX_Datapath/RegisterFile/N25123 ,
         \DLX_Datapath/RegisterFile/N25122 ,
         \DLX_Datapath/RegisterFile/N25121 ,
         \DLX_Datapath/RegisterFile/N25120 ,
         \DLX_Datapath/RegisterFile/N25119 ,
         \DLX_Datapath/RegisterFile/N25118 ,
         \DLX_Datapath/RegisterFile/N25117 ,
         \DLX_Datapath/RegisterFile/N25116 ,
         \DLX_Datapath/RegisterFile/N25115 ,
         \DLX_Datapath/RegisterFile/N25114 ,
         \DLX_Datapath/RegisterFile/N25113 ,
         \DLX_Datapath/RegisterFile/N25112 ,
         \DLX_Datapath/RegisterFile/N25111 ,
         \DLX_Datapath/RegisterFile/N25110 ,
         \DLX_Datapath/RegisterFile/N25109 ,
         \DLX_Datapath/RegisterFile/N25108 ,
         \DLX_Datapath/RegisterFile/N25107 ,
         \DLX_Datapath/RegisterFile/N25106 ,
         \DLX_Datapath/RegisterFile/N25105 ,
         \DLX_Datapath/RegisterFile/N25104 ,
         \DLX_Datapath/RegisterFile/N25103 ,
         \DLX_Datapath/RegisterFile/N25102 ,
         \DLX_Datapath/RegisterFile/N25101 ,
         \DLX_Datapath/RegisterFile/N25100 ,
         \DLX_Datapath/RegisterFile/N25099 ,
         \DLX_Datapath/RegisterFile/N25097 ,
         \DLX_Datapath/RegisterFile/N25094 ,
         \DLX_Datapath/RegisterFile/N25093 ,
         \DLX_Datapath/RegisterFile/N25092 ,
         \DLX_Datapath/RegisterFile/N25091 ,
         \DLX_Datapath/RegisterFile/N25090 ,
         \DLX_Datapath/RegisterFile/N25089 ,
         \DLX_Datapath/RegisterFile/N25088 ,
         \DLX_Datapath/RegisterFile/N25087 ,
         \DLX_Datapath/RegisterFile/N25086 ,
         \DLX_Datapath/RegisterFile/N25085 ,
         \DLX_Datapath/RegisterFile/N25084 ,
         \DLX_Datapath/RegisterFile/N25083 ,
         \DLX_Datapath/RegisterFile/N25081 ,
         \DLX_Datapath/RegisterFile/N25079 ,
         \DLX_Datapath/RegisterFile/N25078 ,
         \DLX_Datapath/RegisterFile/N25076 ,
         \DLX_Datapath/RegisterFile/N25074 ,
         \DLX_Datapath/RegisterFile/N25072 ,
         \DLX_Datapath/RegisterFile/N25071 ,
         \DLX_Datapath/RegisterFile/N25070 ,
         \DLX_Datapath/RegisterFile/N25069 ,
         \DLX_Datapath/RegisterFile/N25067 ,
         \DLX_Datapath/RegisterFile/N25066 ,
         \DLX_Datapath/RegisterFile/N25065 ,
         \DLX_Datapath/RegisterFile/N25064 ,
         \DLX_Datapath/RegisterFile/N25063 ,
         \DLX_Datapath/RegisterFile/N25062 ,
         \DLX_Datapath/RegisterFile/N25061 ,
         \DLX_Datapath/RegisterFile/N25060 ,
         \DLX_Datapath/RegisterFile/N25059 ,
         \DLX_Datapath/RegisterFile/N25058 ,
         \DLX_Datapath/RegisterFile/N25057 ,
         \DLX_Datapath/RegisterFile/N25056 ,
         \DLX_Datapath/RegisterFile/N25055 ,
         \DLX_Datapath/RegisterFile/N25054 ,
         \DLX_Datapath/RegisterFile/N25053 ,
         \DLX_Datapath/RegisterFile/N25052 ,
         \DLX_Datapath/RegisterFile/N25051 ,
         \DLX_Datapath/RegisterFile/N25050 ,
         \DLX_Datapath/RegisterFile/N25049 ,
         \DLX_Datapath/RegisterFile/N25048 ,
         \DLX_Datapath/RegisterFile/N25047 ,
         \DLX_Datapath/RegisterFile/N25046 ,
         \DLX_Datapath/RegisterFile/N25045 ,
         \DLX_Datapath/RegisterFile/N25044 ,
         \DLX_Datapath/RegisterFile/N25043 ,
         \DLX_Datapath/RegisterFile/N25042 ,
         \DLX_Datapath/RegisterFile/N25041 ,
         \DLX_Datapath/RegisterFile/N25040 ,
         \DLX_Datapath/RegisterFile/N25039 ,
         \DLX_Datapath/RegisterFile/N25038 ,
         \DLX_Datapath/RegisterFile/N25037 ,
         \DLX_Datapath/RegisterFile/N25036 ,
         \DLX_Datapath/RegisterFile/N25035 ,
         \DLX_Datapath/RegisterFile/N25033 ,
         \DLX_Datapath/RegisterFile/N25030 ,
         \DLX_Datapath/RegisterFile/N25029 ,
         \DLX_Datapath/RegisterFile/N25028 ,
         \DLX_Datapath/RegisterFile/N25027 ,
         \DLX_Datapath/RegisterFile/N25026 ,
         \DLX_Datapath/RegisterFile/N25025 ,
         \DLX_Datapath/RegisterFile/N25024 ,
         \DLX_Datapath/RegisterFile/N25023 ,
         \DLX_Datapath/RegisterFile/N25022 ,
         \DLX_Datapath/RegisterFile/N25021 ,
         \DLX_Datapath/RegisterFile/N25020 ,
         \DLX_Datapath/RegisterFile/N25019 ,
         \DLX_Datapath/RegisterFile/N25015 ,
         \DLX_Datapath/RegisterFile/N25014 ,
         \DLX_Datapath/RegisterFile/N25012 ,
         \DLX_Datapath/RegisterFile/N25011 ,
         \DLX_Datapath/RegisterFile/N25010 ,
         \DLX_Datapath/RegisterFile/N25009 ,
         \DLX_Datapath/RegisterFile/N25008 ,
         \DLX_Datapath/RegisterFile/N25007 ,
         \DLX_Datapath/RegisterFile/N25003 ,
         \DLX_Datapath/RegisterFile/N25002 ,
         \DLX_Datapath/RegisterFile/N25001 ,
         \DLX_Datapath/RegisterFile/N25000 ,
         \DLX_Datapath/RegisterFile/N24999 ,
         \DLX_Datapath/RegisterFile/N24998 ,
         \DLX_Datapath/RegisterFile/N24997 ,
         \DLX_Datapath/RegisterFile/N24996 ,
         \DLX_Datapath/RegisterFile/N24995 ,
         \DLX_Datapath/RegisterFile/N24994 ,
         \DLX_Datapath/RegisterFile/N24993 ,
         \DLX_Datapath/RegisterFile/N24992 ,
         \DLX_Datapath/RegisterFile/N24991 ,
         \DLX_Datapath/RegisterFile/N24990 ,
         \DLX_Datapath/RegisterFile/N24989 ,
         \DLX_Datapath/RegisterFile/N24988 ,
         \DLX_Datapath/RegisterFile/N24987 ,
         \DLX_Datapath/RegisterFile/N24986 ,
         \DLX_Datapath/RegisterFile/N24985 ,
         \DLX_Datapath/RegisterFile/N24984 ,
         \DLX_Datapath/RegisterFile/N24983 ,
         \DLX_Datapath/RegisterFile/N24982 ,
         \DLX_Datapath/RegisterFile/N24981 ,
         \DLX_Datapath/RegisterFile/N24980 ,
         \DLX_Datapath/RegisterFile/N24979 ,
         \DLX_Datapath/RegisterFile/N24978 ,
         \DLX_Datapath/RegisterFile/N24977 ,
         \DLX_Datapath/RegisterFile/N24976 ,
         \DLX_Datapath/RegisterFile/N24975 ,
         \DLX_Datapath/RegisterFile/N24974 ,
         \DLX_Datapath/RegisterFile/N24973 ,
         \DLX_Datapath/RegisterFile/N24972 ,
         \DLX_Datapath/RegisterFile/N24971 ,
         \DLX_Datapath/RegisterFile/N24969 ,
         \DLX_Datapath/RegisterFile/N24968 ,
         \DLX_Datapath/RegisterFile/N24966 ,
         \DLX_Datapath/RegisterFile/N24965 ,
         \DLX_Datapath/RegisterFile/N24963 ,
         \DLX_Datapath/RegisterFile/N24962 ,
         \DLX_Datapath/RegisterFile/N24961 ,
         \DLX_Datapath/RegisterFile/N24960 ,
         \DLX_Datapath/RegisterFile/N24959 ,
         \DLX_Datapath/RegisterFile/N24958 ,
         \DLX_Datapath/RegisterFile/N24957 ,
         \DLX_Datapath/RegisterFile/N24956 ,
         \DLX_Datapath/RegisterFile/N24955 ,
         \DLX_Datapath/RegisterFile/N24953 ,
         \DLX_Datapath/RegisterFile/N24951 ,
         \DLX_Datapath/RegisterFile/N24950 ,
         \DLX_Datapath/RegisterFile/N24948 ,
         \DLX_Datapath/RegisterFile/N24946 ,
         \DLX_Datapath/RegisterFile/N24944 ,
         \DLX_Datapath/RegisterFile/N24943 ,
         \DLX_Datapath/RegisterFile/N24942 ,
         \DLX_Datapath/RegisterFile/N24941 ,
         \DLX_Datapath/RegisterFile/N24939 ,
         \DLX_Datapath/RegisterFile/N24938 ,
         \DLX_Datapath/RegisterFile/N24937 ,
         \DLX_Datapath/RegisterFile/N24936 ,
         \DLX_Datapath/RegisterFile/N24935 ,
         \DLX_Datapath/RegisterFile/N24934 ,
         \DLX_Datapath/RegisterFile/N24933 ,
         \DLX_Datapath/RegisterFile/N24932 ,
         \DLX_Datapath/RegisterFile/N24931 ,
         \DLX_Datapath/RegisterFile/N24930 ,
         \DLX_Datapath/RegisterFile/N24929 ,
         \DLX_Datapath/RegisterFile/N24928 ,
         \DLX_Datapath/RegisterFile/N24927 ,
         \DLX_Datapath/RegisterFile/N24926 ,
         \DLX_Datapath/RegisterFile/N24925 ,
         \DLX_Datapath/RegisterFile/N24924 ,
         \DLX_Datapath/RegisterFile/N24923 ,
         \DLX_Datapath/RegisterFile/N24922 ,
         \DLX_Datapath/RegisterFile/N24921 ,
         \DLX_Datapath/RegisterFile/N24920 ,
         \DLX_Datapath/RegisterFile/N24919 ,
         \DLX_Datapath/RegisterFile/N24918 ,
         \DLX_Datapath/RegisterFile/N24917 ,
         \DLX_Datapath/RegisterFile/N24916 ,
         \DLX_Datapath/RegisterFile/N24915 ,
         \DLX_Datapath/RegisterFile/N24914 ,
         \DLX_Datapath/RegisterFile/N24913 ,
         \DLX_Datapath/RegisterFile/N24912 ,
         \DLX_Datapath/RegisterFile/N24911 ,
         \DLX_Datapath/RegisterFile/N24910 ,
         \DLX_Datapath/RegisterFile/N24909 ,
         \DLX_Datapath/RegisterFile/N24908 ,
         \DLX_Datapath/RegisterFile/N24907 ,
         \DLX_Datapath/RegisterFile/N24906 ,
         \DLX_Datapath/RegisterFile/N24905 ,
         \DLX_Datapath/RegisterFile/N24904 ,
         \DLX_Datapath/RegisterFile/N24903 ,
         \DLX_Datapath/RegisterFile/N24902 ,
         \DLX_Datapath/RegisterFile/N24901 ,
         \DLX_Datapath/RegisterFile/N24900 ,
         \DLX_Datapath/RegisterFile/N24898 ,
         \DLX_Datapath/RegisterFile/N24897 ,
         \DLX_Datapath/RegisterFile/N24896 ,
         \DLX_Datapath/RegisterFile/N24895 ,
         \DLX_Datapath/RegisterFile/N24894 ,
         \DLX_Datapath/RegisterFile/N24893 ,
         \DLX_Datapath/RegisterFile/N24892 ,
         \DLX_Datapath/RegisterFile/N24891 ,
         \DLX_Datapath/RegisterFile/N24890 ,
         \DLX_Datapath/RegisterFile/N24889 ,
         \DLX_Datapath/RegisterFile/N24888 ,
         \DLX_Datapath/RegisterFile/N24887 ,
         \DLX_Datapath/RegisterFile/N24886 ,
         \DLX_Datapath/RegisterFile/N24885 ,
         \DLX_Datapath/RegisterFile/N24884 ,
         \DLX_Datapath/RegisterFile/N24883 ,
         \DLX_Datapath/RegisterFile/N24882 ,
         \DLX_Datapath/RegisterFile/N24881 ,
         \DLX_Datapath/RegisterFile/N24880 ,
         \DLX_Datapath/RegisterFile/N24879 ,
         \DLX_Datapath/RegisterFile/N24878 ,
         \DLX_Datapath/RegisterFile/N24877 ,
         \DLX_Datapath/RegisterFile/N24876 ,
         \DLX_Datapath/RegisterFile/N24875 ,
         \DLX_Datapath/RegisterFile/N24874 ,
         \DLX_Datapath/RegisterFile/N24873 ,
         \DLX_Datapath/RegisterFile/N24872 ,
         \DLX_Datapath/RegisterFile/N24871 ,
         \DLX_Datapath/RegisterFile/N24870 ,
         \DLX_Datapath/RegisterFile/N24869 ,
         \DLX_Datapath/RegisterFile/N24868 ,
         \DLX_Datapath/RegisterFile/N24867 ,
         \DLX_Datapath/RegisterFile/N24866 ,
         \DLX_Datapath/RegisterFile/N24865 ,
         \DLX_Datapath/RegisterFile/N24864 ,
         \DLX_Datapath/RegisterFile/N24863 ,
         \DLX_Datapath/RegisterFile/N24862 ,
         \DLX_Datapath/RegisterFile/N24861 ,
         \DLX_Datapath/RegisterFile/N24860 ,
         \DLX_Datapath/RegisterFile/N24859 ,
         \DLX_Datapath/RegisterFile/N24858 ,
         \DLX_Datapath/RegisterFile/N24857 ,
         \DLX_Datapath/RegisterFile/N24856 ,
         \DLX_Datapath/RegisterFile/N24855 ,
         \DLX_Datapath/RegisterFile/N24854 ,
         \DLX_Datapath/RegisterFile/N24853 ,
         \DLX_Datapath/RegisterFile/N24852 ,
         \DLX_Datapath/RegisterFile/N24851 ,
         \DLX_Datapath/RegisterFile/N24850 ,
         \DLX_Datapath/RegisterFile/N24849 ,
         \DLX_Datapath/RegisterFile/N24848 ,
         \DLX_Datapath/RegisterFile/N24847 ,
         \DLX_Datapath/RegisterFile/N24846 ,
         \DLX_Datapath/RegisterFile/N24845 ,
         \DLX_Datapath/RegisterFile/N24844 ,
         \DLX_Datapath/RegisterFile/N24843 ,
         \DLX_Datapath/RegisterFile/N24842 ,
         \DLX_Datapath/RegisterFile/N24841 ,
         \DLX_Datapath/RegisterFile/N24840 ,
         \DLX_Datapath/RegisterFile/N24838 ,
         \DLX_Datapath/RegisterFile/N24837 ,
         \DLX_Datapath/RegisterFile/N24836 ,
         \DLX_Datapath/RegisterFile/N24835 ,
         \DLX_Datapath/RegisterFile/N24834 ,
         \DLX_Datapath/RegisterFile/N24833 ,
         \DLX_Datapath/RegisterFile/N24832 ,
         \DLX_Datapath/RegisterFile/N24829 ,
         \DLX_Datapath/RegisterFile/N24828 ,
         \DLX_Datapath/RegisterFile/N24827 ,
         \DLX_Datapath/RegisterFile/N24825 ,
         \DLX_Datapath/RegisterFile/N24823 ,
         \DLX_Datapath/RegisterFile/N24822 ,
         \DLX_Datapath/RegisterFile/N24820 ,
         \DLX_Datapath/RegisterFile/N24819 ,
         \DLX_Datapath/RegisterFile/N24818 ,
         \DLX_Datapath/RegisterFile/N24816 ,
         \DLX_Datapath/RegisterFile/N24815 ,
         \DLX_Datapath/RegisterFile/N24814 ,
         \DLX_Datapath/RegisterFile/N24813 ,
         \DLX_Datapath/RegisterFile/N24812 ,
         \DLX_Datapath/RegisterFile/N24811 ,
         \DLX_Datapath/RegisterFile/N24810 ,
         \DLX_Datapath/RegisterFile/N24809 ,
         \DLX_Datapath/RegisterFile/N24808 ,
         \DLX_Datapath/RegisterFile/N24807 ,
         \DLX_Datapath/RegisterFile/N24806 ,
         \DLX_Datapath/RegisterFile/N24805 ,
         \DLX_Datapath/RegisterFile/N24804 ,
         \DLX_Datapath/RegisterFile/N24803 ,
         \DLX_Datapath/RegisterFile/N24802 ,
         \DLX_Datapath/RegisterFile/N24801 ,
         \DLX_Datapath/RegisterFile/N24800 ,
         \DLX_Datapath/RegisterFile/N24799 ,
         \DLX_Datapath/RegisterFile/N24798 ,
         \DLX_Datapath/RegisterFile/N24797 ,
         \DLX_Datapath/RegisterFile/N24796 ,
         \DLX_Datapath/RegisterFile/N24795 ,
         \DLX_Datapath/RegisterFile/N24794 ,
         \DLX_Datapath/RegisterFile/N24793 ,
         \DLX_Datapath/RegisterFile/N24792 ,
         \DLX_Datapath/RegisterFile/N24791 ,
         \DLX_Datapath/RegisterFile/N24790 ,
         \DLX_Datapath/RegisterFile/N24789 ,
         \DLX_Datapath/RegisterFile/N24788 ,
         \DLX_Datapath/RegisterFile/N24787 ,
         \DLX_Datapath/RegisterFile/N24786 ,
         \DLX_Datapath/RegisterFile/N24785 ,
         \DLX_Datapath/RegisterFile/N24784 ,
         \DLX_Datapath/RegisterFile/N24783 ,
         \DLX_Datapath/RegisterFile/N24782 ,
         \DLX_Datapath/RegisterFile/N24781 ,
         \DLX_Datapath/RegisterFile/N24780 ,
         \DLX_Datapath/RegisterFile/N24779 ,
         \DLX_Datapath/RegisterFile/N24778 ,
         \DLX_Datapath/RegisterFile/N24777 ,
         \DLX_Datapath/RegisterFile/N24776 ,
         \DLX_Datapath/RegisterFile/N24774 ,
         \DLX_Datapath/RegisterFile/N24773 ,
         \DLX_Datapath/RegisterFile/N24772 ,
         \DLX_Datapath/RegisterFile/N24771 ,
         \DLX_Datapath/RegisterFile/N24770 ,
         \DLX_Datapath/RegisterFile/N24769 ,
         \DLX_Datapath/RegisterFile/N24768 ,
         \DLX_Datapath/RegisterFile/N24767 ,
         \DLX_Datapath/RegisterFile/N24765 ,
         \DLX_Datapath/RegisterFile/N24764 ,
         \DLX_Datapath/RegisterFile/N24763 ,
         \DLX_Datapath/RegisterFile/N24759 ,
         \DLX_Datapath/RegisterFile/N24758 ,
         \DLX_Datapath/RegisterFile/N24754 ,
         \DLX_Datapath/RegisterFile/N24753 ,
         \DLX_Datapath/RegisterFile/N24752 ,
         \DLX_Datapath/RegisterFile/N24751 ,
         \DLX_Datapath/RegisterFile/N24749 ,
         \DLX_Datapath/RegisterFile/N24747 ,
         \DLX_Datapath/RegisterFile/N24746 ,
         \DLX_Datapath/RegisterFile/N24745 ,
         \DLX_Datapath/RegisterFile/N24744 ,
         \DLX_Datapath/RegisterFile/N24743 ,
         \DLX_Datapath/RegisterFile/N24742 ,
         \DLX_Datapath/RegisterFile/N24741 ,
         \DLX_Datapath/RegisterFile/N24740 ,
         \DLX_Datapath/RegisterFile/N24739 ,
         \DLX_Datapath/RegisterFile/N24738 ,
         \DLX_Datapath/RegisterFile/N24737 ,
         \DLX_Datapath/RegisterFile/N24736 ,
         \DLX_Datapath/RegisterFile/N24735 ,
         \DLX_Datapath/RegisterFile/N24734 ,
         \DLX_Datapath/RegisterFile/N24733 ,
         \DLX_Datapath/RegisterFile/N24732 ,
         \DLX_Datapath/RegisterFile/N24731 ,
         \DLX_Datapath/RegisterFile/N24730 ,
         \DLX_Datapath/RegisterFile/N24729 ,
         \DLX_Datapath/RegisterFile/N24728 ,
         \DLX_Datapath/RegisterFile/N24727 ,
         \DLX_Datapath/RegisterFile/N24726 ,
         \DLX_Datapath/RegisterFile/N24725 ,
         \DLX_Datapath/RegisterFile/N24724 ,
         \DLX_Datapath/RegisterFile/N24723 ,
         \DLX_Datapath/RegisterFile/N24722 ,
         \DLX_Datapath/RegisterFile/N24721 ,
         \DLX_Datapath/RegisterFile/N24720 ,
         \DLX_Datapath/RegisterFile/N24719 ,
         \DLX_Datapath/RegisterFile/N24718 ,
         \DLX_Datapath/RegisterFile/N24717 ,
         \DLX_Datapath/RegisterFile/N24716 ,
         \DLX_Datapath/RegisterFile/N24715 ,
         \DLX_Datapath/RegisterFile/N24713 ,
         \DLX_Datapath/RegisterFile/N24712 ,
         \DLX_Datapath/RegisterFile/N24709 ,
         \DLX_Datapath/RegisterFile/N24707 ,
         \DLX_Datapath/RegisterFile/N24706 ,
         \DLX_Datapath/RegisterFile/N24704 ,
         \DLX_Datapath/RegisterFile/N24701 ,
         \DLX_Datapath/RegisterFile/N24700 ,
         \DLX_Datapath/RegisterFile/N24699 ,
         \DLX_Datapath/RegisterFile/N24697 ,
         \DLX_Datapath/RegisterFile/N24696 ,
         \DLX_Datapath/RegisterFile/N24695 ,
         \DLX_Datapath/RegisterFile/N24694 ,
         \DLX_Datapath/RegisterFile/N24690 ,
         \DLX_Datapath/RegisterFile/N24689 ,
         \DLX_Datapath/RegisterFile/N24688 ,
         \DLX_Datapath/RegisterFile/N24687 ,
         \DLX_Datapath/RegisterFile/N24686 ,
         \DLX_Datapath/RegisterFile/N24685 ,
         \DLX_Datapath/RegisterFile/N24683 ,
         \DLX_Datapath/RegisterFile/N24682 ,
         \DLX_Datapath/RegisterFile/N24681 ,
         \DLX_Datapath/RegisterFile/N24680 ,
         \DLX_Datapath/RegisterFile/N24679 ,
         \DLX_Datapath/RegisterFile/N24678 ,
         \DLX_Datapath/RegisterFile/N24677 ,
         \DLX_Datapath/RegisterFile/N24676 ,
         \DLX_Datapath/RegisterFile/N24675 ,
         \DLX_Datapath/RegisterFile/N24674 ,
         \DLX_Datapath/RegisterFile/N24673 ,
         \DLX_Datapath/RegisterFile/N24672 ,
         \DLX_Datapath/RegisterFile/N24671 ,
         \DLX_Datapath/RegisterFile/N24670 ,
         \DLX_Datapath/RegisterFile/N24669 ,
         \DLX_Datapath/RegisterFile/N24668 ,
         \DLX_Datapath/RegisterFile/N24667 ,
         \DLX_Datapath/RegisterFile/N24666 ,
         \DLX_Datapath/RegisterFile/N24665 ,
         \DLX_Datapath/RegisterFile/N24664 ,
         \DLX_Datapath/RegisterFile/N24663 ,
         \DLX_Datapath/RegisterFile/N24662 ,
         \DLX_Datapath/RegisterFile/N24661 ,
         \DLX_Datapath/RegisterFile/N24660 ,
         \DLX_Datapath/RegisterFile/N24659 ,
         \DLX_Datapath/RegisterFile/N24658 ,
         \DLX_Datapath/RegisterFile/N24657 ,
         \DLX_Datapath/RegisterFile/N24656 ,
         \DLX_Datapath/RegisterFile/N24655 ,
         \DLX_Datapath/RegisterFile/N24654 ,
         \DLX_Datapath/RegisterFile/N24653 ,
         \DLX_Datapath/RegisterFile/N24652 ,
         \DLX_Datapath/RegisterFile/N24651 ,
         \DLX_Datapath/RegisterFile/N24650 ,
         \DLX_Datapath/RegisterFile/N24649 ,
         \DLX_Datapath/RegisterFile/N24648 ,
         \DLX_Datapath/RegisterFile/N24647 ,
         \DLX_Datapath/RegisterFile/N24646 ,
         \DLX_Datapath/RegisterFile/N24645 ,
         \DLX_Datapath/RegisterFile/N24644 ,
         \DLX_Datapath/RegisterFile/N24643 ,
         \DLX_Datapath/RegisterFile/N24642 ,
         \DLX_Datapath/RegisterFile/N24641 ,
         \DLX_Datapath/RegisterFile/N24640 ,
         \DLX_Datapath/RegisterFile/N24639 ,
         \DLX_Datapath/RegisterFile/N24638 ,
         \DLX_Datapath/RegisterFile/N24637 ,
         \DLX_Datapath/RegisterFile/N24636 ,
         \DLX_Datapath/RegisterFile/N24635 ,
         \DLX_Datapath/RegisterFile/N24632 ,
         \DLX_Datapath/RegisterFile/N24631 ,
         \DLX_Datapath/RegisterFile/N24630 ,
         \DLX_Datapath/RegisterFile/N24628 ,
         \DLX_Datapath/RegisterFile/N24625 ,
         \DLX_Datapath/RegisterFile/N24624 ,
         \DLX_Datapath/RegisterFile/N24619 ,
         \DLX_Datapath/RegisterFile/N24618 ,
         \DLX_Datapath/RegisterFile/N24617 ,
         \DLX_Datapath/RegisterFile/N24616 ,
         \DLX_Datapath/RegisterFile/N24615 ,
         \DLX_Datapath/RegisterFile/N24614 ,
         \DLX_Datapath/RegisterFile/N24613 ,
         \DLX_Datapath/RegisterFile/N24612 ,
         \DLX_Datapath/RegisterFile/N24611 ,
         \DLX_Datapath/RegisterFile/N24610 ,
         \DLX_Datapath/RegisterFile/N24609 ,
         \DLX_Datapath/RegisterFile/N24608 ,
         \DLX_Datapath/RegisterFile/N24607 ,
         \DLX_Datapath/RegisterFile/N24606 ,
         \DLX_Datapath/RegisterFile/N24605 ,
         \DLX_Datapath/RegisterFile/N24604 ,
         \DLX_Datapath/RegisterFile/N24603 ,
         \DLX_Datapath/RegisterFile/N24602 ,
         \DLX_Datapath/RegisterFile/N24601 ,
         \DLX_Datapath/RegisterFile/N24600 ,
         \DLX_Datapath/RegisterFile/N24599 ,
         \DLX_Datapath/RegisterFile/N24598 ,
         \DLX_Datapath/RegisterFile/N24597 ,
         \DLX_Datapath/RegisterFile/N24596 ,
         \DLX_Datapath/RegisterFile/N24595 ,
         \DLX_Datapath/RegisterFile/N24594 ,
         \DLX_Datapath/RegisterFile/N24593 ,
         \DLX_Datapath/RegisterFile/N24592 ,
         \DLX_Datapath/RegisterFile/N24591 ,
         \DLX_Datapath/RegisterFile/N24590 ,
         \DLX_Datapath/RegisterFile/N24589 ,
         \DLX_Datapath/RegisterFile/N24588 ,
         \DLX_Datapath/RegisterFile/N24587 ,
         \DLX_Datapath/RegisterFile/N24586 ,
         \DLX_Datapath/RegisterFile/N24585 ,
         \DLX_Datapath/RegisterFile/N24583 ,
         \DLX_Datapath/RegisterFile/N24581 ,
         \DLX_Datapath/RegisterFile/N24580 ,
         \DLX_Datapath/RegisterFile/N24579 ,
         \DLX_Datapath/RegisterFile/N24578 ,
         \DLX_Datapath/RegisterFile/N24576 ,
         \DLX_Datapath/RegisterFile/N24573 ,
         \DLX_Datapath/RegisterFile/N24572 ,
         \DLX_Datapath/RegisterFile/N24571 ,
         \DLX_Datapath/RegisterFile/N24569 ,
         \DLX_Datapath/RegisterFile/N24567 ,
         \DLX_Datapath/RegisterFile/N24566 ,
         \DLX_Datapath/RegisterFile/N24564 ,
         \DLX_Datapath/RegisterFile/N24563 ,
         \DLX_Datapath/RegisterFile/N24562 ,
         \DLX_Datapath/RegisterFile/N24560 ,
         \DLX_Datapath/RegisterFile/N24559 ,
         \DLX_Datapath/RegisterFile/N24558 ,
         \DLX_Datapath/RegisterFile/N24557 ,
         \DLX_Datapath/RegisterFile/N24555 ,
         \DLX_Datapath/RegisterFile/N24554 ,
         \DLX_Datapath/RegisterFile/N24553 ,
         \DLX_Datapath/RegisterFile/N24552 ,
         \DLX_Datapath/RegisterFile/N24551 ,
         \DLX_Datapath/RegisterFile/N24550 ,
         \DLX_Datapath/RegisterFile/N24549 ,
         \DLX_Datapath/RegisterFile/N24548 ,
         \DLX_Datapath/RegisterFile/N24547 ,
         \DLX_Datapath/RegisterFile/N24546 ,
         \DLX_Datapath/RegisterFile/N24545 ,
         \DLX_Datapath/RegisterFile/N24544 ,
         \DLX_Datapath/RegisterFile/N24543 ,
         \DLX_Datapath/RegisterFile/N24542 ,
         \DLX_Datapath/RegisterFile/N24541 ,
         \DLX_Datapath/RegisterFile/N24540 ,
         \DLX_Datapath/RegisterFile/N24539 ,
         \DLX_Datapath/RegisterFile/N24538 ,
         \DLX_Datapath/RegisterFile/N24537 ,
         \DLX_Datapath/RegisterFile/N24536 ,
         \DLX_Datapath/RegisterFile/N24535 ,
         \DLX_Datapath/RegisterFile/N24534 ,
         \DLX_Datapath/RegisterFile/N24533 ,
         \DLX_Datapath/RegisterFile/N24532 ,
         \DLX_Datapath/RegisterFile/N24531 ,
         \DLX_Datapath/RegisterFile/N24530 ,
         \DLX_Datapath/RegisterFile/N24529 ,
         \DLX_Datapath/RegisterFile/N24528 ,
         \DLX_Datapath/RegisterFile/N24527 ,
         \DLX_Datapath/RegisterFile/N24526 ,
         \DLX_Datapath/RegisterFile/N24525 ,
         \DLX_Datapath/RegisterFile/N24524 ,
         \DLX_Datapath/RegisterFile/N24523 ,
         \DLX_Datapath/RegisterFile/N24522 ,
         \DLX_Datapath/RegisterFile/N24521 ,
         \DLX_Datapath/RegisterFile/N24520 ,
         \DLX_Datapath/RegisterFile/N24519 ,
         \DLX_Datapath/RegisterFile/N24518 ,
         \DLX_Datapath/RegisterFile/N24517 ,
         \DLX_Datapath/RegisterFile/N24516 ,
         \DLX_Datapath/RegisterFile/N24515 ,
         \DLX_Datapath/RegisterFile/N24514 ,
         \DLX_Datapath/RegisterFile/N24513 ,
         \DLX_Datapath/RegisterFile/N24512 ,
         \DLX_Datapath/RegisterFile/N24511 ,
         \DLX_Datapath/RegisterFile/N24510 ,
         \DLX_Datapath/RegisterFile/N24509 ,
         \DLX_Datapath/RegisterFile/N24508 ,
         \DLX_Datapath/RegisterFile/N24507 ,
         \DLX_Datapath/RegisterFile/N24506 ,
         \DLX_Datapath/RegisterFile/N24505 ,
         \DLX_Datapath/RegisterFile/N24504 ,
         \DLX_Datapath/RegisterFile/N24503 ,
         \DLX_Datapath/RegisterFile/N24502 ,
         \DLX_Datapath/RegisterFile/N24501 ,
         \DLX_Datapath/RegisterFile/N24500 ,
         \DLX_Datapath/RegisterFile/N24499 ,
         \DLX_Datapath/RegisterFile/N24498 ,
         \DLX_Datapath/RegisterFile/N24497 ,
         \DLX_Datapath/RegisterFile/N24496 ,
         \DLX_Datapath/RegisterFile/N24495 ,
         \DLX_Datapath/RegisterFile/N24494 ,
         \DLX_Datapath/RegisterFile/N24493 ,
         \DLX_Datapath/RegisterFile/N24492 ,
         \DLX_Datapath/RegisterFile/N24491 ,
         \DLX_Datapath/RegisterFile/N24490 ,
         \DLX_Datapath/RegisterFile/N24489 ,
         \DLX_Datapath/RegisterFile/N24488 ,
         \DLX_Datapath/RegisterFile/N24487 ,
         \DLX_Datapath/RegisterFile/N24486 ,
         \DLX_Datapath/RegisterFile/N24485 ,
         \DLX_Datapath/RegisterFile/N24484 ,
         \DLX_Datapath/RegisterFile/N24483 ,
         \DLX_Datapath/RegisterFile/N24482 ,
         \DLX_Datapath/RegisterFile/N24481 ,
         \DLX_Datapath/RegisterFile/N24480 ,
         \DLX_Datapath/RegisterFile/N24479 ,
         \DLX_Datapath/RegisterFile/N24478 ,
         \DLX_Datapath/RegisterFile/N24477 ,
         \DLX_Datapath/RegisterFile/N24476 ,
         \DLX_Datapath/RegisterFile/N24475 ,
         \DLX_Datapath/RegisterFile/N24474 ,
         \DLX_Datapath/RegisterFile/N24473 ,
         \DLX_Datapath/RegisterFile/N24472 ,
         \DLX_Datapath/RegisterFile/N24471 ,
         \DLX_Datapath/RegisterFile/N24470 ,
         \DLX_Datapath/RegisterFile/N24469 ,
         \DLX_Datapath/RegisterFile/N24468 ,
         \DLX_Datapath/RegisterFile/N24467 ,
         \DLX_Datapath/RegisterFile/N24466 ,
         \DLX_Datapath/RegisterFile/N24465 ,
         \DLX_Datapath/RegisterFile/N24464 ,
         \DLX_Datapath/RegisterFile/N24463 ,
         \DLX_Datapath/RegisterFile/N24462 ,
         \DLX_Datapath/RegisterFile/N24461 ,
         \DLX_Datapath/RegisterFile/N24460 ,
         \DLX_Datapath/RegisterFile/N24459 ,
         \DLX_Datapath/RegisterFile/N24457 ,
         \DLX_Datapath/RegisterFile/N24456 ,
         \DLX_Datapath/RegisterFile/N24455 ,
         \DLX_Datapath/RegisterFile/N24453 ,
         \DLX_Datapath/RegisterFile/N24451 ,
         \DLX_Datapath/RegisterFile/N24450 ,
         \DLX_Datapath/RegisterFile/N24448 ,
         \DLX_Datapath/RegisterFile/N24445 ,
         \DLX_Datapath/RegisterFile/N24444 ,
         \DLX_Datapath/RegisterFile/N24443 ,
         \DLX_Datapath/RegisterFile/N24441 ,
         \DLX_Datapath/RegisterFile/N24439 ,
         \DLX_Datapath/RegisterFile/N24438 ,
         \DLX_Datapath/RegisterFile/N24436 ,
         \DLX_Datapath/RegisterFile/N24435 ,
         \DLX_Datapath/RegisterFile/N24434 ,
         \DLX_Datapath/RegisterFile/N24432 ,
         \DLX_Datapath/RegisterFile/N24431 ,
         \DLX_Datapath/RegisterFile/N24430 ,
         \DLX_Datapath/RegisterFile/N24429 ,
         \DLX_Datapath/RegisterFile/N24427 ,
         \DLX_Datapath/RegisterFile/N24426 ,
         \DLX_Datapath/RegisterFile/N24425 ,
         \DLX_Datapath/RegisterFile/N24424 ,
         \DLX_Datapath/RegisterFile/N24423 ,
         \DLX_Datapath/RegisterFile/N24422 ,
         \DLX_Datapath/RegisterFile/N24421 ,
         \DLX_Datapath/RegisterFile/N24420 ,
         \DLX_Datapath/RegisterFile/N24419 ,
         \DLX_Datapath/RegisterFile/N24418 ,
         \DLX_Datapath/RegisterFile/N24417 ,
         \DLX_Datapath/RegisterFile/N24416 ,
         \DLX_Datapath/RegisterFile/N24415 ,
         \DLX_Datapath/RegisterFile/N24414 ,
         \DLX_Datapath/RegisterFile/N24413 ,
         \DLX_Datapath/RegisterFile/N24412 ,
         \DLX_Datapath/RegisterFile/N24411 ,
         \DLX_Datapath/RegisterFile/N24410 ,
         \DLX_Datapath/RegisterFile/N24409 ,
         \DLX_Datapath/RegisterFile/N24408 ,
         \DLX_Datapath/RegisterFile/N24407 ,
         \DLX_Datapath/RegisterFile/N24406 ,
         \DLX_Datapath/RegisterFile/N24405 ,
         \DLX_Datapath/RegisterFile/N24404 ,
         \DLX_Datapath/RegisterFile/N24403 ,
         \DLX_Datapath/RegisterFile/N24402 ,
         \DLX_Datapath/RegisterFile/N24401 ,
         \DLX_Datapath/RegisterFile/N24400 ,
         \DLX_Datapath/RegisterFile/N24399 ,
         \DLX_Datapath/RegisterFile/N24398 ,
         \DLX_Datapath/RegisterFile/N24397 ,
         \DLX_Datapath/RegisterFile/N24396 ,
         \DLX_Datapath/RegisterFile/N24395 ,
         \DLX_Datapath/RegisterFile/N24393 ,
         \DLX_Datapath/RegisterFile/N24392 ,
         \DLX_Datapath/RegisterFile/N24391 ,
         \DLX_Datapath/RegisterFile/N24390 ,
         \DLX_Datapath/RegisterFile/N24389 ,
         \DLX_Datapath/RegisterFile/N24388 ,
         \DLX_Datapath/RegisterFile/N24387 ,
         \DLX_Datapath/RegisterFile/N24386 ,
         \DLX_Datapath/RegisterFile/N24385 ,
         \DLX_Datapath/RegisterFile/N24384 ,
         \DLX_Datapath/RegisterFile/N24383 ,
         \DLX_Datapath/RegisterFile/N24382 ,
         \DLX_Datapath/RegisterFile/N24381 ,
         \DLX_Datapath/RegisterFile/N24380 ,
         \DLX_Datapath/RegisterFile/N24379 ,
         \DLX_Datapath/RegisterFile/N24377 ,
         \DLX_Datapath/RegisterFile/N24375 ,
         \DLX_Datapath/RegisterFile/N24374 ,
         \DLX_Datapath/RegisterFile/N24372 ,
         \DLX_Datapath/RegisterFile/N24371 ,
         \DLX_Datapath/RegisterFile/N24370 ,
         \DLX_Datapath/RegisterFile/N24368 ,
         \DLX_Datapath/RegisterFile/N24365 ,
         \DLX_Datapath/RegisterFile/N24363 ,
         \DLX_Datapath/RegisterFile/N24362 ,
         \DLX_Datapath/RegisterFile/N24361 ,
         \DLX_Datapath/RegisterFile/N24360 ,
         \DLX_Datapath/RegisterFile/N24359 ,
         \DLX_Datapath/RegisterFile/N24358 ,
         \DLX_Datapath/RegisterFile/N24357 ,
         \DLX_Datapath/RegisterFile/N24356 ,
         \DLX_Datapath/RegisterFile/N24355 ,
         \DLX_Datapath/RegisterFile/N24354 ,
         \DLX_Datapath/RegisterFile/N24353 ,
         \DLX_Datapath/RegisterFile/N24352 ,
         \DLX_Datapath/RegisterFile/N24351 ,
         \DLX_Datapath/RegisterFile/N24350 ,
         \DLX_Datapath/RegisterFile/N24349 ,
         \DLX_Datapath/RegisterFile/N24348 ,
         \DLX_Datapath/RegisterFile/N24347 ,
         \DLX_Datapath/RegisterFile/N24346 ,
         \DLX_Datapath/RegisterFile/N24345 ,
         \DLX_Datapath/RegisterFile/N24344 ,
         \DLX_Datapath/RegisterFile/N24343 ,
         \DLX_Datapath/RegisterFile/N24342 ,
         \DLX_Datapath/RegisterFile/N24341 ,
         \DLX_Datapath/RegisterFile/N24340 ,
         \DLX_Datapath/RegisterFile/N24339 ,
         \DLX_Datapath/RegisterFile/N24338 ,
         \DLX_Datapath/RegisterFile/N24337 ,
         \DLX_Datapath/RegisterFile/N24336 ,
         \DLX_Datapath/RegisterFile/N24335 ,
         \DLX_Datapath/RegisterFile/N24334 ,
         \DLX_Datapath/RegisterFile/N24333 ,
         \DLX_Datapath/RegisterFile/N24332 ,
         \DLX_Datapath/RegisterFile/N24331 ,
         \DLX_Datapath/RegisterFile/N24330 ,
         \DLX_Datapath/RegisterFile/N24329 ,
         \DLX_Datapath/RegisterFile/N24328 ,
         \DLX_Datapath/RegisterFile/N24327 ,
         \DLX_Datapath/RegisterFile/N24326 ,
         \DLX_Datapath/RegisterFile/N24325 ,
         \DLX_Datapath/RegisterFile/N24324 ,
         \DLX_Datapath/RegisterFile/N24323 ,
         \DLX_Datapath/RegisterFile/N24322 ,
         \DLX_Datapath/RegisterFile/N24320 ,
         \DLX_Datapath/RegisterFile/N24318 ,
         \DLX_Datapath/RegisterFile/N24317 ,
         \DLX_Datapath/RegisterFile/N24316 ,
         \DLX_Datapath/RegisterFile/N24315 ,
         \DLX_Datapath/RegisterFile/N24311 ,
         \DLX_Datapath/RegisterFile/N24310 ,
         \DLX_Datapath/RegisterFile/N24308 ,
         \DLX_Datapath/RegisterFile/N24307 ,
         \DLX_Datapath/RegisterFile/N24306 ,
         \DLX_Datapath/RegisterFile/N24304 ,
         \DLX_Datapath/RegisterFile/N24303 ,
         \DLX_Datapath/RegisterFile/N24302 ,
         \DLX_Datapath/RegisterFile/N24301 ,
         \DLX_Datapath/RegisterFile/N24299 ,
         \DLX_Datapath/RegisterFile/N24298 ,
         \DLX_Datapath/RegisterFile/N24297 ,
         \DLX_Datapath/RegisterFile/N24296 ,
         \DLX_Datapath/RegisterFile/N24295 ,
         \DLX_Datapath/RegisterFile/N24294 ,
         \DLX_Datapath/RegisterFile/N24293 ,
         \DLX_Datapath/RegisterFile/N24292 ,
         \DLX_Datapath/RegisterFile/N24291 ,
         \DLX_Datapath/RegisterFile/N24290 ,
         \DLX_Datapath/RegisterFile/N24289 ,
         \DLX_Datapath/RegisterFile/N24288 ,
         \DLX_Datapath/RegisterFile/N24287 ,
         \DLX_Datapath/RegisterFile/N24286 ,
         \DLX_Datapath/RegisterFile/N24285 ,
         \DLX_Datapath/RegisterFile/N24284 ,
         \DLX_Datapath/RegisterFile/N24283 ,
         \DLX_Datapath/RegisterFile/N24282 ,
         \DLX_Datapath/RegisterFile/N24281 ,
         \DLX_Datapath/RegisterFile/N24280 ,
         \DLX_Datapath/RegisterFile/N24279 ,
         \DLX_Datapath/RegisterFile/N24278 ,
         \DLX_Datapath/RegisterFile/N24277 ,
         \DLX_Datapath/RegisterFile/N24276 ,
         \DLX_Datapath/RegisterFile/N24275 ,
         \DLX_Datapath/RegisterFile/N24274 ,
         \DLX_Datapath/RegisterFile/N24273 ,
         \DLX_Datapath/RegisterFile/N24272 ,
         \DLX_Datapath/RegisterFile/N24271 ,
         \DLX_Datapath/RegisterFile/N24270 ,
         \DLX_Datapath/RegisterFile/N24269 ,
         \DLX_Datapath/RegisterFile/N24268 ,
         \DLX_Datapath/RegisterFile/N24267 ,
         \DLX_Datapath/RegisterFile/N24266 ,
         \DLX_Datapath/RegisterFile/N24265 ,
         \DLX_Datapath/RegisterFile/N24264 ,
         \DLX_Datapath/RegisterFile/N24263 ,
         \DLX_Datapath/RegisterFile/N24262 ,
         \DLX_Datapath/RegisterFile/N24261 ,
         \DLX_Datapath/RegisterFile/N24260 ,
         \DLX_Datapath/RegisterFile/N24259 ,
         \DLX_Datapath/RegisterFile/N24258 ,
         \DLX_Datapath/RegisterFile/N24257 ,
         \DLX_Datapath/RegisterFile/N24256 ,
         \DLX_Datapath/RegisterFile/N24255 ,
         \DLX_Datapath/RegisterFile/N24254 ,
         \DLX_Datapath/RegisterFile/N24253 ,
         \DLX_Datapath/RegisterFile/N24252 ,
         \DLX_Datapath/RegisterFile/N24251 ,
         \DLX_Datapath/RegisterFile/N24250 ,
         \DLX_Datapath/RegisterFile/N24249 ,
         \DLX_Datapath/RegisterFile/N24248 ,
         \DLX_Datapath/RegisterFile/N24247 ,
         \DLX_Datapath/RegisterFile/N24246 ,
         \DLX_Datapath/RegisterFile/N24245 ,
         \DLX_Datapath/RegisterFile/N24244 ,
         \DLX_Datapath/RegisterFile/N24243 ,
         \DLX_Datapath/RegisterFile/N24242 ,
         \DLX_Datapath/RegisterFile/N24241 ,
         \DLX_Datapath/RegisterFile/N24240 ,
         \DLX_Datapath/RegisterFile/N24239 ,
         \DLX_Datapath/RegisterFile/N24238 ,
         \DLX_Datapath/RegisterFile/N24237 ,
         \DLX_Datapath/RegisterFile/N24236 ,
         \DLX_Datapath/RegisterFile/N24235 ,
         \DLX_Datapath/RegisterFile/N24234 ,
         \DLX_Datapath/RegisterFile/N24233 ,
         \DLX_Datapath/RegisterFile/N24232 ,
         \DLX_Datapath/RegisterFile/N24231 ,
         \DLX_Datapath/RegisterFile/N24230 ,
         \DLX_Datapath/RegisterFile/N24229 ,
         \DLX_Datapath/RegisterFile/N24228 ,
         \DLX_Datapath/RegisterFile/N24227 ,
         \DLX_Datapath/RegisterFile/N24226 ,
         \DLX_Datapath/RegisterFile/N24225 ,
         \DLX_Datapath/RegisterFile/N24224 ,
         \DLX_Datapath/RegisterFile/N24223 ,
         \DLX_Datapath/RegisterFile/N24222 ,
         \DLX_Datapath/RegisterFile/N24221 ,
         \DLX_Datapath/RegisterFile/N24220 ,
         \DLX_Datapath/RegisterFile/N24219 ,
         \DLX_Datapath/RegisterFile/N24218 ,
         \DLX_Datapath/RegisterFile/N24217 ,
         \DLX_Datapath/RegisterFile/N24216 ,
         \DLX_Datapath/RegisterFile/N24215 ,
         \DLX_Datapath/RegisterFile/N24214 ,
         \DLX_Datapath/RegisterFile/N24213 ,
         \DLX_Datapath/RegisterFile/N24212 ,
         \DLX_Datapath/RegisterFile/N24211 ,
         \DLX_Datapath/RegisterFile/N24210 ,
         \DLX_Datapath/RegisterFile/N24209 ,
         \DLX_Datapath/RegisterFile/N24208 ,
         \DLX_Datapath/RegisterFile/N24207 ,
         \DLX_Datapath/RegisterFile/N24206 ,
         \DLX_Datapath/RegisterFile/N24205 ,
         \DLX_Datapath/RegisterFile/N24204 ,
         \DLX_Datapath/RegisterFile/N24203 ,
         \DLX_Datapath/RegisterFile/N24201 ,
         \DLX_Datapath/RegisterFile/N24200 ,
         \DLX_Datapath/RegisterFile/N24199 ,
         \DLX_Datapath/RegisterFile/N24198 ,
         \DLX_Datapath/RegisterFile/N24197 ,
         \DLX_Datapath/RegisterFile/N24196 ,
         \DLX_Datapath/RegisterFile/N24195 ,
         \DLX_Datapath/RegisterFile/N24194 ,
         \DLX_Datapath/RegisterFile/N24193 ,
         \DLX_Datapath/RegisterFile/N24192 ,
         \DLX_Datapath/RegisterFile/N24191 ,
         \DLX_Datapath/RegisterFile/N24190 ,
         \DLX_Datapath/RegisterFile/N24189 ,
         \DLX_Datapath/RegisterFile/N24188 ,
         \DLX_Datapath/RegisterFile/N24187 ,
         \DLX_Datapath/RegisterFile/N24183 ,
         \DLX_Datapath/RegisterFile/N24182 ,
         \DLX_Datapath/RegisterFile/N24180 ,
         \DLX_Datapath/RegisterFile/N24179 ,
         \DLX_Datapath/RegisterFile/N24178 ,
         \DLX_Datapath/RegisterFile/N24176 ,
         \DLX_Datapath/RegisterFile/N24175 ,
         \DLX_Datapath/RegisterFile/N24174 ,
         \DLX_Datapath/RegisterFile/N24173 ,
         \DLX_Datapath/RegisterFile/N24171 ,
         \DLX_Datapath/RegisterFile/N24170 ,
         \DLX_Datapath/RegisterFile/N24169 ,
         \DLX_Datapath/RegisterFile/N24168 ,
         \DLX_Datapath/RegisterFile/N24167 ,
         \DLX_Datapath/RegisterFile/N24166 ,
         \DLX_Datapath/RegisterFile/N24165 ,
         \DLX_Datapath/RegisterFile/N24164 ,
         \DLX_Datapath/RegisterFile/N24163 ,
         \DLX_Datapath/RegisterFile/N24162 ,
         \DLX_Datapath/RegisterFile/N24161 ,
         \DLX_Datapath/RegisterFile/N24160 ,
         \DLX_Datapath/RegisterFile/N24159 ,
         \DLX_Datapath/RegisterFile/N24158 ,
         \DLX_Datapath/RegisterFile/N24157 ,
         \DLX_Datapath/RegisterFile/N24156 ,
         \DLX_Datapath/RegisterFile/N24155 ,
         \DLX_Datapath/RegisterFile/N24154 ,
         \DLX_Datapath/RegisterFile/N24153 ,
         \DLX_Datapath/RegisterFile/N24152 ,
         \DLX_Datapath/RegisterFile/N24151 ,
         \DLX_Datapath/RegisterFile/N24150 ,
         \DLX_Datapath/RegisterFile/N24149 ,
         \DLX_Datapath/RegisterFile/N24148 ,
         \DLX_Datapath/RegisterFile/N24147 ,
         \DLX_Datapath/RegisterFile/N24146 ,
         \DLX_Datapath/RegisterFile/N24145 ,
         \DLX_Datapath/RegisterFile/N24144 ,
         \DLX_Datapath/RegisterFile/N24143 ,
         \DLX_Datapath/RegisterFile/N24142 ,
         \DLX_Datapath/RegisterFile/N24141 ,
         \DLX_Datapath/RegisterFile/N24140 ,
         \DLX_Datapath/RegisterFile/N24139 ,
         \DLX_Datapath/RegisterFile/N24138 ,
         \DLX_Datapath/RegisterFile/N24137 ,
         \DLX_Datapath/RegisterFile/N24136 ,
         \DLX_Datapath/RegisterFile/N24135 ,
         \DLX_Datapath/RegisterFile/N24134 ,
         \DLX_Datapath/RegisterFile/N24133 ,
         \DLX_Datapath/RegisterFile/N24132 ,
         \DLX_Datapath/RegisterFile/N24131 ,
         \DLX_Datapath/RegisterFile/N24130 ,
         \DLX_Datapath/RegisterFile/N24129 ,
         \DLX_Datapath/RegisterFile/N24128 ,
         \DLX_Datapath/RegisterFile/N24127 ,
         \DLX_Datapath/RegisterFile/N24126 ,
         \DLX_Datapath/RegisterFile/N24125 ,
         \DLX_Datapath/RegisterFile/N24124 ,
         \DLX_Datapath/RegisterFile/N24123 ,
         \DLX_Datapath/RegisterFile/N24118 ,
         \DLX_Datapath/RegisterFile/N24116 ,
         \DLX_Datapath/RegisterFile/N24115 ,
         \DLX_Datapath/RegisterFile/N24114 ,
         \DLX_Datapath/RegisterFile/N24110 ,
         \DLX_Datapath/RegisterFile/N24107 ,
         \DLX_Datapath/RegisterFile/N24106 ,
         \DLX_Datapath/RegisterFile/N24105 ,
         \DLX_Datapath/RegisterFile/N24104 ,
         \DLX_Datapath/RegisterFile/N24103 ,
         \DLX_Datapath/RegisterFile/N24102 ,
         \DLX_Datapath/RegisterFile/N24101 ,
         \DLX_Datapath/RegisterFile/N24100 ,
         \DLX_Datapath/RegisterFile/N24099 ,
         \DLX_Datapath/RegisterFile/N24098 ,
         \DLX_Datapath/RegisterFile/N24097 ,
         \DLX_Datapath/RegisterFile/N24096 ,
         \DLX_Datapath/RegisterFile/N24095 ,
         \DLX_Datapath/RegisterFile/N24094 ,
         \DLX_Datapath/RegisterFile/N24093 ,
         \DLX_Datapath/RegisterFile/N24092 ,
         \DLX_Datapath/RegisterFile/N24091 ,
         \DLX_Datapath/RegisterFile/N24090 ,
         \DLX_Datapath/RegisterFile/N24089 ,
         \DLX_Datapath/RegisterFile/N24088 ,
         \DLX_Datapath/RegisterFile/N24087 ,
         \DLX_Datapath/RegisterFile/N24086 ,
         \DLX_Datapath/RegisterFile/N24085 ,
         \DLX_Datapath/RegisterFile/N24084 ,
         \DLX_Datapath/RegisterFile/N24083 ,
         \DLX_Datapath/RegisterFile/N24082 ,
         \DLX_Datapath/RegisterFile/N24081 ,
         \DLX_Datapath/RegisterFile/N24080 ,
         \DLX_Datapath/RegisterFile/N24079 ,
         \DLX_Datapath/RegisterFile/N24078 ,
         \DLX_Datapath/RegisterFile/N24077 ,
         \DLX_Datapath/RegisterFile/N24076 ,
         \DLX_Datapath/RegisterFile/N24075 ,
         \DLX_Datapath/RegisterFile/N24073 ,
         \DLX_Datapath/RegisterFile/N24072 ,
         \DLX_Datapath/RegisterFile/N24071 ,
         \DLX_Datapath/RegisterFile/N24069 ,
         \DLX_Datapath/RegisterFile/N24067 ,
         \DLX_Datapath/RegisterFile/N24066 ,
         \DLX_Datapath/RegisterFile/N24065 ,
         \DLX_Datapath/RegisterFile/N24064 ,
         \DLX_Datapath/RegisterFile/N24063 ,
         \DLX_Datapath/RegisterFile/N24061 ,
         \DLX_Datapath/RegisterFile/N24060 ,
         \DLX_Datapath/RegisterFile/N24059 ,
         \DLX_Datapath/RegisterFile/N24054 ,
         \DLX_Datapath/RegisterFile/N24052 ,
         \DLX_Datapath/RegisterFile/N24051 ,
         \DLX_Datapath/RegisterFile/N24050 ,
         \DLX_Datapath/RegisterFile/N24048 ,
         \DLX_Datapath/RegisterFile/N24047 ,
         \DLX_Datapath/RegisterFile/N24046 ,
         \DLX_Datapath/RegisterFile/N24045 ,
         \DLX_Datapath/RegisterFile/N24043 ,
         \DLX_Datapath/RegisterFile/N24042 ,
         \DLX_Datapath/RegisterFile/N24041 ,
         \DLX_Datapath/RegisterFile/N24040 ,
         \DLX_Datapath/RegisterFile/N24039 ,
         \DLX_Datapath/RegisterFile/N24038 ,
         \DLX_Datapath/RegisterFile/N24037 ,
         \DLX_Datapath/RegisterFile/N24036 ,
         \DLX_Datapath/RegisterFile/N24035 ,
         \DLX_Datapath/RegisterFile/N24034 ,
         \DLX_Datapath/RegisterFile/N24033 ,
         \DLX_Datapath/RegisterFile/N24032 ,
         \DLX_Datapath/RegisterFile/N24031 ,
         \DLX_Datapath/RegisterFile/N24030 ,
         \DLX_Datapath/RegisterFile/N24029 ,
         \DLX_Datapath/RegisterFile/N24028 ,
         \DLX_Datapath/RegisterFile/N24027 ,
         \DLX_Datapath/RegisterFile/N24026 ,
         \DLX_Datapath/RegisterFile/N24025 ,
         \DLX_Datapath/RegisterFile/N24024 ,
         \DLX_Datapath/RegisterFile/N24023 ,
         \DLX_Datapath/RegisterFile/N24022 ,
         \DLX_Datapath/RegisterFile/N24021 ,
         \DLX_Datapath/RegisterFile/N24020 ,
         \DLX_Datapath/RegisterFile/N24019 ,
         \DLX_Datapath/RegisterFile/N24018 ,
         \DLX_Datapath/RegisterFile/N24017 ,
         \DLX_Datapath/RegisterFile/N24016 ,
         \DLX_Datapath/RegisterFile/N24015 ,
         \DLX_Datapath/RegisterFile/N24014 ,
         \DLX_Datapath/RegisterFile/N24013 ,
         \DLX_Datapath/RegisterFile/N24012 ,
         \DLX_Datapath/RegisterFile/N24011 ,
         \DLX_Datapath/RegisterFile/N24010 ,
         \DLX_Datapath/RegisterFile/N24009 ,
         \DLX_Datapath/RegisterFile/N24008 ,
         \DLX_Datapath/RegisterFile/N24007 ,
         \DLX_Datapath/RegisterFile/N24006 ,
         \DLX_Datapath/RegisterFile/N24005 ,
         \DLX_Datapath/RegisterFile/N24004 ,
         \DLX_Datapath/RegisterFile/N24003 ,
         \DLX_Datapath/RegisterFile/N24002 ,
         \DLX_Datapath/RegisterFile/N24001 ,
         \DLX_Datapath/RegisterFile/N24000 ,
         \DLX_Datapath/RegisterFile/N23999 ,
         \DLX_Datapath/RegisterFile/N23998 ,
         \DLX_Datapath/RegisterFile/N23997 ,
         \DLX_Datapath/RegisterFile/N23996 ,
         \DLX_Datapath/RegisterFile/N23995 ,
         \DLX_Datapath/RegisterFile/N23994 ,
         \DLX_Datapath/RegisterFile/N23993 ,
         \DLX_Datapath/RegisterFile/N23992 ,
         \DLX_Datapath/RegisterFile/N23991 ,
         \DLX_Datapath/RegisterFile/N23990 ,
         \DLX_Datapath/RegisterFile/N23989 ,
         \DLX_Datapath/RegisterFile/N23988 ,
         \DLX_Datapath/RegisterFile/N23987 ,
         \DLX_Datapath/RegisterFile/N23986 ,
         \DLX_Datapath/RegisterFile/N23985 ,
         \DLX_Datapath/RegisterFile/N23984 ,
         \DLX_Datapath/RegisterFile/N23983 ,
         \DLX_Datapath/RegisterFile/N23982 ,
         \DLX_Datapath/RegisterFile/N23981 ,
         \DLX_Datapath/RegisterFile/N23980 ,
         \DLX_Datapath/RegisterFile/N23979 ,
         \DLX_Datapath/RegisterFile/N23978 ,
         \DLX_Datapath/RegisterFile/N23977 ,
         \DLX_Datapath/RegisterFile/N23976 ,
         \DLX_Datapath/RegisterFile/N23975 ,
         \DLX_Datapath/RegisterFile/N23974 ,
         \DLX_Datapath/RegisterFile/N23973 ,
         \DLX_Datapath/RegisterFile/N23972 ,
         \DLX_Datapath/RegisterFile/N23971 ,
         \DLX_Datapath/RegisterFile/N23970 ,
         \DLX_Datapath/RegisterFile/N23969 ,
         \DLX_Datapath/RegisterFile/N23968 ,
         \DLX_Datapath/RegisterFile/N23967 ,
         \DLX_Datapath/RegisterFile/N23966 ,
         \DLX_Datapath/RegisterFile/N23965 ,
         \DLX_Datapath/RegisterFile/N23964 ,
         \DLX_Datapath/RegisterFile/N23963 ,
         \DLX_Datapath/RegisterFile/N23962 ,
         \DLX_Datapath/RegisterFile/N23961 ,
         \DLX_Datapath/RegisterFile/N23960 ,
         \DLX_Datapath/RegisterFile/N23959 ,
         \DLX_Datapath/RegisterFile/N23958 ,
         \DLX_Datapath/RegisterFile/N23957 ,
         \DLX_Datapath/RegisterFile/N23956 ,
         \DLX_Datapath/RegisterFile/N23955 ,
         \DLX_Datapath/RegisterFile/N23954 ,
         \DLX_Datapath/RegisterFile/N23953 ,
         \DLX_Datapath/RegisterFile/N23952 ,
         \DLX_Datapath/RegisterFile/N23951 ,
         \DLX_Datapath/RegisterFile/N23950 ,
         \DLX_Datapath/RegisterFile/N23949 ,
         \DLX_Datapath/RegisterFile/N23948 ,
         \DLX_Datapath/RegisterFile/N23947 ,
         \DLX_Datapath/RegisterFile/N23945 ,
         \DLX_Datapath/RegisterFile/N23944 ,
         \DLX_Datapath/RegisterFile/N23943 ,
         \DLX_Datapath/RegisterFile/N23941 ,
         \DLX_Datapath/RegisterFile/N23939 ,
         \DLX_Datapath/RegisterFile/N23938 ,
         \DLX_Datapath/RegisterFile/N23936 ,
         \DLX_Datapath/RegisterFile/N23933 ,
         \DLX_Datapath/RegisterFile/N23932 ,
         \DLX_Datapath/RegisterFile/N23931 ,
         \DLX_Datapath/RegisterFile/N23929 ,
         \DLX_Datapath/RegisterFile/N23926 ,
         \DLX_Datapath/RegisterFile/N23924 ,
         \DLX_Datapath/RegisterFile/N23923 ,
         \DLX_Datapath/RegisterFile/N23922 ,
         \DLX_Datapath/RegisterFile/N23920 ,
         \DLX_Datapath/RegisterFile/N23919 ,
         \DLX_Datapath/RegisterFile/N23918 ,
         \DLX_Datapath/RegisterFile/N23917 ,
         \DLX_Datapath/RegisterFile/N23915 ,
         \DLX_Datapath/RegisterFile/N23914 ,
         \DLX_Datapath/RegisterFile/N23913 ,
         \DLX_Datapath/RegisterFile/N23912 ,
         \DLX_Datapath/RegisterFile/N23911 ,
         \DLX_Datapath/RegisterFile/N23910 ,
         \DLX_Datapath/RegisterFile/N23909 ,
         \DLX_Datapath/RegisterFile/N23908 ,
         \DLX_Datapath/RegisterFile/N23907 ,
         \DLX_Datapath/RegisterFile/N23906 ,
         \DLX_Datapath/RegisterFile/N23905 ,
         \DLX_Datapath/RegisterFile/N23904 ,
         \DLX_Datapath/RegisterFile/N23903 ,
         \DLX_Datapath/RegisterFile/N23902 ,
         \DLX_Datapath/RegisterFile/N23901 ,
         \DLX_Datapath/RegisterFile/N23900 ,
         \DLX_Datapath/RegisterFile/N23899 ,
         \DLX_Datapath/RegisterFile/N23898 ,
         \DLX_Datapath/RegisterFile/N23897 ,
         \DLX_Datapath/RegisterFile/N23896 ,
         \DLX_Datapath/RegisterFile/N23895 ,
         \DLX_Datapath/RegisterFile/N23894 ,
         \DLX_Datapath/RegisterFile/N23893 ,
         \DLX_Datapath/RegisterFile/N23892 ,
         \DLX_Datapath/RegisterFile/N23891 ,
         \DLX_Datapath/RegisterFile/N23890 ,
         \DLX_Datapath/RegisterFile/N23889 ,
         \DLX_Datapath/RegisterFile/N23888 ,
         \DLX_Datapath/RegisterFile/N23887 ,
         \DLX_Datapath/RegisterFile/N23886 ,
         \DLX_Datapath/RegisterFile/N23885 ,
         \DLX_Datapath/RegisterFile/N23884 ,
         \DLX_Datapath/RegisterFile/N23883 ,
         \DLX_Datapath/RegisterFile/N23881 ,
         \DLX_Datapath/RegisterFile/N23880 ,
         \DLX_Datapath/RegisterFile/N23879 ,
         \DLX_Datapath/RegisterFile/N23878 ,
         \DLX_Datapath/RegisterFile/N23877 ,
         \DLX_Datapath/RegisterFile/N23876 ,
         \DLX_Datapath/RegisterFile/N23875 ,
         \DLX_Datapath/RegisterFile/N23874 ,
         \DLX_Datapath/RegisterFile/N23873 ,
         \DLX_Datapath/RegisterFile/N23872 ,
         \DLX_Datapath/RegisterFile/N23871 ,
         \DLX_Datapath/RegisterFile/N23870 ,
         \DLX_Datapath/RegisterFile/N23869 ,
         \DLX_Datapath/RegisterFile/N23868 ,
         \DLX_Datapath/RegisterFile/N23867 ,
         \DLX_Datapath/RegisterFile/N23865 ,
         \DLX_Datapath/RegisterFile/N23862 ,
         \DLX_Datapath/RegisterFile/N23860 ,
         \DLX_Datapath/RegisterFile/N23859 ,
         \DLX_Datapath/RegisterFile/N23858 ,
         \DLX_Datapath/RegisterFile/N23856 ,
         \DLX_Datapath/RegisterFile/N23854 ,
         \DLX_Datapath/RegisterFile/N23851 ,
         \DLX_Datapath/RegisterFile/N23850 ,
         \DLX_Datapath/RegisterFile/N23849 ,
         \DLX_Datapath/RegisterFile/N23848 ,
         \DLX_Datapath/RegisterFile/N23847 ,
         \DLX_Datapath/RegisterFile/N23846 ,
         \DLX_Datapath/RegisterFile/N23845 ,
         \DLX_Datapath/RegisterFile/N23844 ,
         \DLX_Datapath/RegisterFile/N23843 ,
         \DLX_Datapath/RegisterFile/N23842 ,
         \DLX_Datapath/RegisterFile/N23841 ,
         \DLX_Datapath/RegisterFile/N23840 ,
         \DLX_Datapath/RegisterFile/N23839 ,
         \DLX_Datapath/RegisterFile/N23838 ,
         \DLX_Datapath/RegisterFile/N23837 ,
         \DLX_Datapath/RegisterFile/N23836 ,
         \DLX_Datapath/RegisterFile/N23835 ,
         \DLX_Datapath/RegisterFile/N23834 ,
         \DLX_Datapath/RegisterFile/N23833 ,
         \DLX_Datapath/RegisterFile/N23832 ,
         \DLX_Datapath/RegisterFile/N23831 ,
         \DLX_Datapath/RegisterFile/N23830 ,
         \DLX_Datapath/RegisterFile/N23829 ,
         \DLX_Datapath/RegisterFile/N23828 ,
         \DLX_Datapath/RegisterFile/N23827 ,
         \DLX_Datapath/RegisterFile/N23826 ,
         \DLX_Datapath/RegisterFile/N23825 ,
         \DLX_Datapath/RegisterFile/N23824 ,
         \DLX_Datapath/RegisterFile/N23823 ,
         \DLX_Datapath/RegisterFile/N23822 ,
         \DLX_Datapath/RegisterFile/N23821 ,
         \DLX_Datapath/RegisterFile/N23820 ,
         \DLX_Datapath/RegisterFile/N23819 ,
         \DLX_Datapath/RegisterFile/N23818 ,
         \DLX_Datapath/RegisterFile/N23817 ,
         \DLX_Datapath/RegisterFile/N23816 ,
         \DLX_Datapath/RegisterFile/N23814 ,
         \DLX_Datapath/RegisterFile/N23813 ,
         \DLX_Datapath/RegisterFile/N23812 ,
         \DLX_Datapath/RegisterFile/N23811 ,
         \DLX_Datapath/RegisterFile/N23810 ,
         \DLX_Datapath/RegisterFile/N23809 ,
         \DLX_Datapath/RegisterFile/N23808 ,
         \DLX_Datapath/RegisterFile/N23807 ,
         \DLX_Datapath/RegisterFile/N23805 ,
         \DLX_Datapath/RegisterFile/N23803 ,
         \DLX_Datapath/RegisterFile/N23799 ,
         \DLX_Datapath/RegisterFile/N23798 ,
         \DLX_Datapath/RegisterFile/N23797 ,
         \DLX_Datapath/RegisterFile/N23795 ,
         \DLX_Datapath/RegisterFile/N23794 ,
         \DLX_Datapath/RegisterFile/N23793 ,
         \DLX_Datapath/RegisterFile/N23792 ,
         \DLX_Datapath/RegisterFile/N23791 ,
         \DLX_Datapath/RegisterFile/N23790 ,
         \DLX_Datapath/RegisterFile/N23789 ,
         \DLX_Datapath/RegisterFile/N23787 ,
         \DLX_Datapath/RegisterFile/N23786 ,
         \DLX_Datapath/RegisterFile/N23785 ,
         \DLX_Datapath/RegisterFile/N23784 ,
         \DLX_Datapath/RegisterFile/N23783 ,
         \DLX_Datapath/RegisterFile/N23782 ,
         \DLX_Datapath/RegisterFile/N23781 ,
         \DLX_Datapath/RegisterFile/N23780 ,
         \DLX_Datapath/RegisterFile/N23779 ,
         \DLX_Datapath/RegisterFile/N23778 ,
         \DLX_Datapath/RegisterFile/N23777 ,
         \DLX_Datapath/RegisterFile/N23776 ,
         \DLX_Datapath/RegisterFile/N23775 ,
         \DLX_Datapath/RegisterFile/N23774 ,
         \DLX_Datapath/RegisterFile/N23773 ,
         \DLX_Datapath/RegisterFile/N23772 ,
         \DLX_Datapath/RegisterFile/N23771 ,
         \DLX_Datapath/RegisterFile/N23770 ,
         \DLX_Datapath/RegisterFile/N23769 ,
         \DLX_Datapath/RegisterFile/N23768 ,
         \DLX_Datapath/RegisterFile/N23767 ,
         \DLX_Datapath/RegisterFile/N23766 ,
         \DLX_Datapath/RegisterFile/N23765 ,
         \DLX_Datapath/RegisterFile/N23764 ,
         \DLX_Datapath/RegisterFile/N23763 ,
         \DLX_Datapath/RegisterFile/N23762 ,
         \DLX_Datapath/RegisterFile/N23761 ,
         \DLX_Datapath/RegisterFile/N23760 ,
         \DLX_Datapath/RegisterFile/N23759 ,
         \DLX_Datapath/RegisterFile/N23758 ,
         \DLX_Datapath/RegisterFile/N23757 ,
         \DLX_Datapath/RegisterFile/N23756 ,
         \DLX_Datapath/RegisterFile/N23755 ,
         \DLX_Datapath/RegisterFile/N23754 ,
         \DLX_Datapath/RegisterFile/N23753 ,
         \DLX_Datapath/RegisterFile/N23750 ,
         \DLX_Datapath/RegisterFile/N23749 ,
         \DLX_Datapath/RegisterFile/N23748 ,
         \DLX_Datapath/RegisterFile/N23747 ,
         \DLX_Datapath/RegisterFile/N23746 ,
         \DLX_Datapath/RegisterFile/N23745 ,
         \DLX_Datapath/RegisterFile/N23744 ,
         \DLX_Datapath/RegisterFile/N23743 ,
         \DLX_Datapath/RegisterFile/N23742 ,
         \DLX_Datapath/RegisterFile/N23741 ,
         \DLX_Datapath/RegisterFile/N23740 ,
         \DLX_Datapath/RegisterFile/N23739 ,
         \DLX_Datapath/RegisterFile/N23735 ,
         \DLX_Datapath/RegisterFile/N23732 ,
         \DLX_Datapath/RegisterFile/N23731 ,
         \DLX_Datapath/RegisterFile/N23730 ,
         \DLX_Datapath/RegisterFile/N23729 ,
         \DLX_Datapath/RegisterFile/N23728 ,
         \DLX_Datapath/RegisterFile/N23727 ,
         \DLX_Datapath/RegisterFile/N23726 ,
         \DLX_Datapath/RegisterFile/N23725 ,
         \DLX_Datapath/RegisterFile/N23723 ,
         \DLX_Datapath/RegisterFile/N23722 ,
         \DLX_Datapath/RegisterFile/N23721 ,
         \DLX_Datapath/RegisterFile/N23720 ,
         \DLX_Datapath/RegisterFile/N23719 ,
         \DLX_Datapath/RegisterFile/N23718 ,
         \DLX_Datapath/RegisterFile/N23717 ,
         \DLX_Datapath/RegisterFile/N23716 ,
         \DLX_Datapath/RegisterFile/N23715 ,
         \DLX_Datapath/RegisterFile/N23714 ,
         \DLX_Datapath/RegisterFile/N23713 ,
         \DLX_Datapath/RegisterFile/N23712 ,
         \DLX_Datapath/RegisterFile/N23711 ,
         \DLX_Datapath/RegisterFile/N23710 ,
         \DLX_Datapath/RegisterFile/N23709 ,
         \DLX_Datapath/RegisterFile/N23708 ,
         \DLX_Datapath/RegisterFile/N23707 ,
         \DLX_Datapath/RegisterFile/N23706 ,
         \DLX_Datapath/RegisterFile/N23705 ,
         \DLX_Datapath/RegisterFile/N23704 ,
         \DLX_Datapath/RegisterFile/N23703 ,
         \DLX_Datapath/RegisterFile/N23702 ,
         \DLX_Datapath/RegisterFile/N23701 ,
         \DLX_Datapath/RegisterFile/N23700 ,
         \DLX_Datapath/RegisterFile/N23699 ,
         \DLX_Datapath/RegisterFile/N23698 ,
         \DLX_Datapath/RegisterFile/N23697 ,
         \DLX_Datapath/RegisterFile/N23696 ,
         \DLX_Datapath/RegisterFile/N23695 ,
         \DLX_Datapath/RegisterFile/N23694 ,
         \DLX_Datapath/RegisterFile/N23693 ,
         \DLX_Datapath/RegisterFile/N23692 ,
         \DLX_Datapath/RegisterFile/N23691 ,
         \DLX_Datapath/RegisterFile/N23690 ,
         \DLX_Datapath/RegisterFile/N23689 ,
         \DLX_Datapath/RegisterFile/N23688 ,
         \DLX_Datapath/RegisterFile/N23687 ,
         \DLX_Datapath/RegisterFile/N23686 ,
         \DLX_Datapath/RegisterFile/N23685 ,
         \DLX_Datapath/RegisterFile/N23684 ,
         \DLX_Datapath/RegisterFile/N23683 ,
         \DLX_Datapath/RegisterFile/N23682 ,
         \DLX_Datapath/RegisterFile/N23681 ,
         \DLX_Datapath/RegisterFile/N23680 ,
         \DLX_Datapath/RegisterFile/N23679 ,
         \DLX_Datapath/RegisterFile/N23678 ,
         \DLX_Datapath/RegisterFile/N23677 ,
         \DLX_Datapath/RegisterFile/N23676 ,
         \DLX_Datapath/RegisterFile/N23675 ,
         \DLX_Datapath/RegisterFile/N23674 ,
         \DLX_Datapath/RegisterFile/N23673 ,
         \DLX_Datapath/RegisterFile/N23672 ,
         \DLX_Datapath/RegisterFile/N23671 ,
         \DLX_Datapath/RegisterFile/N23670 ,
         \DLX_Datapath/RegisterFile/N23669 ,
         \DLX_Datapath/RegisterFile/N23668 ,
         \DLX_Datapath/RegisterFile/N23667 ,
         \DLX_Datapath/RegisterFile/N23666 ,
         \DLX_Datapath/RegisterFile/N23665 ,
         \DLX_Datapath/RegisterFile/N23664 ,
         \DLX_Datapath/RegisterFile/N23663 ,
         \DLX_Datapath/RegisterFile/N23662 ,
         \DLX_Datapath/RegisterFile/N23661 ,
         \DLX_Datapath/RegisterFile/N23660 ,
         \DLX_Datapath/RegisterFile/N23659 ,
         \DLX_Datapath/RegisterFile/N23658 ,
         \DLX_Datapath/RegisterFile/N23657 ,
         \DLX_Datapath/RegisterFile/N23656 ,
         \DLX_Datapath/RegisterFile/N23655 ,
         \DLX_Datapath/RegisterFile/N23654 ,
         \DLX_Datapath/RegisterFile/N23653 ,
         \DLX_Datapath/RegisterFile/N23652 ,
         \DLX_Datapath/RegisterFile/N23651 ,
         \DLX_Datapath/RegisterFile/N23650 ,
         \DLX_Datapath/RegisterFile/N23649 ,
         \DLX_Datapath/RegisterFile/N23648 ,
         \DLX_Datapath/RegisterFile/N23647 ,
         \DLX_Datapath/RegisterFile/N23646 ,
         \DLX_Datapath/RegisterFile/N23645 ,
         \DLX_Datapath/RegisterFile/N23644 ,
         \DLX_Datapath/RegisterFile/N23643 ,
         \DLX_Datapath/RegisterFile/N23642 ,
         \DLX_Datapath/RegisterFile/N23641 ,
         \DLX_Datapath/RegisterFile/N23640 ,
         \DLX_Datapath/RegisterFile/N23639 ,
         \DLX_Datapath/RegisterFile/N23638 ,
         \DLX_Datapath/RegisterFile/N23637 ,
         \DLX_Datapath/RegisterFile/N23636 ,
         \DLX_Datapath/RegisterFile/N23635 ,
         \DLX_Datapath/RegisterFile/N23634 ,
         \DLX_Datapath/RegisterFile/N23633 ,
         \DLX_Datapath/RegisterFile/N23632 ,
         \DLX_Datapath/RegisterFile/N23631 ,
         \DLX_Datapath/RegisterFile/N23630 ,
         \DLX_Datapath/RegisterFile/N23629 ,
         \DLX_Datapath/RegisterFile/N23628 ,
         \DLX_Datapath/RegisterFile/N23627 ,
         \DLX_Datapath/RegisterFile/N23626 ,
         \DLX_Datapath/RegisterFile/N23625 ,
         \DLX_Datapath/RegisterFile/N23624 ,
         \DLX_Datapath/RegisterFile/N23623 ,
         \DLX_Datapath/RegisterFile/N23622 ,
         \DLX_Datapath/RegisterFile/N23621 ,
         \DLX_Datapath/RegisterFile/N23620 ,
         \DLX_Datapath/RegisterFile/N23619 ,
         \DLX_Datapath/RegisterFile/N23618 ,
         \DLX_Datapath/RegisterFile/N23617 ,
         \DLX_Datapath/RegisterFile/N23615 ,
         \DLX_Datapath/RegisterFile/N23614 ,
         \DLX_Datapath/RegisterFile/N23613 ,
         \DLX_Datapath/RegisterFile/N23612 ,
         \DLX_Datapath/RegisterFile/N23611 ,
         \DLX_Datapath/RegisterFile/N23610 ,
         \DLX_Datapath/RegisterFile/N23609 ,
         \DLX_Datapath/RegisterFile/N23608 ,
         \DLX_Datapath/RegisterFile/N23607 ,
         \DLX_Datapath/RegisterFile/N23606 ,
         \DLX_Datapath/RegisterFile/N23605 ,
         \DLX_Datapath/RegisterFile/N23604 ,
         \DLX_Datapath/RegisterFile/N23603 ,
         \DLX_Datapath/RegisterFile/N23602 ,
         \DLX_Datapath/RegisterFile/N23601 ,
         \DLX_Datapath/RegisterFile/N23600 ,
         \DLX_Datapath/RegisterFile/N23599 ,
         \DLX_Datapath/RegisterFile/N23598 ,
         \DLX_Datapath/RegisterFile/N23597 ,
         \DLX_Datapath/RegisterFile/N23596 ,
         \DLX_Datapath/RegisterFile/N23595 ,
         \DLX_Datapath/RegisterFile/N23594 ,
         \DLX_Datapath/RegisterFile/N23593 ,
         \DLX_Datapath/RegisterFile/N23592 ,
         \DLX_Datapath/RegisterFile/N23591 ,
         \DLX_Datapath/RegisterFile/N23590 ,
         \DLX_Datapath/RegisterFile/N23589 ,
         \DLX_Datapath/RegisterFile/N23588 ,
         \DLX_Datapath/RegisterFile/N23587 ,
         \DLX_Datapath/RegisterFile/N23586 ,
         \DLX_Datapath/RegisterFile/N23585 ,
         \DLX_Datapath/RegisterFile/N23584 ,
         \DLX_Datapath/RegisterFile/N23583 ,
         \DLX_Datapath/RegisterFile/N23582 ,
         \DLX_Datapath/RegisterFile/N23581 ,
         \DLX_Datapath/RegisterFile/N23580 ,
         \DLX_Datapath/RegisterFile/N23579 ,
         \DLX_Datapath/RegisterFile/N23578 ,
         \DLX_Datapath/RegisterFile/N23577 ,
         \DLX_Datapath/RegisterFile/N23576 ,
         \DLX_Datapath/RegisterFile/N23575 ,
         \DLX_Datapath/RegisterFile/N23574 ,
         \DLX_Datapath/RegisterFile/N23573 ,
         \DLX_Datapath/RegisterFile/N23572 ,
         \DLX_Datapath/RegisterFile/N23571 ,
         \DLX_Datapath/RegisterFile/N23570 ,
         \DLX_Datapath/RegisterFile/N23569 ,
         \DLX_Datapath/RegisterFile/N23568 ,
         \DLX_Datapath/RegisterFile/N23567 ,
         \DLX_Datapath/RegisterFile/N23566 ,
         \DLX_Datapath/RegisterFile/N23565 ,
         \DLX_Datapath/RegisterFile/N23564 ,
         \DLX_Datapath/RegisterFile/N23563 ,
         \DLX_Datapath/RegisterFile/N23561 ,
         \DLX_Datapath/RegisterFile/N23560 ,
         \DLX_Datapath/RegisterFile/N23558 ,
         \DLX_Datapath/RegisterFile/N23557 ,
         \DLX_Datapath/RegisterFile/N23556 ,
         \DLX_Datapath/RegisterFile/N23555 ,
         \DLX_Datapath/RegisterFile/N23554 ,
         \DLX_Datapath/RegisterFile/N23553 ,
         \DLX_Datapath/RegisterFile/N23552 ,
         \DLX_Datapath/RegisterFile/N23551 ,
         \DLX_Datapath/RegisterFile/N23550 ,
         \DLX_Datapath/RegisterFile/N23549 ,
         \DLX_Datapath/RegisterFile/N23548 ,
         \DLX_Datapath/RegisterFile/N23547 ,
         \DLX_Datapath/RegisterFile/N23543 ,
         \DLX_Datapath/RegisterFile/N23542 ,
         \DLX_Datapath/RegisterFile/N23539 ,
         \DLX_Datapath/RegisterFile/N23538 ,
         \DLX_Datapath/RegisterFile/N23536 ,
         \DLX_Datapath/RegisterFile/N23535 ,
         \DLX_Datapath/RegisterFile/N23534 ,
         \DLX_Datapath/RegisterFile/N23533 ,
         \DLX_Datapath/RegisterFile/N23531 ,
         \DLX_Datapath/RegisterFile/N23530 ,
         \DLX_Datapath/RegisterFile/N23529 ,
         \DLX_Datapath/RegisterFile/N23528 ,
         \DLX_Datapath/RegisterFile/N23527 ,
         \DLX_Datapath/RegisterFile/N23526 ,
         \DLX_Datapath/RegisterFile/N23525 ,
         \DLX_Datapath/RegisterFile/N23524 ,
         \DLX_Datapath/RegisterFile/N23523 ,
         \DLX_Datapath/RegisterFile/N23522 ,
         \DLX_Datapath/RegisterFile/N23521 ,
         \DLX_Datapath/RegisterFile/N23520 ,
         \DLX_Datapath/RegisterFile/N23519 ,
         \DLX_Datapath/RegisterFile/N23518 ,
         \DLX_Datapath/RegisterFile/N23517 ,
         \DLX_Datapath/RegisterFile/N23516 ,
         \DLX_Datapath/RegisterFile/N23515 ,
         \DLX_Datapath/RegisterFile/N23514 ,
         \DLX_Datapath/RegisterFile/N23513 ,
         \DLX_Datapath/RegisterFile/N23512 ,
         \DLX_Datapath/RegisterFile/N23511 ,
         \DLX_Datapath/RegisterFile/N23510 ,
         \DLX_Datapath/RegisterFile/N23509 ,
         \DLX_Datapath/RegisterFile/N23508 ,
         \DLX_Datapath/RegisterFile/N23507 ,
         \DLX_Datapath/RegisterFile/N23506 ,
         \DLX_Datapath/RegisterFile/N23505 ,
         \DLX_Datapath/RegisterFile/N23504 ,
         \DLX_Datapath/RegisterFile/N23503 ,
         \DLX_Datapath/RegisterFile/N23502 ,
         \DLX_Datapath/RegisterFile/N23501 ,
         \DLX_Datapath/RegisterFile/N23500 ,
         \DLX_Datapath/RegisterFile/N23499 ,
         \DLX_Datapath/RegisterFile/N23498 ,
         \DLX_Datapath/RegisterFile/N23497 ,
         \DLX_Datapath/RegisterFile/N23496 ,
         \DLX_Datapath/RegisterFile/N23494 ,
         \DLX_Datapath/RegisterFile/N23492 ,
         \DLX_Datapath/RegisterFile/N23491 ,
         \DLX_Datapath/RegisterFile/N23489 ,
         \DLX_Datapath/RegisterFile/N23486 ,
         \DLX_Datapath/RegisterFile/N23479 ,
         \DLX_Datapath/RegisterFile/N23476 ,
         \DLX_Datapath/RegisterFile/N23474 ,
         \DLX_Datapath/RegisterFile/N23473 ,
         \DLX_Datapath/RegisterFile/N23472 ,
         \DLX_Datapath/RegisterFile/N23471 ,
         \DLX_Datapath/RegisterFile/N23469 ,
         \DLX_Datapath/RegisterFile/N23467 ,
         \DLX_Datapath/RegisterFile/N23466 ,
         \DLX_Datapath/RegisterFile/N23465 ,
         \DLX_Datapath/RegisterFile/N23464 ,
         \DLX_Datapath/RegisterFile/N23463 ,
         \DLX_Datapath/RegisterFile/N23462 ,
         \DLX_Datapath/RegisterFile/N23461 ,
         \DLX_Datapath/RegisterFile/N23460 ,
         \DLX_Datapath/RegisterFile/N23459 ,
         \DLX_Datapath/RegisterFile/N23458 ,
         \DLX_Datapath/RegisterFile/N23457 ,
         \DLX_Datapath/RegisterFile/N23456 ,
         \DLX_Datapath/RegisterFile/N23455 ,
         \DLX_Datapath/RegisterFile/N23454 ,
         \DLX_Datapath/RegisterFile/N23453 ,
         \DLX_Datapath/RegisterFile/N23452 ,
         \DLX_Datapath/RegisterFile/N23451 ,
         \DLX_Datapath/RegisterFile/N23450 ,
         \DLX_Datapath/RegisterFile/N23449 ,
         \DLX_Datapath/RegisterFile/N23448 ,
         \DLX_Datapath/RegisterFile/N23447 ,
         \DLX_Datapath/RegisterFile/N23446 ,
         \DLX_Datapath/RegisterFile/N23445 ,
         \DLX_Datapath/RegisterFile/N23444 ,
         \DLX_Datapath/RegisterFile/N23443 ,
         \DLX_Datapath/RegisterFile/N23442 ,
         \DLX_Datapath/RegisterFile/N23441 ,
         \DLX_Datapath/RegisterFile/N23440 ,
         \DLX_Datapath/RegisterFile/N23439 ,
         \DLX_Datapath/RegisterFile/N23438 ,
         \DLX_Datapath/RegisterFile/N23437 ,
         \DLX_Datapath/RegisterFile/N23436 ,
         \DLX_Datapath/RegisterFile/N23435 ,
         \DLX_Datapath/RegisterFile/N23434 ,
         \DLX_Datapath/RegisterFile/N23433 ,
         \DLX_Datapath/RegisterFile/N23432 ,
         \DLX_Datapath/RegisterFile/N23431 ,
         \DLX_Datapath/RegisterFile/N23430 ,
         \DLX_Datapath/RegisterFile/N23429 ,
         \DLX_Datapath/RegisterFile/N23428 ,
         \DLX_Datapath/RegisterFile/N23427 ,
         \DLX_Datapath/RegisterFile/N23426 ,
         \DLX_Datapath/RegisterFile/N23425 ,
         \DLX_Datapath/RegisterFile/N23424 ,
         \DLX_Datapath/RegisterFile/N23423 ,
         \DLX_Datapath/RegisterFile/N23422 ,
         \DLX_Datapath/RegisterFile/N23421 ,
         \DLX_Datapath/RegisterFile/N23420 ,
         \DLX_Datapath/RegisterFile/N23419 ,
         \DLX_Datapath/RegisterFile/N23418 ,
         \DLX_Datapath/RegisterFile/N23417 ,
         \DLX_Datapath/RegisterFile/N23416 ,
         \DLX_Datapath/RegisterFile/N23415 ,
         \DLX_Datapath/RegisterFile/N23414 ,
         \DLX_Datapath/RegisterFile/N23413 ,
         \DLX_Datapath/RegisterFile/N23412 ,
         \DLX_Datapath/RegisterFile/N23411 ,
         \DLX_Datapath/RegisterFile/N23410 ,
         \DLX_Datapath/RegisterFile/N23409 ,
         \DLX_Datapath/RegisterFile/N23408 ,
         \DLX_Datapath/RegisterFile/N23407 ,
         \DLX_Datapath/RegisterFile/N23406 ,
         \DLX_Datapath/RegisterFile/N23405 ,
         \DLX_Datapath/RegisterFile/N23404 ,
         \DLX_Datapath/RegisterFile/N23403 ,
         \DLX_Datapath/RegisterFile/N23402 ,
         \DLX_Datapath/RegisterFile/N23401 ,
         \DLX_Datapath/RegisterFile/N23400 ,
         \DLX_Datapath/RegisterFile/N23399 ,
         \DLX_Datapath/RegisterFile/N23398 ,
         \DLX_Datapath/RegisterFile/N23397 ,
         \DLX_Datapath/RegisterFile/N23396 ,
         \DLX_Datapath/RegisterFile/N23395 ,
         \DLX_Datapath/RegisterFile/N23394 ,
         \DLX_Datapath/RegisterFile/N23393 ,
         \DLX_Datapath/RegisterFile/N23392 ,
         \DLX_Datapath/RegisterFile/N23391 ,
         \DLX_Datapath/RegisterFile/N23390 ,
         \DLX_Datapath/RegisterFile/N23389 ,
         \DLX_Datapath/RegisterFile/N23388 ,
         \DLX_Datapath/RegisterFile/N23387 ,
         \DLX_Datapath/RegisterFile/N23386 ,
         \DLX_Datapath/RegisterFile/N23385 ,
         \DLX_Datapath/RegisterFile/N23384 ,
         \DLX_Datapath/RegisterFile/N23383 ,
         \DLX_Datapath/RegisterFile/N23382 ,
         \DLX_Datapath/RegisterFile/N23381 ,
         \DLX_Datapath/RegisterFile/N23380 ,
         \DLX_Datapath/RegisterFile/N23379 ,
         \DLX_Datapath/RegisterFile/N23378 ,
         \DLX_Datapath/RegisterFile/N23377 ,
         \DLX_Datapath/RegisterFile/N23376 ,
         \DLX_Datapath/RegisterFile/N23375 ,
         \DLX_Datapath/RegisterFile/N23374 ,
         \DLX_Datapath/RegisterFile/N23373 ,
         \DLX_Datapath/RegisterFile/N23372 ,
         \DLX_Datapath/RegisterFile/N23371 ,
         \DLX_Datapath/RegisterFile/N23370 ,
         \DLX_Datapath/RegisterFile/N23369 ,
         \DLX_Datapath/RegisterFile/N23368 ,
         \DLX_Datapath/RegisterFile/N23367 ,
         \DLX_Datapath/RegisterFile/N23365 ,
         \DLX_Datapath/RegisterFile/N23364 ,
         \DLX_Datapath/RegisterFile/N23363 ,
         \DLX_Datapath/RegisterFile/N23361 ,
         \DLX_Datapath/RegisterFile/N23358 ,
         \DLX_Datapath/RegisterFile/N23356 ,
         \DLX_Datapath/RegisterFile/N23355 ,
         \DLX_Datapath/RegisterFile/N23351 ,
         \DLX_Datapath/RegisterFile/N23347 ,
         \DLX_Datapath/RegisterFile/N23346 ,
         \DLX_Datapath/RegisterFile/N23344 ,
         \DLX_Datapath/RegisterFile/N23343 ,
         \DLX_Datapath/RegisterFile/N23341 ,
         \DLX_Datapath/RegisterFile/N23339 ,
         \DLX_Datapath/RegisterFile/N23338 ,
         \DLX_Datapath/RegisterFile/N23337 ,
         \DLX_Datapath/RegisterFile/N23336 ,
         \DLX_Datapath/RegisterFile/N23335 ,
         \DLX_Datapath/RegisterFile/N23334 ,
         \DLX_Datapath/RegisterFile/N23333 ,
         \DLX_Datapath/RegisterFile/N23332 ,
         \DLX_Datapath/RegisterFile/N23331 ,
         \DLX_Datapath/RegisterFile/N23330 ,
         \DLX_Datapath/RegisterFile/N23329 ,
         \DLX_Datapath/RegisterFile/N23328 ,
         \DLX_Datapath/RegisterFile/N23327 ,
         \DLX_Datapath/RegisterFile/N23326 ,
         \DLX_Datapath/RegisterFile/N23325 ,
         \DLX_Datapath/RegisterFile/N23324 ,
         \DLX_Datapath/RegisterFile/N23323 ,
         \DLX_Datapath/RegisterFile/N23322 ,
         \DLX_Datapath/RegisterFile/N23321 ,
         \DLX_Datapath/RegisterFile/N23320 ,
         \DLX_Datapath/RegisterFile/N23319 ,
         \DLX_Datapath/RegisterFile/N23318 ,
         \DLX_Datapath/RegisterFile/N23317 ,
         \DLX_Datapath/RegisterFile/N23316 ,
         \DLX_Datapath/RegisterFile/N23315 ,
         \DLX_Datapath/RegisterFile/N23314 ,
         \DLX_Datapath/RegisterFile/N23313 ,
         \DLX_Datapath/RegisterFile/N23312 ,
         \DLX_Datapath/RegisterFile/N23311 ,
         \DLX_Datapath/RegisterFile/N23310 ,
         \DLX_Datapath/RegisterFile/N23309 ,
         \DLX_Datapath/RegisterFile/N23308 ,
         \DLX_Datapath/RegisterFile/N23307 ,
         \DLX_Datapath/RegisterFile/N23306 ,
         \DLX_Datapath/RegisterFile/N23305 ,
         \DLX_Datapath/RegisterFile/N23304 ,
         \DLX_Datapath/RegisterFile/N23303 ,
         \DLX_Datapath/RegisterFile/N23301 ,
         \DLX_Datapath/RegisterFile/N23299 ,
         \DLX_Datapath/RegisterFile/N23298 ,
         \DLX_Datapath/RegisterFile/N23297 ,
         \DLX_Datapath/RegisterFile/N23296 ,
         \DLX_Datapath/RegisterFile/N23295 ,
         \DLX_Datapath/RegisterFile/N23294 ,
         \DLX_Datapath/RegisterFile/N23293 ,
         \DLX_Datapath/RegisterFile/N23292 ,
         \DLX_Datapath/RegisterFile/N23291 ,
         \DLX_Datapath/RegisterFile/N23289 ,
         \DLX_Datapath/RegisterFile/N23287 ,
         \DLX_Datapath/RegisterFile/N23286 ,
         \DLX_Datapath/RegisterFile/N23284 ,
         \DLX_Datapath/RegisterFile/N23283 ,
         \DLX_Datapath/RegisterFile/N23282 ,
         \DLX_Datapath/RegisterFile/N23280 ,
         \DLX_Datapath/RegisterFile/N23279 ,
         \DLX_Datapath/RegisterFile/N23278 ,
         \DLX_Datapath/RegisterFile/N23277 ,
         \DLX_Datapath/RegisterFile/N23275 ,
         \DLX_Datapath/RegisterFile/N23274 ,
         \DLX_Datapath/RegisterFile/N23273 ,
         \DLX_Datapath/RegisterFile/N23272 ,
         \DLX_Datapath/RegisterFile/N23271 ,
         \DLX_Datapath/RegisterFile/N23270 ,
         \DLX_Datapath/RegisterFile/N23269 ,
         \DLX_Datapath/RegisterFile/N23268 ,
         \DLX_Datapath/RegisterFile/N23267 ,
         \DLX_Datapath/RegisterFile/N23266 ,
         \DLX_Datapath/RegisterFile/N23265 ,
         \DLX_Datapath/RegisterFile/N23264 ,
         \DLX_Datapath/RegisterFile/N23263 ,
         \DLX_Datapath/RegisterFile/N23262 ,
         \DLX_Datapath/RegisterFile/N23261 ,
         \DLX_Datapath/RegisterFile/N23260 ,
         \DLX_Datapath/RegisterFile/N23259 ,
         \DLX_Datapath/RegisterFile/N23258 ,
         \DLX_Datapath/RegisterFile/N23257 ,
         \DLX_Datapath/RegisterFile/N23256 ,
         \DLX_Datapath/RegisterFile/N23255 ,
         \DLX_Datapath/RegisterFile/N23254 ,
         \DLX_Datapath/RegisterFile/N23253 ,
         \DLX_Datapath/RegisterFile/N23252 ,
         \DLX_Datapath/RegisterFile/N23251 ,
         \DLX_Datapath/RegisterFile/N23250 ,
         \DLX_Datapath/RegisterFile/N23249 ,
         \DLX_Datapath/RegisterFile/N23248 ,
         \DLX_Datapath/RegisterFile/N23247 ,
         \DLX_Datapath/RegisterFile/N23246 ,
         \DLX_Datapath/RegisterFile/N23245 ,
         \DLX_Datapath/RegisterFile/N23244 ,
         \DLX_Datapath/RegisterFile/N23243 ,
         \DLX_Datapath/RegisterFile/N23242 ,
         \DLX_Datapath/RegisterFile/N23241 ,
         \DLX_Datapath/RegisterFile/N23240 ,
         \DLX_Datapath/RegisterFile/N23239 ,
         \DLX_Datapath/RegisterFile/N23238 ,
         \DLX_Datapath/RegisterFile/N23237 ,
         \DLX_Datapath/RegisterFile/N23236 ,
         \DLX_Datapath/RegisterFile/N23235 ,
         \DLX_Datapath/RegisterFile/N23234 ,
         \DLX_Datapath/RegisterFile/N23233 ,
         \DLX_Datapath/RegisterFile/N23232 ,
         \DLX_Datapath/RegisterFile/N23231 ,
         \DLX_Datapath/RegisterFile/N23230 ,
         \DLX_Datapath/RegisterFile/N23229 ,
         \DLX_Datapath/RegisterFile/N23228 ,
         \DLX_Datapath/RegisterFile/N23227 ,
         \DLX_Datapath/RegisterFile/N23226 ,
         \DLX_Datapath/RegisterFile/N23225 ,
         \DLX_Datapath/RegisterFile/N23224 ,
         \DLX_Datapath/RegisterFile/N23223 ,
         \DLX_Datapath/RegisterFile/N23222 ,
         \DLX_Datapath/RegisterFile/N23221 ,
         \DLX_Datapath/RegisterFile/N23220 ,
         \DLX_Datapath/RegisterFile/N23219 ,
         \DLX_Datapath/RegisterFile/N23218 ,
         \DLX_Datapath/RegisterFile/N23217 ,
         \DLX_Datapath/RegisterFile/N23216 ,
         \DLX_Datapath/RegisterFile/N23215 ,
         \DLX_Datapath/RegisterFile/N23214 ,
         \DLX_Datapath/RegisterFile/N23213 ,
         \DLX_Datapath/RegisterFile/N23212 ,
         \DLX_Datapath/RegisterFile/N23211 ,
         \DLX_Datapath/RegisterFile/N23210 ,
         \DLX_Datapath/RegisterFile/N23209 ,
         \DLX_Datapath/RegisterFile/N23208 ,
         \DLX_Datapath/RegisterFile/N23207 ,
         \DLX_Datapath/RegisterFile/N23206 ,
         \DLX_Datapath/RegisterFile/N23205 ,
         \DLX_Datapath/RegisterFile/N23204 ,
         \DLX_Datapath/RegisterFile/N23203 ,
         \DLX_Datapath/RegisterFile/N23202 ,
         \DLX_Datapath/RegisterFile/N23201 ,
         \DLX_Datapath/RegisterFile/N23200 ,
         \DLX_Datapath/RegisterFile/N23199 ,
         \DLX_Datapath/RegisterFile/N23198 ,
         \DLX_Datapath/RegisterFile/N23197 ,
         \DLX_Datapath/RegisterFile/N23196 ,
         \DLX_Datapath/RegisterFile/N23195 ,
         \DLX_Datapath/RegisterFile/N23194 ,
         \DLX_Datapath/RegisterFile/N23193 ,
         \DLX_Datapath/RegisterFile/N23192 ,
         \DLX_Datapath/RegisterFile/N23191 ,
         \DLX_Datapath/RegisterFile/N23190 ,
         \DLX_Datapath/RegisterFile/N23189 ,
         \DLX_Datapath/RegisterFile/N23188 ,
         \DLX_Datapath/RegisterFile/N23187 ,
         \DLX_Datapath/RegisterFile/N23186 ,
         \DLX_Datapath/RegisterFile/N23185 ,
         \DLX_Datapath/RegisterFile/N23184 ,
         \DLX_Datapath/RegisterFile/N23183 ,
         \DLX_Datapath/RegisterFile/N23182 ,
         \DLX_Datapath/RegisterFile/N23181 ,
         \DLX_Datapath/RegisterFile/N23180 ,
         \DLX_Datapath/RegisterFile/N23179 ,
         \DLX_Datapath/RegisterFile/N23178 ,
         \DLX_Datapath/RegisterFile/N23177 ,
         \DLX_Datapath/RegisterFile/N23176 ,
         \DLX_Datapath/RegisterFile/N23174 ,
         \DLX_Datapath/RegisterFile/N23173 ,
         \DLX_Datapath/RegisterFile/N23172 ,
         \DLX_Datapath/RegisterFile/N23171 ,
         \DLX_Datapath/RegisterFile/N23170 ,
         \DLX_Datapath/RegisterFile/N23169 ,
         \DLX_Datapath/RegisterFile/N23168 ,
         \DLX_Datapath/RegisterFile/N23167 ,
         \DLX_Datapath/RegisterFile/N23166 ,
         \DLX_Datapath/RegisterFile/N23165 ,
         \DLX_Datapath/RegisterFile/N23163 ,
         \DLX_Datapath/RegisterFile/N23162 ,
         \DLX_Datapath/RegisterFile/N23161 ,
         \DLX_Datapath/RegisterFile/N23160 ,
         \DLX_Datapath/RegisterFile/N23159 ,
         \DLX_Datapath/RegisterFile/N23158 ,
         \DLX_Datapath/RegisterFile/N23157 ,
         \DLX_Datapath/RegisterFile/N23156 ,
         \DLX_Datapath/RegisterFile/N23155 ,
         \DLX_Datapath/RegisterFile/N23154 ,
         \DLX_Datapath/RegisterFile/N23153 ,
         \DLX_Datapath/RegisterFile/N23152 ,
         \DLX_Datapath/RegisterFile/N23151 ,
         \DLX_Datapath/RegisterFile/N23150 ,
         \DLX_Datapath/RegisterFile/N23149 ,
         \DLX_Datapath/RegisterFile/N23148 ,
         \DLX_Datapath/RegisterFile/N23147 ,
         \DLX_Datapath/RegisterFile/N23146 ,
         \DLX_Datapath/RegisterFile/N23145 ,
         \DLX_Datapath/RegisterFile/N23144 ,
         \DLX_Datapath/RegisterFile/N23143 ,
         \DLX_Datapath/RegisterFile/N23142 ,
         \DLX_Datapath/RegisterFile/N23141 ,
         \DLX_Datapath/RegisterFile/N23140 ,
         \DLX_Datapath/RegisterFile/N23139 ,
         \DLX_Datapath/RegisterFile/N23138 ,
         \DLX_Datapath/RegisterFile/N23137 ,
         \DLX_Datapath/RegisterFile/N23136 ,
         \DLX_Datapath/RegisterFile/N23135 ,
         \DLX_Datapath/RegisterFile/N23134 ,
         \DLX_Datapath/RegisterFile/N23133 ,
         \DLX_Datapath/RegisterFile/N23132 ,
         \DLX_Datapath/RegisterFile/N23131 ,
         \DLX_Datapath/RegisterFile/N23130 ,
         \DLX_Datapath/RegisterFile/N23129 ,
         \DLX_Datapath/RegisterFile/N23128 ,
         \DLX_Datapath/RegisterFile/N23127 ,
         \DLX_Datapath/RegisterFile/N23126 ,
         \DLX_Datapath/RegisterFile/N23125 ,
         \DLX_Datapath/RegisterFile/N23124 ,
         \DLX_Datapath/RegisterFile/N23123 ,
         \DLX_Datapath/RegisterFile/N23122 ,
         \DLX_Datapath/RegisterFile/N23121 ,
         \DLX_Datapath/RegisterFile/N23120 ,
         \DLX_Datapath/RegisterFile/N23119 ,
         \DLX_Datapath/RegisterFile/N23118 ,
         \DLX_Datapath/RegisterFile/N23117 ,
         \DLX_Datapath/RegisterFile/N23116 ,
         \DLX_Datapath/RegisterFile/N23115 ,
         \DLX_Datapath/RegisterFile/N23114 ,
         \DLX_Datapath/RegisterFile/N23113 ,
         \DLX_Datapath/RegisterFile/N23112 ,
         \DLX_Datapath/RegisterFile/N23111 ,
         \DLX_Datapath/RegisterFile/N23110 ,
         \DLX_Datapath/RegisterFile/N23109 ,
         \DLX_Datapath/RegisterFile/N23108 ,
         \DLX_Datapath/RegisterFile/N23107 ,
         \DLX_Datapath/RegisterFile/N23106 ,
         \DLX_Datapath/RegisterFile/N23104 ,
         \DLX_Datapath/RegisterFile/N23102 ,
         \DLX_Datapath/RegisterFile/N23101 ,
         \DLX_Datapath/RegisterFile/N23100 ,
         \DLX_Datapath/RegisterFile/N23099 ,
         \DLX_Datapath/RegisterFile/N23098 ,
         \DLX_Datapath/RegisterFile/N23097 ,
         \DLX_Datapath/RegisterFile/N23095 ,
         \DLX_Datapath/RegisterFile/N23093 ,
         \DLX_Datapath/RegisterFile/N23092 ,
         \DLX_Datapath/RegisterFile/N23091 ,
         \DLX_Datapath/RegisterFile/N23090 ,
         \DLX_Datapath/RegisterFile/N23089 ,
         \DLX_Datapath/RegisterFile/N23088 ,
         \DLX_Datapath/RegisterFile/N23087 ,
         \DLX_Datapath/RegisterFile/N23086 ,
         \DLX_Datapath/RegisterFile/N23085 ,
         \DLX_Datapath/RegisterFile/N23084 ,
         \DLX_Datapath/RegisterFile/N23083 ,
         \DLX_Datapath/RegisterFile/N23082 ,
         \DLX_Datapath/RegisterFile/N23081 ,
         \DLX_Datapath/RegisterFile/N23080 ,
         \DLX_Datapath/RegisterFile/N23079 ,
         \DLX_Datapath/RegisterFile/N23078 ,
         \DLX_Datapath/RegisterFile/N23077 ,
         \DLX_Datapath/RegisterFile/N23076 ,
         \DLX_Datapath/RegisterFile/N23075 ,
         \DLX_Datapath/RegisterFile/N23074 ,
         \DLX_Datapath/RegisterFile/N23073 ,
         \DLX_Datapath/RegisterFile/N23072 ,
         \DLX_Datapath/RegisterFile/N23071 ,
         \DLX_Datapath/RegisterFile/N23070 ,
         \DLX_Datapath/RegisterFile/N23069 ,
         \DLX_Datapath/RegisterFile/N23068 ,
         \DLX_Datapath/RegisterFile/N23067 ,
         \DLX_Datapath/RegisterFile/N23066 ,
         \DLX_Datapath/RegisterFile/N23065 ,
         \DLX_Datapath/RegisterFile/N23064 ,
         \DLX_Datapath/RegisterFile/N23063 ,
         \DLX_Datapath/RegisterFile/N23062 ,
         \DLX_Datapath/RegisterFile/N23061 ,
         \DLX_Datapath/RegisterFile/N23060 ,
         \DLX_Datapath/RegisterFile/N23059 ,
         \DLX_Datapath/RegisterFile/N23058 ,
         \DLX_Datapath/RegisterFile/N23057 ,
         \DLX_Datapath/RegisterFile/N23056 ,
         \DLX_Datapath/RegisterFile/N23055 ,
         \DLX_Datapath/RegisterFile/N23054 ,
         \DLX_Datapath/RegisterFile/N23053 ,
         \DLX_Datapath/RegisterFile/N23052 ,
         \DLX_Datapath/RegisterFile/N23051 ,
         \DLX_Datapath/RegisterFile/N23050 ,
         \DLX_Datapath/RegisterFile/N23049 ,
         \DLX_Datapath/RegisterFile/N23048 ,
         \DLX_Datapath/RegisterFile/N23047 ,
         \DLX_Datapath/RegisterFile/N23046 ,
         \DLX_Datapath/RegisterFile/N23045 ,
         \DLX_Datapath/RegisterFile/N23043 ,
         \DLX_Datapath/RegisterFile/N23042 ,
         \DLX_Datapath/RegisterFile/N23041 ,
         \DLX_Datapath/RegisterFile/N23040 ,
         \DLX_Datapath/RegisterFile/N23039 ,
         \DLX_Datapath/RegisterFile/N23038 ,
         \DLX_Datapath/RegisterFile/N23037 ,
         \DLX_Datapath/RegisterFile/N23036 ,
         \DLX_Datapath/RegisterFile/N23035 ,
         \DLX_Datapath/RegisterFile/N23034 ,
         \DLX_Datapath/RegisterFile/N23033 ,
         \DLX_Datapath/RegisterFile/N23032 ,
         \DLX_Datapath/RegisterFile/N23031 ,
         \DLX_Datapath/RegisterFile/N23030 ,
         \DLX_Datapath/RegisterFile/N23029 ,
         \DLX_Datapath/RegisterFile/N23028 ,
         \DLX_Datapath/RegisterFile/N23027 ,
         \DLX_Datapath/RegisterFile/N23026 ,
         \DLX_Datapath/RegisterFile/N23024 ,
         \DLX_Datapath/RegisterFile/N23023 ,
         \DLX_Datapath/RegisterFile/N23022 ,
         \DLX_Datapath/RegisterFile/N23021 ,
         \DLX_Datapath/RegisterFile/N23020 ,
         \DLX_Datapath/RegisterFile/N23018 ,
         \DLX_Datapath/RegisterFile/N23017 ,
         \DLX_Datapath/RegisterFile/N23016 ,
         \DLX_Datapath/RegisterFile/N23015 ,
         \DLX_Datapath/RegisterFile/N23014 ,
         \DLX_Datapath/RegisterFile/N23013 ,
         \DLX_Datapath/RegisterFile/N23012 ,
         \DLX_Datapath/RegisterFile/N23011 ,
         \DLX_Datapath/RegisterFile/N23010 ,
         \DLX_Datapath/RegisterFile/N23009 ,
         \DLX_Datapath/RegisterFile/N23008 ,
         \DLX_Datapath/RegisterFile/N23007 ,
         \DLX_Datapath/RegisterFile/N23006 ,
         \DLX_Datapath/RegisterFile/N23005 ,
         \DLX_Datapath/RegisterFile/N23004 ,
         \DLX_Datapath/RegisterFile/N23003 ,
         \DLX_Datapath/RegisterFile/N23002 ,
         \DLX_Datapath/RegisterFile/N23001 ,
         \DLX_Datapath/RegisterFile/N23000 ,
         \DLX_Datapath/RegisterFile/N22999 ,
         \DLX_Datapath/RegisterFile/N22998 ,
         \DLX_Datapath/RegisterFile/N22997 ,
         \DLX_Datapath/RegisterFile/N22996 ,
         \DLX_Datapath/RegisterFile/N22995 ,
         \DLX_Datapath/RegisterFile/N22994 ,
         \DLX_Datapath/RegisterFile/N22993 ,
         \DLX_Datapath/RegisterFile/N22992 ,
         \DLX_Datapath/RegisterFile/N22991 ,
         \DLX_Datapath/RegisterFile/N22990 ,
         \DLX_Datapath/RegisterFile/N22989 ,
         \DLX_Datapath/RegisterFile/N22988 ,
         \DLX_Datapath/RegisterFile/N22987 ,
         \DLX_Datapath/RegisterFile/N22986 ,
         \DLX_Datapath/RegisterFile/N22985 ,
         \DLX_Datapath/RegisterFile/N22984 ,
         \DLX_Datapath/RegisterFile/N22983 ,
         \DLX_Datapath/RegisterFile/N22982 ,
         \DLX_Datapath/RegisterFile/N22981 ,
         \DLX_Datapath/RegisterFile/N22980 ,
         \DLX_Datapath/RegisterFile/N22979 ,
         \DLX_Datapath/RegisterFile/N22978 ,
         \DLX_Datapath/RegisterFile/N22977 ,
         \DLX_Datapath/RegisterFile/N22976 ,
         \DLX_Datapath/RegisterFile/N22974 ,
         \DLX_Datapath/RegisterFile/N22973 ,
         \DLX_Datapath/RegisterFile/N22972 ,
         \DLX_Datapath/RegisterFile/N22971 ,
         \DLX_Datapath/RegisterFile/N22969 ,
         \DLX_Datapath/RegisterFile/N22967 ,
         \DLX_Datapath/RegisterFile/N22966 ,
         \DLX_Datapath/RegisterFile/N22964 ,
         \DLX_Datapath/RegisterFile/N22963 ,
         \DLX_Datapath/RegisterFile/N22962 ,
         \DLX_Datapath/RegisterFile/N22961 ,
         \DLX_Datapath/RegisterFile/N22960 ,
         \DLX_Datapath/RegisterFile/N22959 ,
         \DLX_Datapath/RegisterFile/N22958 ,
         \DLX_Datapath/RegisterFile/N22957 ,
         \DLX_Datapath/RegisterFile/N22954 ,
         \DLX_Datapath/RegisterFile/N22953 ,
         \DLX_Datapath/RegisterFile/N22952 ,
         \DLX_Datapath/RegisterFile/N22951 ,
         \DLX_Datapath/RegisterFile/N22950 ,
         \DLX_Datapath/RegisterFile/N22949 ,
         \DLX_Datapath/RegisterFile/N22948 ,
         \DLX_Datapath/RegisterFile/N22947 ,
         \DLX_Datapath/RegisterFile/N22946 ,
         \DLX_Datapath/RegisterFile/N22945 ,
         \DLX_Datapath/RegisterFile/N22944 ,
         \DLX_Datapath/RegisterFile/N22943 ,
         \DLX_Datapath/RegisterFile/N22942 ,
         \DLX_Datapath/RegisterFile/N22941 ,
         \DLX_Datapath/RegisterFile/N22940 ,
         \DLX_Datapath/RegisterFile/N22939 ,
         \DLX_Datapath/RegisterFile/N22938 ,
         \DLX_Datapath/RegisterFile/N22937 ,
         \DLX_Datapath/RegisterFile/N22936 ,
         \DLX_Datapath/RegisterFile/N22935 ,
         \DLX_Datapath/RegisterFile/N22934 ,
         \DLX_Datapath/RegisterFile/N22933 ,
         \DLX_Datapath/RegisterFile/N22932 ,
         \DLX_Datapath/RegisterFile/N22931 ,
         \DLX_Datapath/RegisterFile/N22930 ,
         \DLX_Datapath/RegisterFile/N22929 ,
         \DLX_Datapath/RegisterFile/N22928 ,
         \DLX_Datapath/RegisterFile/N22927 ,
         \DLX_Datapath/RegisterFile/N22926 ,
         \DLX_Datapath/RegisterFile/N22925 ,
         \DLX_Datapath/RegisterFile/N22924 ,
         \DLX_Datapath/RegisterFile/N22923 ,
         \DLX_Datapath/RegisterFile/N22922 ,
         \DLX_Datapath/RegisterFile/N22921 ,
         \DLX_Datapath/RegisterFile/N22920 ,
         \DLX_Datapath/RegisterFile/N22919 ,
         \DLX_Datapath/RegisterFile/N22918 ,
         \DLX_Datapath/RegisterFile/N22917 ,
         \DLX_Datapath/RegisterFile/N22916 ,
         \DLX_Datapath/RegisterFile/N22915 ,
         \DLX_Datapath/RegisterFile/N22914 ,
         \DLX_Datapath/RegisterFile/N22913 ,
         \DLX_Datapath/RegisterFile/N22912 ,
         \DLX_Datapath/RegisterFile/N22911 ,
         \DLX_Datapath/RegisterFile/N22910 ,
         \DLX_Datapath/RegisterFile/N22909 ,
         \DLX_Datapath/RegisterFile/N22908 ,
         \DLX_Datapath/RegisterFile/N22907 ,
         \DLX_Datapath/RegisterFile/N22905 ,
         \DLX_Datapath/RegisterFile/N22903 ,
         \DLX_Datapath/RegisterFile/N22902 ,
         \DLX_Datapath/RegisterFile/N22900 ,
         \DLX_Datapath/RegisterFile/N22899 ,
         \DLX_Datapath/RegisterFile/N22898 ,
         \DLX_Datapath/RegisterFile/N22896 ,
         \DLX_Datapath/RegisterFile/N22895 ,
         \DLX_Datapath/RegisterFile/N22894 ,
         \DLX_Datapath/RegisterFile/N22893 ,
         \DLX_Datapath/RegisterFile/N22890 ,
         \DLX_Datapath/RegisterFile/N22889 ,
         \DLX_Datapath/RegisterFile/N22888 ,
         \DLX_Datapath/RegisterFile/N22887 ,
         \DLX_Datapath/RegisterFile/N22886 ,
         \DLX_Datapath/RegisterFile/N22885 ,
         \DLX_Datapath/RegisterFile/N22884 ,
         \DLX_Datapath/RegisterFile/N22883 ,
         \DLX_Datapath/RegisterFile/N22882 ,
         \DLX_Datapath/RegisterFile/N22881 ,
         \DLX_Datapath/RegisterFile/N22880 ,
         \DLX_Datapath/RegisterFile/N22879 ,
         \DLX_Datapath/RegisterFile/N22878 ,
         \DLX_Datapath/RegisterFile/N22877 ,
         \DLX_Datapath/RegisterFile/N22876 ,
         \DLX_Datapath/RegisterFile/N22875 ,
         \DLX_Datapath/RegisterFile/N22874 ,
         \DLX_Datapath/RegisterFile/N22873 ,
         \DLX_Datapath/RegisterFile/N22872 ,
         \DLX_Datapath/RegisterFile/N22871 ,
         \DLX_Datapath/RegisterFile/N22870 ,
         \DLX_Datapath/RegisterFile/N22869 ,
         \DLX_Datapath/RegisterFile/N22868 ,
         \DLX_Datapath/RegisterFile/N22867 ,
         \DLX_Datapath/RegisterFile/N22866 ,
         \DLX_Datapath/RegisterFile/N22865 ,
         \DLX_Datapath/RegisterFile/N22864 ,
         \DLX_Datapath/RegisterFile/N22863 ,
         \DLX_Datapath/RegisterFile/N22862 ,
         \DLX_Datapath/RegisterFile/N22861 ,
         \DLX_Datapath/RegisterFile/N22860 ,
         \DLX_Datapath/RegisterFile/N22859 ,
         \DLX_Datapath/RegisterFile/N22858 ,
         \DLX_Datapath/RegisterFile/N22857 ,
         \DLX_Datapath/RegisterFile/N22856 ,
         \DLX_Datapath/RegisterFile/N22855 ,
         \DLX_Datapath/RegisterFile/N22854 ,
         \DLX_Datapath/RegisterFile/N22853 ,
         \DLX_Datapath/RegisterFile/N22852 ,
         \DLX_Datapath/RegisterFile/N22851 ,
         \DLX_Datapath/RegisterFile/N22850 ,
         \DLX_Datapath/RegisterFile/N22849 ,
         \DLX_Datapath/RegisterFile/N22848 ,
         \DLX_Datapath/RegisterFile/N22847 ,
         \DLX_Datapath/RegisterFile/N22846 ,
         \DLX_Datapath/RegisterFile/N22845 ,
         \DLX_Datapath/RegisterFile/N22844 ,
         \DLX_Datapath/RegisterFile/N22843 ,
         \DLX_Datapath/RegisterFile/N22842 ,
         \DLX_Datapath/RegisterFile/N22841 ,
         \DLX_Datapath/RegisterFile/N22840 ,
         \DLX_Datapath/RegisterFile/N22839 ,
         \DLX_Datapath/RegisterFile/N22838 ,
         \DLX_Datapath/RegisterFile/N22837 ,
         \DLX_Datapath/RegisterFile/N22836 ,
         \DLX_Datapath/RegisterFile/N22835 ,
         \DLX_Datapath/RegisterFile/N22834 ,
         \DLX_Datapath/RegisterFile/N22833 ,
         \DLX_Datapath/RegisterFile/N22832 ,
         \DLX_Datapath/RegisterFile/N22831 ,
         \DLX_Datapath/RegisterFile/N22830 ,
         \DLX_Datapath/RegisterFile/N22829 ,
         \DLX_Datapath/RegisterFile/N22828 ,
         \DLX_Datapath/RegisterFile/N22827 ,
         \DLX_Datapath/RegisterFile/N22826 ,
         \DLX_Datapath/RegisterFile/N22825 ,
         \DLX_Datapath/RegisterFile/N22824 ,
         \DLX_Datapath/RegisterFile/N22823 ,
         \DLX_Datapath/RegisterFile/N22822 ,
         \DLX_Datapath/RegisterFile/N22821 ,
         \DLX_Datapath/RegisterFile/N22820 ,
         \DLX_Datapath/RegisterFile/N22819 ,
         \DLX_Datapath/RegisterFile/N22818 ,
         \DLX_Datapath/RegisterFile/N22817 ,
         \DLX_Datapath/RegisterFile/N22816 ,
         \DLX_Datapath/RegisterFile/N22815 ,
         \DLX_Datapath/RegisterFile/N22814 ,
         \DLX_Datapath/RegisterFile/N22813 ,
         \DLX_Datapath/RegisterFile/N22812 ,
         \DLX_Datapath/RegisterFile/N22811 ,
         \DLX_Datapath/RegisterFile/N22810 ,
         \DLX_Datapath/RegisterFile/N22809 ,
         \DLX_Datapath/RegisterFile/N22808 ,
         \DLX_Datapath/RegisterFile/N22807 ,
         \DLX_Datapath/RegisterFile/N22806 ,
         \DLX_Datapath/RegisterFile/N22805 ,
         \DLX_Datapath/RegisterFile/N22804 ,
         \DLX_Datapath/RegisterFile/N22803 ,
         \DLX_Datapath/RegisterFile/N22802 ,
         \DLX_Datapath/RegisterFile/N22801 ,
         \DLX_Datapath/RegisterFile/N22800 ,
         \DLX_Datapath/RegisterFile/N22799 ,
         \DLX_Datapath/RegisterFile/N22798 ,
         \DLX_Datapath/RegisterFile/N22797 ,
         \DLX_Datapath/RegisterFile/N22796 ,
         \DLX_Datapath/RegisterFile/N22795 ,
         \DLX_Datapath/RegisterFile/N22794 ,
         \DLX_Datapath/RegisterFile/N22793 ,
         \DLX_Datapath/RegisterFile/N22792 ,
         \DLX_Datapath/RegisterFile/N22791 ,
         \DLX_Datapath/RegisterFile/N22790 ,
         \DLX_Datapath/RegisterFile/N22789 ,
         \DLX_Datapath/RegisterFile/N22788 ,
         \DLX_Datapath/RegisterFile/N22787 ,
         \DLX_Datapath/RegisterFile/N22786 ,
         \DLX_Datapath/RegisterFile/N22785 ,
         \DLX_Datapath/RegisterFile/N22784 ,
         \DLX_Datapath/RegisterFile/N22783 ,
         \DLX_Datapath/RegisterFile/N22782 ,
         \DLX_Datapath/RegisterFile/N22781 ,
         \DLX_Datapath/RegisterFile/N22780 ,
         \DLX_Datapath/RegisterFile/N22779 ,
         \DLX_Datapath/RegisterFile/N22778 ,
         \DLX_Datapath/RegisterFile/N22777 ,
         \DLX_Datapath/RegisterFile/N22776 ,
         \DLX_Datapath/RegisterFile/N22775 ,
         \DLX_Datapath/RegisterFile/N22774 ,
         \DLX_Datapath/RegisterFile/N22773 ,
         \DLX_Datapath/RegisterFile/N22772 ,
         \DLX_Datapath/RegisterFile/N22771 ,
         \DLX_Datapath/RegisterFile/N22770 ,
         \DLX_Datapath/RegisterFile/N22769 ,
         \DLX_Datapath/RegisterFile/N22768 ,
         \DLX_Datapath/RegisterFile/N22767 ,
         \DLX_Datapath/RegisterFile/N22766 ,
         \DLX_Datapath/RegisterFile/N22765 ,
         \DLX_Datapath/RegisterFile/N22764 ,
         \DLX_Datapath/RegisterFile/N22763 ,
         \DLX_Datapath/RegisterFile/N22762 ,
         \DLX_Datapath/RegisterFile/N22761 ,
         \DLX_Datapath/RegisterFile/N22760 ,
         \DLX_Datapath/RegisterFile/N22759 ,
         \DLX_Datapath/RegisterFile/N22758 ,
         \DLX_Datapath/RegisterFile/N22757 ,
         \DLX_Datapath/RegisterFile/N22756 ,
         \DLX_Datapath/RegisterFile/N22755 ,
         \DLX_Datapath/RegisterFile/N22754 ,
         \DLX_Datapath/RegisterFile/N22753 ,
         \DLX_Datapath/RegisterFile/N22752 ,
         \DLX_Datapath/RegisterFile/N22751 ,
         \DLX_Datapath/RegisterFile/N22750 ,
         \DLX_Datapath/RegisterFile/N22749 ,
         \DLX_Datapath/RegisterFile/N22748 ,
         \DLX_Datapath/RegisterFile/N22747 ,
         \DLX_Datapath/RegisterFile/N22746 ,
         \DLX_Datapath/RegisterFile/N22745 ,
         \DLX_Datapath/RegisterFile/N22744 ,
         \DLX_Datapath/RegisterFile/N22743 ,
         \DLX_Datapath/RegisterFile/N22742 ,
         \DLX_Datapath/RegisterFile/N22741 ,
         \DLX_Datapath/RegisterFile/N22740 ,
         \DLX_Datapath/RegisterFile/N22739 ,
         \DLX_Datapath/RegisterFile/N22738 ,
         \DLX_Datapath/RegisterFile/N22737 ,
         \DLX_Datapath/RegisterFile/N22736 ,
         \DLX_Datapath/RegisterFile/N22735 ,
         \DLX_Datapath/RegisterFile/N22734 ,
         \DLX_Datapath/RegisterFile/N22733 ,
         \DLX_Datapath/RegisterFile/N22732 ,
         \DLX_Datapath/RegisterFile/N22731 ,
         \DLX_Datapath/RegisterFile/N22730 ,
         \DLX_Datapath/RegisterFile/N22729 ,
         \DLX_Datapath/RegisterFile/N22728 ,
         \DLX_Datapath/RegisterFile/N22727 ,
         \DLX_Datapath/RegisterFile/N22726 ,
         \DLX_Datapath/RegisterFile/N22725 ,
         \DLX_Datapath/RegisterFile/N22724 ,
         \DLX_Datapath/RegisterFile/N22723 ,
         \DLX_Datapath/RegisterFile/N22722 ,
         \DLX_Datapath/RegisterFile/N22721 ,
         \DLX_Datapath/RegisterFile/N22720 ,
         \DLX_Datapath/RegisterFile/N22719 ,
         \DLX_Datapath/RegisterFile/N22718 ,
         \DLX_Datapath/RegisterFile/N22717 ,
         \DLX_Datapath/RegisterFile/N22716 ,
         \DLX_Datapath/RegisterFile/N22715 ,
         \DLX_Datapath/RegisterFile/N22714 ,
         \DLX_Datapath/RegisterFile/N22713 ,
         \DLX_Datapath/RegisterFile/N22712 ,
         \DLX_Datapath/RegisterFile/N22711 ,
         \DLX_Datapath/RegisterFile/N22710 ,
         \DLX_Datapath/RegisterFile/N22709 ,
         \DLX_Datapath/RegisterFile/N22708 ,
         \DLX_Datapath/RegisterFile/N22707 ,
         \DLX_Datapath/RegisterFile/N22706 ,
         \DLX_Datapath/RegisterFile/N22705 ,
         \DLX_Datapath/RegisterFile/N22704 ,
         \DLX_Datapath/RegisterFile/N22703 ,
         \DLX_Datapath/RegisterFile/N22702 ,
         \DLX_Datapath/RegisterFile/N22701 ,
         \DLX_Datapath/RegisterFile/N22700 ,
         \DLX_Datapath/RegisterFile/N22699 ,
         \DLX_Datapath/RegisterFile/N22698 ,
         \DLX_Datapath/RegisterFile/N22697 ,
         \DLX_Datapath/RegisterFile/N22696 ,
         \DLX_Datapath/RegisterFile/N22695 ,
         \DLX_Datapath/RegisterFile/N22694 ,
         \DLX_Datapath/RegisterFile/N22693 ,
         \DLX_Datapath/RegisterFile/N22692 ,
         \DLX_Datapath/RegisterFile/N22691 ,
         \DLX_Datapath/RegisterFile/N22690 ,
         \DLX_Datapath/RegisterFile/N22689 ,
         \DLX_Datapath/RegisterFile/N22688 ,
         \DLX_Datapath/RegisterFile/N22687 ,
         \DLX_Datapath/RegisterFile/N22686 ,
         \DLX_Datapath/RegisterFile/N22685 ,
         \DLX_Datapath/RegisterFile/N22684 ,
         \DLX_Datapath/RegisterFile/N22683 ,
         \DLX_Datapath/RegisterFile/N22682 ,
         \DLX_Datapath/RegisterFile/N22681 ,
         \DLX_Datapath/RegisterFile/N22680 ,
         \DLX_Datapath/RegisterFile/N22679 ,
         \DLX_Datapath/RegisterFile/N22678 ,
         \DLX_Datapath/RegisterFile/N22677 ,
         \DLX_Datapath/RegisterFile/N22676 ,
         \DLX_Datapath/RegisterFile/N22675 ,
         \DLX_Datapath/RegisterFile/N22674 ,
         \DLX_Datapath/RegisterFile/N22673 ,
         \DLX_Datapath/RegisterFile/N22672 ,
         \DLX_Datapath/RegisterFile/N22671 ,
         \DLX_Datapath/RegisterFile/N22670 ,
         \DLX_Datapath/RegisterFile/N22669 ,
         \DLX_Datapath/RegisterFile/N22668 ,
         \DLX_Datapath/RegisterFile/N22667 ,
         \DLX_Datapath/RegisterFile/N22666 ,
         \DLX_Datapath/RegisterFile/N22665 ,
         \DLX_Datapath/RegisterFile/N22664 ,
         \DLX_Datapath/RegisterFile/N22663 ,
         \DLX_Datapath/RegisterFile/N22662 ,
         \DLX_Datapath/RegisterFile/N22661 ,
         \DLX_Datapath/RegisterFile/N22660 ,
         \DLX_Datapath/RegisterFile/N22659 ,
         \DLX_Datapath/RegisterFile/N22657 ,
         \DLX_Datapath/RegisterFile/N22656 ,
         \DLX_Datapath/RegisterFile/N22655 ,
         \DLX_Datapath/RegisterFile/N22654 ,
         \DLX_Datapath/RegisterFile/N22653 ,
         \DLX_Datapath/RegisterFile/N22652 ,
         \DLX_Datapath/RegisterFile/N22651 ,
         \DLX_Datapath/RegisterFile/N22650 ,
         \DLX_Datapath/RegisterFile/N22649 ,
         \DLX_Datapath/RegisterFile/N22648 ,
         \DLX_Datapath/RegisterFile/N22647 ,
         \DLX_Datapath/RegisterFile/N22646 ,
         \DLX_Datapath/RegisterFile/N22645 ,
         \DLX_Datapath/RegisterFile/N22644 ,
         \DLX_Datapath/RegisterFile/N22643 ,
         \DLX_Datapath/RegisterFile/N22642 ,
         \DLX_Datapath/RegisterFile/N22641 ,
         \DLX_Datapath/RegisterFile/N22640 ,
         \DLX_Datapath/RegisterFile/N22639 ,
         \DLX_Datapath/RegisterFile/N22638 ,
         \DLX_Datapath/RegisterFile/N22637 ,
         \DLX_Datapath/RegisterFile/N22635 ,
         \DLX_Datapath/RegisterFile/N22634 ,
         \DLX_Datapath/RegisterFile/N22633 ,
         \DLX_Datapath/RegisterFile/N22632 ,
         \DLX_Datapath/RegisterFile/N22631 ,
         \DLX_Datapath/RegisterFile/N22630 ,
         \DLX_Datapath/RegisterFile/N22629 ,
         \DLX_Datapath/RegisterFile/N22628 ,
         \DLX_Datapath/RegisterFile/N22627 ,
         \DLX_Datapath/RegisterFile/N22626 ,
         \DLX_Datapath/RegisterFile/N22625 ,
         \DLX_Datapath/RegisterFile/N22624 ,
         \DLX_Datapath/RegisterFile/N22623 ,
         \DLX_Datapath/RegisterFile/N22622 ,
         \DLX_Datapath/RegisterFile/N22621 ,
         \DLX_Datapath/RegisterFile/N22620 ,
         \DLX_Datapath/RegisterFile/N22619 ,
         \DLX_Datapath/RegisterFile/N22618 ,
         \DLX_Datapath/RegisterFile/N22617 ,
         \DLX_Datapath/RegisterFile/N22616 ,
         \DLX_Datapath/RegisterFile/N22615 ,
         \DLX_Datapath/RegisterFile/N22614 ,
         \DLX_Datapath/RegisterFile/N22613 ,
         \DLX_Datapath/RegisterFile/N22612 ,
         \DLX_Datapath/RegisterFile/N22611 ,
         \DLX_Datapath/RegisterFile/N22610 ,
         \DLX_Datapath/RegisterFile/N22609 ,
         \DLX_Datapath/RegisterFile/N22608 ,
         \DLX_Datapath/RegisterFile/N22607 ,
         \DLX_Datapath/RegisterFile/N22606 ,
         \DLX_Datapath/RegisterFile/N22605 ,
         \DLX_Datapath/RegisterFile/N22604 ,
         \DLX_Datapath/RegisterFile/N22603 ,
         \DLX_Datapath/RegisterFile/N22602 ,
         \DLX_Datapath/RegisterFile/N22601 ,
         \DLX_Datapath/RegisterFile/N22600 ,
         \DLX_Datapath/RegisterFile/N22599 ,
         \DLX_Datapath/RegisterFile/N22598 ,
         \DLX_Datapath/RegisterFile/N22597 ,
         \DLX_Datapath/RegisterFile/N22596 ,
         \DLX_Datapath/RegisterFile/N22595 ,
         \DLX_Datapath/RegisterFile/N22594 ,
         \DLX_Datapath/RegisterFile/N22593 ,
         \DLX_Datapath/RegisterFile/N22592 ,
         \DLX_Datapath/RegisterFile/N22591 ,
         \DLX_Datapath/RegisterFile/N22590 ,
         \DLX_Datapath/RegisterFile/N22589 ,
         \DLX_Datapath/RegisterFile/N22588 ,
         \DLX_Datapath/RegisterFile/N22587 ,
         \DLX_Datapath/RegisterFile/N22586 ,
         \DLX_Datapath/RegisterFile/N22585 ,
         \DLX_Datapath/RegisterFile/N22584 ,
         \DLX_Datapath/RegisterFile/N22583 ,
         \DLX_Datapath/RegisterFile/N22582 ,
         \DLX_Datapath/RegisterFile/N22581 ,
         \DLX_Datapath/RegisterFile/N22580 ,
         \DLX_Datapath/RegisterFile/N22579 ,
         \DLX_Datapath/RegisterFile/N22577 ,
         \DLX_Datapath/RegisterFile/N22576 ,
         \DLX_Datapath/RegisterFile/N22575 ,
         \DLX_Datapath/RegisterFile/N22574 ,
         \DLX_Datapath/RegisterFile/N22572 ,
         \DLX_Datapath/RegisterFile/N22571 ,
         \DLX_Datapath/RegisterFile/N22570 ,
         \DLX_Datapath/RegisterFile/N22569 ,
         \DLX_Datapath/RegisterFile/N22568 ,
         \DLX_Datapath/RegisterFile/N22567 ,
         \DLX_Datapath/RegisterFile/N22566 ,
         \DLX_Datapath/RegisterFile/N22565 ,
         \DLX_Datapath/RegisterFile/N22564 ,
         \DLX_Datapath/RegisterFile/N22563 ,
         \DLX_Datapath/RegisterFile/N22562 ,
         \DLX_Datapath/RegisterFile/N22561 ,
         \DLX_Datapath/RegisterFile/N22560 ,
         \DLX_Datapath/RegisterFile/N22559 ,
         \DLX_Datapath/RegisterFile/N22558 ,
         \DLX_Datapath/RegisterFile/N22557 ,
         \DLX_Datapath/RegisterFile/N22556 ,
         \DLX_Datapath/RegisterFile/N22555 ,
         \DLX_Datapath/RegisterFile/N22554 ,
         \DLX_Datapath/RegisterFile/N22553 ,
         \DLX_Datapath/RegisterFile/N22552 ,
         \DLX_Datapath/RegisterFile/N22551 ,
         \DLX_Datapath/RegisterFile/N22550 ,
         \DLX_Datapath/RegisterFile/N22549 ,
         \DLX_Datapath/RegisterFile/N22548 ,
         \DLX_Datapath/RegisterFile/N22547 ,
         \DLX_Datapath/RegisterFile/N22545 ,
         \DLX_Datapath/RegisterFile/N22544 ,
         \DLX_Datapath/RegisterFile/N22543 ,
         \DLX_Datapath/RegisterFile/N22542 ,
         \DLX_Datapath/RegisterFile/N22541 ,
         \DLX_Datapath/RegisterFile/N22540 ,
         \DLX_Datapath/RegisterFile/N22539 , \DLX_Datapath/RegisterFile/N9337 ,
         \DLX_Datapath/RegisterFile/old_CWP2[1] ,
         \DLX_Datapath/RegisterFile/old_CWP2[2] ,
         \DLX_Datapath/ArithLogUnit/N193 , \DLX_Datapath/ArithLogUnit/N187 ,
         \DLX_Datapath/ArithLogUnit/N180 , \DLX_Datapath/ArithLogUnit/N179 ,
         \DLX_Datapath/ArithLogUnit/N178 , \DLX_Datapath/ArithLogUnit/N177 ,
         \DLX_Datapath/ArithLogUnit/N176 , \DLX_Datapath/ArithLogUnit/N175 ,
         \DLX_Datapath/ArithLogUnit/N174 , \DLX_Datapath/ArithLogUnit/N173 ,
         \DLX_Datapath/ArithLogUnit/N172 , \DLX_Datapath/ArithLogUnit/N171 ,
         \DLX_Datapath/ArithLogUnit/N170 , \DLX_Datapath/ArithLogUnit/N169 ,
         \DLX_Datapath/ArithLogUnit/N168 , \DLX_Datapath/ArithLogUnit/N167 ,
         \DLX_Datapath/ArithLogUnit/N166 , \DLX_Datapath/ArithLogUnit/N165 ,
         \DLX_Datapath/ArithLogUnit/N164 , \DLX_Datapath/ArithLogUnit/N163 ,
         \DLX_Datapath/ArithLogUnit/N162 , \DLX_Datapath/ArithLogUnit/N161 ,
         \DLX_Datapath/ArithLogUnit/N160 , \DLX_Datapath/ArithLogUnit/N159 ,
         \DLX_Datapath/ArithLogUnit/N158 , \DLX_Datapath/ArithLogUnit/N157 ,
         \DLX_Datapath/ArithLogUnit/N156 , \DLX_Datapath/ArithLogUnit/N155 ,
         \DLX_Datapath/ArithLogUnit/N154 , \DLX_Datapath/ArithLogUnit/N153 ,
         \DLX_Datapath/ArithLogUnit/N152 , \DLX_Datapath/ArithLogUnit/N151 ,
         \DLX_Datapath/ArithLogUnit/N150 , \DLX_Datapath/ArithLogUnit/N149 ,
         \DLX_Datapath/ArithLogUnit/N148 , \DLX_Datapath/ArithLogUnit/N147 ,
         \DLX_Datapath/ArithLogUnit/N146 , \DLX_Datapath/ArithLogUnit/N145 ,
         \DLX_Datapath/ArithLogUnit/N141 , \DLX_Datapath/ArithLogUnit/N140 ,
         \DLX_Datapath/ArithLogUnit/N139 , \DLX_Datapath/ArithLogUnit/N138 ,
         \DLX_Datapath/ArithLogUnit/N137 , \DLX_Datapath/ArithLogUnit/N136 ,
         \DLX_Datapath/ArithLogUnit/N135 , \DLX_Datapath/ArithLogUnit/N134 ,
         \DLX_Datapath/ArithLogUnit/N133 , \DLX_Datapath/ArithLogUnit/N132 ,
         \DLX_Datapath/ArithLogUnit/N131 , \DLX_Datapath/ArithLogUnit/N130 ,
         \DLX_Datapath/ArithLogUnit/N129 , \DLX_Datapath/ArithLogUnit/N128 ,
         \DLX_Datapath/ArithLogUnit/N127 , \DLX_Datapath/ArithLogUnit/N126 ,
         \DLX_Datapath/ArithLogUnit/N125 , \DLX_Datapath/ArithLogUnit/N124 ,
         \DLX_Datapath/ArithLogUnit/N123 , \DLX_Datapath/ArithLogUnit/N122 ,
         \DLX_Datapath/ArithLogUnit/N121 , \DLX_Datapath/ArithLogUnit/N120 ,
         \DLX_Datapath/ArithLogUnit/N119 , \DLX_Datapath/ArithLogUnit/N118 ,
         \DLX_Datapath/ArithLogUnit/N117 , \DLX_Datapath/ArithLogUnit/N116 ,
         \DLX_Datapath/ArithLogUnit/N115 , \DLX_Datapath/ArithLogUnit/N114 ,
         \DLX_Datapath/ArithLogUnit/N113 , \DLX_Datapath/ArithLogUnit/N112 ,
         \DLX_Datapath/ArithLogUnit/useBorrow_cmp ,
         \DLX_Datapath/ArithLogUnit/Cout_cmp ,
         \DLX_Datapath/ArithLogUnit/Cin_add ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[1] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[16] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[17] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[0] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[16] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[17] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ,
         \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N103 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N102 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N101 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N100 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N99 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N98 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N97 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N96 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N95 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N94 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N93 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N92 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N91 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N90 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N89 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N88 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N87 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N86 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N85 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N84 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N83 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N82 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N81 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N80 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N79 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N78 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N77 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N76 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N75 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N74 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N73 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N72 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N71 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N70 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N69 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N68 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N67 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N66 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N65 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N64 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N63 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N62 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N61 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N60 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N59 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N58 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N57 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N56 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N55 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N54 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N53 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N52 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N51 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N50 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N49 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N48 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N47 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N46 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N45 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N44 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N43 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N42 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N41 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N40 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N39 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N38 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N37 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N36 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N35 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N34 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N33 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N32 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N31 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N30 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N29 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N28 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N27 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N26 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N25 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N24 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N23 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N22 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N21 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N20 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N19 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N18 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N17 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N16 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N15 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N14 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N13 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N12 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N11 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N10 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N9 ,
         \DLX_Datapath/ArithLogUnit/ALU_shift/N8 ,
         \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/S_1[1] ,
         \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/S_0[1] ,
         \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_0/S_0[1] ,
         \DLX_ControlUnit/N2798 , \DLX_ControlUnit/N2789 ,
         \DLX_ControlUnit/N2787 , \DLX_ControlUnit/N2785 , n54614, n54616,
         n54618, n54620, n54623, n57378, n57379, n57380, n57381, n57382,
         n57390, n57393, n57424, n57425, n57426, n57427, n57428, n57429,
         n57430, n57431, n58565, n58570, n58575, n58577, n58588, n58592,
         n58594, n58596, n58604, n58609, n58614, n58618, n58624, n58629,
         n58632, n58635, n58643, n58647, n58651, n58653, n58656, n58664,
         n58669, n58671, n58673, n58680, n58682, n58685, n58688, n58691,
         n58698, n58713, n58720, n58722, n58724, n58728, n58746, n58769,
         n58770, n58771, n58772, n58773, n58774, n58775, n58776, n58777,
         n58778, n58779, n58780, n58781, n58782, n58783, n58784, n58785,
         n58786, n58787, n58788, n58789, n58790, n58791, n58792, n58793,
         n58794, n58795, n58796, n58797, n58798, n58799, n58800, n58833,
         n58834, n58835, n58836, n58837, n58838, n58839, n58840, n58841,
         n58842, n58843, n58844, n58845, n58846, n58847, n58848, n58849,
         n58850, n58851, n58852, n58853, n58854, n58855, n58856, n58857,
         n58858, n58859, n58860, n58861, n58862, n58863, n58864, n58865,
         n58866, n58867, n58868, n58869, n58870, n58871, n58872, n58873,
         n58874, n58875, n58876, n58878, n58879, n58880, n58881, n58883,
         n58884, n58885, n58886, n58888, n58890, n58891, n58892, n58893,
         n58894, n58895, n58896, n58897, n58898, n58899, n58901, n58902,
         n58903, n58905, n58907, n58909, n58910, n58911, n58912, n58913,
         n58914, n58915, n58917, n58918, n58919, n58920, n58922, n58923,
         n58924, n58925, n58927, n58928, n58929, n58931, n58932, n58933,
         n58934, n58935, n58937, n58938, n58939, n58940, n58942, n58943,
         n58945, n58946, n58948, n58949, n58950, n58951, n58952, n58953,
         n58954, n58955, n58957, n58958, n58959, n58961, n58963, n58964,
         n58966, n58967, n58968, n58969, n58970, n58971, n58972, n58974,
         n58975, n58976, n58977, n58979, n58981, n58983, n58984, n58985,
         n58986, n58987, n58988, n58990, n58992, n58993, n58995, n58996,
         n58998, n58999, n59001, n59002, n59003, n59004, n59005, n59006,
         n59008, n59009, n59012, n59013, n59019, n59020, n59021, n59022,
         n59023, n59024, n59025, n59026, n59027, n59028, n59029, n59030,
         n59031, n59032, n59033, n59034, n59035, n59036, n59037, n59038,
         n59039, n59040, n59041, n59042, n59043, n59044, n59045, n59046,
         n59047, n59048, n59049, n59050, n59053, n59054, n59057, n59058,
         n59059, n59060, n59061, n59068, n59069, n59070, n59071, n59072,
         n59073, n59077, n59078, n59080, n59081, n59082, n59084, n59085,
         n59088, n59090, n59093, n59098, n59216, n59217, n59218, n59219,
         n59220, n59323, n59325, n59326, n59327, n59328, n59329, n59330,
         n59331, n59332, n59333, n59334, n59335, n59336, n59337, n59338,
         n59339, n59340, n59341, n59342, n59343, n59344, n59345, n59346,
         n59347, n59348, n59349, n59350, n59415, n59417, n59419, n59420,
         n59421, n59422, n59423, n59435, n59441, n59442, n59443, n59444,
         n59445, n59451, n59452, n59453, n59454, n59471, n59472, n59477,
         n59478, n59514, n59515, n59516, n59517, n59518, n60158, n60159,
         n60161, n60162, n60163, n60164, n60165, n60166, n60167, n60168,
         n60169, n60170, n60171, n60172, n60173, n60174, n60175, n60176,
         n60177, n60178, n60179, n60180, n60181, n60182, n60183, n60184,
         n60185, n60186, n60187, n60188, n60189, n60190, n60191, n60192,
         n60193, n60194, n60195, n60196, n60197, n60198, n60199, n60200,
         n60201, n60202, n60203, n60204, n60205, n60206, n60207, n60208,
         n60209, n60210, n60211, n60212, n60213, n60214, n60215, n60216,
         n60217, n60218, n60219, n60220, n60221, n60222, n60223, n60224,
         n60225, n60226, n60227, n60228, n60229, n60270, n60271, n60272,
         n60273, n60290, n60291, n60292, n60293, n60294, n60295, n60296,
         n60297, n60298, n60299, n60300, n60301, n60302, n60303, n60304,
         n60305, n60306, n60307, n60308, n60309, n60310, n60311, n60312,
         n60313, n60314, n60315, n60316, n60317, n60318, n60319, n60320,
         n60321, n60322, n60323, n60324, n60325, n60327, n60328, n60329,
         n60330, n60331, n60332, n60333, n60334, n60335, n60336, n60337,
         n60338, n60339, n60340, n60341, n60342, n60343, n60344, n60345,
         n60346, n60347, n60348, n60349, n60350, n60351, n60352, n60353,
         n60354, n60355, n60356, n60358, n60360, n60362, n60364, n60365,
         n60366, n60367, n60368, n60369, n60370, n60371, n60372, n60373,
         n60374, n60375, n60376, n60377, n60442, n60443,
         \dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[1] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[2] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[3] ,
         \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[2] ,
         \add_0_root_r2411/carry[7] , \add_0_root_r2411/carry[6] ,
         \add_0_root_sub_0_root_DLX_Datapath/RegisterFile/add_172/carry[6] ,
         \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ,
         net2410613, net2411291, net2411318, net2465147, net2465245,
         net2465244, net2465273, net2465400, n61539, n61540, n61666, n61670,
         n61799, n61904, n62027, n62182, n62183, n62185, n62189, n62190,
         n62191, n62194, n62196, n62197, n62198, n62199, n62200, n62201,
         n62202, n62204, n62212, n62245, n62247, n62496, n62573, n62574,
         n62661, n62662, n62664, n64126, n64127, n64246, n64247, n64266,
         n64267, n64652, n64655, n66263, n69283, n69289, n69292, n69303,
         n69307, n69313, n69315, n69319, n69321, n69322, n69323, n69324,
         n69325, n69326, n69330, n69339, n69340, n69343, n69346, n69347,
         n69348, n69349, n69350, n69351, n69352, n69353, n69354, n69355,
         n69356, n69357, n69358, n69359, n69362, n69369, n69377, n69378,
         n69379, n69380, n69381, n69382, n69413, n69414, n69415, n69416,
         n69417, n69424, n69425, n69426, n69429, n69430, n69459, n69460,
         n69463, n69464, n69465, n69466, n69469, n69470, n69483, n69484,
         n69486, n69490, n69492, n69498, n69503, n69507, n69509, n69511,
         n69514, n69515, n69519, n69521, n69524, n69526, n69529, n69538,
         n69541, n69543, n69545, n69549, n69553, n69555, n69560, n69561,
         n69564, n69567, n69571, n69577, n69578, n69581, n69583, n69588,
         n69589, n69591, n69595, n69597, n69603, n69612, n69614, n69616,
         n69620, n69624, n69626, n69629, n69631, n69634, n69643, n69646,
         n69648, n69654, n69658, n69660, n69665, n69666, n69682, n69683,
         n69688, n69689, n69694, n69697, n69698, n69699, n69700, n69701,
         n69702, n69703, n69704, n69705, n69706, n69707, n69708, n69709,
         n69710, n69711, n69712, n69713, n69714, n69715, n69716, n69717,
         n69718, n69719, n69720, n69721, n69722, n69723, n69724, n69725,
         n69726, n69727, n69728, n69729, n69730, n69765, n69784, n69785,
         n69786, n69787, n69788, n69789, n69790, n69791, n69792, n69793,
         n69794, n69795, n69796, n69797, n69798, n69799, n69800, n69801,
         n69802, n69975, n69991, n69994, n69998, n70000, n70006, n70015,
         n70017, n70019, n70023, n70027, n70029, n70032, n70034, n70037,
         n70046, n70049, n70051, n70057, n70061, n70063, n70068, n70069,
         n70085, n70086, n70091, n70097, n70098, n70105, n70107, n70108,
         n70110, n70125, n70127, n70130, n70142, n70147, n70151, n70153,
         n70159, n70168, n70170, n70172, n70176, n70180, n70182, n70185,
         n70187, n70190, n70199, n70202, n70204, n70206, n70208, n70209,
         n70210, n70214, n70216, n70221, n70222, n70225, n70228, n70238,
         n70239, n70242, n70244, n70249, n70250, n70251, n70258, n70260,
         n70261, n70263, n70278, n70280, n70283, n70291, n70295, n70297,
         n70303, n70304, n70308, n70312, n70314, n70316, n70317, n70320,
         n70321, n70324, n70326, n70329, n70330, n70331, n70334, n70342,
         n70343, n70346, n70348, n70350, n70354, n70355, n70358, n70360,
         n70363, n70364, n70365, n70366, n70367, n70369, n70372, n70376,
         n70382, n70383, n70386, n70388, n70394, n70395, n70402, n70404,
         n70405, n70407, n70422, n70424, n70427, n70433, n70437, n70439,
         n70445, n70446, n70450, n70454, n70456, n70458, n70461, n70462,
         n70463, n70466, n70468, n70470, n70471, n70472, n70473, n70474,
         n70476, n70484, n70485, n70488, n70490, n70492, n70494, n70496,
         n70497, n70500, n70502, n70506, n70507, n70508, n70511, n70514,
         n70518, n70524, n70525, n70530, n70535, n70536, n70537, n70544,
         n70546, n70547, n70549, n70564, n70566, n70569, n70575, n70576,
         n70577, n70580, n70584, n70586, n70592, n70601, n70603, n70605,
         n70609, n70613, n70615, n70618, n70619, n70620, n70623, n70631,
         n70632, n70635, n70637, n70639, n70643, n70647, n70649, n70652,
         n70654, n70655, n70656, n70658, n70664, n70671, n70672, n70675,
         n70677, n70683, n70684, n70691, n70693, n70694, n70696, n70711,
         n70713, n70717, n70726, n70729, n70733, n70735, n70741, n70750,
         n70752, n70754, n70758, n70762, n70764, n70767, n70769, n70772,
         n70781, n70784, n70786, n70792, n70796, n70798, n70803, n70804,
         n70820, n70821, n70826, n70832, n70833, n70840, n70842, n70843,
         n70845, n70860, n70862, n70872, n70880, n70882, n70884, n70888,
         n70892, n70894, n70900, n70909, n70911, n70913, n70917, n70921,
         n70923, n70926, n70928, n70931, n70940, n70943, n70945, n70951,
         n70955, n70957, n70962, n70963, n70979, n70980, n70985, n70991,
         n70992, n70999, n71001, n71002, n71004, n71019, n71021, n71026,
         n71033, n71037, n71039, n71045, n71054, n71056, n71058, n71062,
         n71066, n71068, n71071, n71073, n71076, n71085, n71088, n71090,
         n71096, n71100, n71102, n71107, n71108, n71124, n71125, n71130,
         n71136, n71137, n71144, n71146, n71147, n71149, n71164, n71166,
         n71169, n71179, n71182, n71186, n71188, n71194, n71203, n71205,
         n71207, n71211, n71215, n71217, n71220, n71222, n71225, n71234,
         n71237, n71239, n71245, n71249, n71251, n71256, n71257, n71262,
         n71266, n71273, n71274, n71279, n71285, n71286, n71293, n71295,
         n71296, n71298, n71313, n71315, n71325, n71327, n71329, n71331,
         n71335, n71337, n71343, n71352, n71354, n71356, n71360, n71364,
         n71366, n71369, n71371, n71374, n71383, n71386, n71388, n71394,
         n71398, n71400, n71405, n71406, n71422, n71423, n71428, n71429,
         n71434, n71435, n71442, n71444, n71445, n71447, n71462, n71464,
         n71469, n71482, n71486, n71488, n71494, n71503, n71505, n71507,
         n71511, n71515, n71517, n71520, n71522, n71525, n71534, n71537,
         n71539, n71545, n71549, n71551, n71556, n71557, n71573, n71574,
         n71579, n71585, n71586, n71593, n71595, n71596, n71598, n71613,
         n71615, n71618, n71626, n71630, n71632, n71638, n71647, n71649,
         n71651, n71655, n71659, n71661, n71664, n71666, n71669, n71678,
         n71681, n71683, n71689, n71693, n71695, n71700, n71701, n71717,
         n71718, n71723, n71729, n71730, n71737, n71739, n71740, n71742,
         n71757, n71759, n71762, n71772, n71775, n71779, n71781, n71787,
         n71796, n71798, n71800, n71804, n71808, n71810, n71813, n71815,
         n71818, n71827, n71830, n71832, n71838, n71842, n71844, n71849,
         n71850, n71866, n71867, n71872, n71878, n71879, n71886, n71888,
         n71889, n71891, n71906, n71908, n71913, n71922, n71924, n71926,
         n71929, n71933, n71935, n71941, n71950, n71952, n71954, n71958,
         n71962, n71964, n71967, n71969, n71972, n71981, n71984, n71986,
         n71992, n71996, n71997, n71998, n72003, n72004, n72020, n72021,
         n72026, n72032, n72033, n72040, n72042, n72043, n72045, n72060,
         n72062, n72065, n72073, n72077, n72079, n72085, n72094, n72096,
         n72098, n72102, n72106, n72108, n72111, n72113, n72116, n72125,
         n72128, n72130, n72136, n72140, n72142, n72147, n72148, n72164,
         n72165, n72170, n72171, n72176, n72177, n72184, n72186, n72187,
         n72189, n72204, n72206, n72209, n72224, n72228, n72230, n72236,
         n72245, n72247, n72249, n72253, n72257, n72259, n72262, n72264,
         n72267, n72276, n72279, n72281, n72287, n72291, n72293, n72298,
         n72299, n72315, n72316, n72321, n72327, n72328, n72335, n72337,
         n72338, n72340, n72355, n72357, n72362, n72370, n72372, n72375,
         n72379, n72381, n72387, n72396, n72398, n72400, n72404, n72408,
         n72410, n72413, n72415, n72418, n72427, n72430, n72432, n72438,
         n72442, n72444, n72449, n72450, n72466, n72467, n72472, n72478,
         n72479, n72486, n72488, n72489, n72491, n72506, n72508, n72511,
         n72523, n72527, n72529, n72535, n72544, n72546, n72548, n72552,
         n72556, n72558, n72561, n72563, n72566, n72575, n72578, n72580,
         n72586, n72590, n72592, n72597, n72598, n72600, n72603, n72607,
         n72614, n72615, n72620, n72626, n72627, n72634, n72636, n72637,
         n72639, n72654, n72656, n72661, n72665, n72669, n72671, n72677,
         n72686, n72688, n72690, n72694, n72698, n72700, n72703, n72705,
         n72708, n72717, n72720, n72722, n72728, n72732, n72734, n72739,
         n72740, n72745, n72756, n72757, n72762, n72768, n72769, n72776,
         n72778, n72779, n72781, n72796, n72798, n72803, n72808, n72830,
         n72833, n72837, n72839, n72845, n72854, n72856, n72858, n72862,
         n72866, n72868, n72871, n72873, n72876, n72885, n72888, n72890,
         n72896, n72900, n72902, n72907, n72908, n72924, n72925, n72930,
         n72936, n72937, n72944, n72946, n72947, n72949, n72964, n72966,
         n72969, n72978, n72980, n72983, n72987, n72989, n72995, n73004,
         n73006, n73008, n73012, n73016, n73017, n73018, n73021, n73023,
         n73026, n73035, n73038, n73040, n73046, n73050, n73052, n73057,
         n73058, n73074, n73075, n73080, n73086, n73087, n73094, n73096,
         n73097, n73099, n73114, n73116, n73120, n73125, n73129, n73131,
         n73137, n73146, n73148, n73150, n73154, n73158, n73159, n73160,
         n73163, n73165, n73168, n73177, n73180, n73182, n73188, n73192,
         n73194, n73199, n73200, n73216, n73217, n73222, n73228, n73229,
         n73236, n73238, n73239, n73241, n73256, n73258, n73263, n73267,
         n73271, n73273, n73279, n73288, n73290, n73292, n73296, n73300,
         n73301, n73302, n73305, n73307, n73310, n73319, n73322, n73324,
         n73330, n73334, n73336, n73341, n73342, n73358, n73359, n73364,
         n73370, n73371, n73378, n73380, n73381, n73383, n73398, n73400,
         n73405, n73411, n73414, n73418, n73420, n73426, n73435, n73437,
         n73439, n73442, n73443, n73447, n73448, n73449, n73452, n73454,
         n73457, n73461, n73466, n73469, n73471, n73476, n73477, n73481,
         n73483, n73484, n73488, n73489, n73505, n73506, n73511, n73517,
         n73518, n73525, n73527, n73528, n73530, n73545, n73547, n73552,
         n73558, n73560, n73563, n73567, n73569, n73575, n73584, n73586,
         n73588, n73591, n73592, n73596, n73597, n73598, n73601, n73603,
         n73606, n73615, n73618, n73620, n73625, n73626, n73627, n73630,
         n73632, n73637, n73638, n73654, n73655, n73660, n73666, n73667,
         n73674, n73676, n73677, n73679, n73694, n73696, n73699, n73710,
         n73714, n73716, n73722, n73731, n73733, n73735, n73738, n73739,
         n73743, n73744, n73745, n73748, n73750, n73753, n73757, n73762,
         n73765, n73767, n73772, n73773, n73777, n73779, n73780, n73784,
         n73785, n73801, n73802, n73805, n73807, n73812, n73813, n73814,
         n73821, n73823, n73824, n73826, n73841, n73843, n73847, n73851,
         n73855, n73857, n73863, n73872, n73874, n73876, n73879, n73880,
         n73884, n73885, n73886, n73889, n73891, n73894, n73903, n73906,
         n73908, n73913, n73914, n73918, n73920, n73925, n73926, n73942,
         n73943, n73953, n73954, n73955, n73962, n73964, n73965, n73967,
         n73982, n73984, n73988, n73993, n73997, n73999, n74005, n74014,
         n74016, n74018, n74021, n74022, n74026, n74028, n74031, n74032,
         n74033, n74036, n74044, n74045, n74048, n74050, n74052, n74055,
         n74056, n74057, n74060, n74061, n74062, n74065, n74067, n74068,
         n74069, n74071, n74077, n74084, n74085, n74088, n74090, n74095,
         n74096, n74097, n74104, n74106, n74107, n74109, n74124, n74126,
         n74130, n74134, n74138, n74140, n74146, n74155, n74157, n74159,
         n74162, n74163, n74167, n74169, n74172, n74174, n74177, n74186,
         n74189, n74191, n74196, n74197, n74201, n74203, n74206, n74208,
         n74209, n74210, n74212, n74218, n74225, n74226, n74229, n74231,
         n74237, n74238, n74245, n74247, n74248, n74250, n74265, n74267,
         n74270, n74274, n74278, n74280, n74286, n74295, n74297, n74299,
         n74302, n74303, n74307, n74309, n74312, n74314, n74317, n74319,
         n74326, n74329, n74331, n74336, n74337, n74338, n74341, n74342,
         n74343, n74348, n74349, n74365, n74366, n74371, n74377, n74378,
         n74385, n74387, n74388, n74390, n74405, n74407, n74410, n79652,
         n79653, n79654, n79655, n79656, n79657, n79658, n79659, n79660,
         n79661, n79662, n79663, n79664, n79665, n79666, n79667, n79668,
         n79669, n79670, n79671, n79672, n79673, n79674, n79675, n79676,
         n79677, n79678, n79679, n79680, n79681, n79682, n79683, n79684,
         n79685, n79686, n79687, n79688, n79689, n79690, n79691, n79692,
         n79693, n79694, n79695, n79696, n79697, n79698, n79699, n79700,
         n79701, n79702, n79703, n79704, n79705, n79706, n79707, n79708,
         n79709, n79710, n79711, n79712, n79713, n79714, n79715, n79716,
         n79717, n79718, n79719, n79720, n79721, n79722, n79723, n79724,
         n79725, n79726, n79727, n79728, n79729, n79730, n79731, n79732,
         n79733, n79734, n79735, n79736, n79737, n79738, n79739, n79740,
         n79741, n79743, n79744, n79745, n79746, n79747, n79748, n79749,
         n79750, n79751, n79752, n79753, n79754, n79755, n79756, n79757,
         n79758, n79759, n79760, n79761, n79762, n79763, n79764, n79765,
         n79766, n79767, n79768, n79769, n79770, n79771, n79772, n79773,
         n79774, n79775, n79776, n79778, n79779, n79780, n79781, n79782,
         n79783, n79784, n79785, n79786, n79787, n79788, n79789, n79790,
         n79791, n79792, n79793, n79794, n79795, n79796, n79797, n79798,
         n79799, n79800, n79801, n79802, n79803, n79804, n79805, n79806,
         n79807, n79808, n79809, n79811, n79812, n79813, n79814, n79815,
         n79816, n79817, n79818, n79819, n79820, n79821, n79822, n79823,
         n79824, n79825, n79826, n79827, n79828, n79829, n79830, n79831,
         n79832, n79833, n79834, n79835, n79836, n79837, n79838, n79839,
         n79840, n79841, n79842, n79844, n79845, n79846, n79847, n79848,
         n79849, n79850, n79851, n79852, n79853, n79854, n79855, n79856,
         n79857, n79858, n79859, n79860, n79861, n79862, n79863, n79864,
         n79865, n79866, n79867, n79868, n79869, n79870, n79871, n79872,
         n79873, n79874, n79875, n79877, n79878, n79879, n79880, n79881,
         n79882, n79883, n79884, n79885, n79886, n79887, n79888, n79889,
         n79890, n79891, n79892, n79893, n79894, n79895, n79896, n79897,
         n79898, n79899, n79900, n79901, n79902, n79903, n79904, n79905,
         n79906, n79907, n79908, n79910, n79911, n79912, n79913, n79914,
         n79915, n79916, n79917, n79918, n79919, n79920, n79921, n79922,
         n79923, n79924, n79925, n79926, n79927, n79928, n79929, n79930,
         n79931, n79932, n79933, n79934, n79935, n79936, n79937, n79938,
         n79939, n79940, n79941, n79943, n79944, n79945, n79946, n79947,
         n79948, n79949, n79950, n79951, n79952, n79953, n79954, n79955,
         n79956, n79957, n79958, n79959, n79960, n79961, n79962, n79963,
         n79964, n79965, n79966, n79967, n79968, n79969, n79970, n79971,
         n79972, n79973, n79974, n79975, n79976, n79977, n79978, n79979,
         n79980, n79981, n79982, n79983, n79984, n79985, n79986, n79987,
         n79988, n79989, n79990, n79991, n79992, n79993, n79994, n79995,
         n79996, n79997, n79998, n79999, n80000, n80001, n80002, n80003,
         n80004, n80005, n80006, n80007, n80008, n80009, n80010, n80011,
         n80012, n80013, n80014, n80015, n80016, n80017, n80018, n80019,
         n80020, n80021, n80022, n80023, n80024, n80025, n80026, n80027,
         n80028, n80029, n80030, n80031, n80032, n80033, n80034, n80035,
         n80036, n80037, n80038, n80039, n80040, n80041, n80042, n80043,
         n80044, n80045, n80046, n80047, n80048, n80049, n80050, n80051,
         n80052, n80053, n80054, n80055, n80056, n80057, n80058, n80059,
         n80060, n80061, n80062, n80063, n80064, n80065, n80066, n80067,
         n80068, n80069, n80070, n80071, n80072, n80073, n80074, n80075,
         n80076, n80077, n80078, n80079, n80080, n80081, n80082, n80083,
         n80084, n80085, n80086, n80087, n80088, n80089, n80090, n80091,
         n80092, n80093, n80094, n80095, n80096, n80097, n80098, n80099,
         n80100, n80101, n80103, n80104, n80105, n80106, n80107, n80108,
         n80109, n80110, n80111, n80112, n80113, n80114, n80115, n80116,
         n80117, n80118, n80119, n80120, n80121, n80122, n80123, n80124,
         n80125, n80126, n80127, n80128, n80129, n80130, n80131, n80132,
         n80133, n80134, n80135, n80136, n80137, n80138, n80139, n80140,
         n80141, n80142, n80143, n80144, n80145, n80146, n80147, n80148,
         n80149, n80150, n80151, n80152, n80153, n80154, n80155, n80156,
         n80157, n80158, n80159, n80160, n80161, n80162, n80163, n80164,
         n80165, n80166, n80167, n80168, n80169, n80170, n80171, n80172,
         n80173, n80174, n80175, n80176, n80177, n80178, n80179, n80180,
         n80181, n80182, n80183, n80184, n80185, n80186, n80188, n80189,
         n80190, n80191, n80192, n80193, n80194, n80195, n80196, n80197,
         n80198, n80199, n80200, n80201, n80202, n80203, n80204, n80205,
         n80206, n80207, n80208, n80209, n80210, n80211, n80212, n80213,
         n80214, n80215, n80216, n80217, n80218, n80219, n80220, n80221,
         n80222, n80223, n80224, n80225, n80226, n80227, n80228, n80229,
         n80230, n80231, n80232, n80233, n80234, n80235, n80236, n80237,
         n80238, n80239, n80240, n80241, n80242, n80243, n80244, n80245,
         n80246, n80247, n80248, n80249, n80250, n80251, n80252, n80253,
         n80254, n80255, n80256, n80257, n80258, n80259, n80260, n80261,
         n80262, n80263, n80264, n80265, n80266, n80267, n80268, n80269,
         n80270, n80271, n80272, n80273, n80274, n80275, n80276, n80277,
         n80278, n80279, n80280, n80281, n80282, n80283, n80284, n80285,
         n80286, n80287, n80288, n80289, n80290, n80291, n80292, n80293,
         n80294, n80295, n80296, n80297, n80298, n80299, n80300, n80301,
         n80302, n80303, n80304, n80305, n80306, n80307, n80308, n80309,
         n80310, n80311, n80312, n80313, n80314, n80315, n80316, n80317,
         n80318, n80319, n80320, n80321, n80322, n80323, n80324, n80325,
         n80326, n80327, n80328, n80329, n80330, n80331, n80332, n80333,
         n80334, n80335, n80336, n80337, n80338, n80339, n80340, n80341,
         n80342, n80343, n80344, n80345, n80346, n80347, n80348, n80349,
         n80350, n80351, n80352, n80353, n80354, n80355, n80356, n80357,
         n80358, n80359, n80360, n80361, n80362, n80363, n80364, n80365,
         n80366, n80367, n80368, n80369, n80370, n80371, n80372, n80373,
         n80374, n80375, n80376, n80377, n80378, n80379, n80380, n80381,
         n80382, n80383, n80384, n80385, n80386, n80387, n80388, n80389,
         n80390, n80391, n80392, n80393, n80394, n80395, n80396, n80397,
         n80398, n80399, n80400, n80401, n80402, n80403, n80404, n80405,
         n80406, n80407, n80408, n80409, n80410, n80411, n80412, n80413,
         n80414, n80415, n80416, n80417, n80418, n80419, n80420, n80421,
         n80422, n80423, n80424, n80425, n80426, n80427, n80428, n80429,
         n80430, n80431, n80432, n80433, n80434, n80435, n80436, n80437,
         n80438, n80439, n80440, n80441, n80442, n80443, n80444, n80445,
         n80446, n80447, n80448, n80449, n80450, n80451, n80452, n80453,
         n80454, n80455, n80456, n80457, n80458, n80459, n80460, n80461,
         n80462, n80463, n80464, n80465, n80466, n80467, n80468, n80469,
         n80470, n80471, n80472, n80473, n80474, n80475, n80476, n80477,
         n80478, n80479, n80480, n80481, n80482, n80483, n80484, n80485,
         n80486, n80487, n80488, n80489, n80490, n80491, n80492, n80493,
         n80494, n80495, n80496, n80497, n80498, n80499, n80500, n80501,
         n80502, n80503, n80504, n80505, n80506, n80507, n80508, n80509,
         n80510, n80511, n80512, n80513, n80514, n80515, n80516, n80517,
         n80518, n80519, n80520, n80521, n80522, n80523, n80524, n80525,
         n80526, n80527, n80528, n80529, n80530, n80531, n80532, n80533,
         n80534, n80535, n80536, n80537, n80538, n80539, n80540, n80541,
         n80542, n80543, n80544, n80545, n80546, n80547, n80548, n80549,
         n80550, n80551, n80552, n80553, n80554, n80555, n80556, n80557,
         n80558, n80559, n80560, n80561, n80562, n80563, n80564, n80565,
         n80566, n80567, n80568, n80569, n80570, n80571, n80572, n80573,
         n80574, n80575, n80576, n80577, n80578, n80579, n80580, n80581,
         n80582, n80583, n80584, n80585, n80586, n80587, n80588, n80589,
         n80590, n80591, n80592, n80593, n80594, n80595, n80596, n80597,
         n80598, n80599, n80600, n80601, n80602, n80603, n80604, n80605,
         n80606, n80607, n80608, n80609, n80610, n80611, n80612, n80613,
         n80614, n80615, n80616, n80617, n80618, n80619, n80620, n80621,
         n80622, n80623, n80624, n80625, n80626, n80627, n80628, n80629,
         n80630, n80631, n80632, n80633, n80634, n80635, n80636, n80637,
         n80638, n80639, n80640, n80641, n80642, n80643, n80644, n80645,
         n80646, n80647, n80648, n80649, n80650, n80651, n80652, n80653,
         n80654, n80655, n80656, n80657, n80658, n80659, n80660, n80661,
         n80662, n80663, n80664, n80665, n80666, n80667, n80668, n80669,
         n80670, n80671, n80672, n80673, n80674, n80675, n80676, n80677,
         n80678, n80679, n80680, n80681, n80682, n80683, n80684, n80685,
         n80686, n80687, n80688, n80689, n80690, n80691, n80692, n80693,
         n80694, n80695, n80696, n80697, n80698, n80699, n80700, n80701,
         n80702, n80703, n80704, n80705, n80706, n80707, n80708, n80709,
         n80710, n80711, n80712, n80713, n80714, n80715, n80716, n80717,
         n80718, n80719, n80720, n80721, n80722, n80723, n80724, n80725,
         n80726, n80727, n80728, n80729, n80730, n80731, n80732, n80733,
         n80734, n80735, n80736, n80737, n80738, n80739, n80740, n80741,
         n80742, n80743, n80744, n80745, n80746, n80747, n80748, n80749,
         n80750, n80751, n80752, n80753, n80754, n80755, n80756, n80757,
         n80758, n80759, n80760, n80761, n80762, n80763, n80764, n80765,
         n80766, n80767, n80768, n80769, n80770, n80771, n80772, n80773,
         n80774, n80775, n80776, n80777, n80778, n80779, n80780, n80781,
         n80782, n80783, n80784, n80785, n80786, n80787, n80788, n80789,
         n80790, n80791, n80792, n80793, n80794, n80795, n80796, n80797,
         n80798, n80799, n80800, n80801, n80802, n80803, n80804, n80805,
         n80806, n80807, n80808, n80809, n80810, n80811, n80812, n80813,
         n80814, n80815, n80816, n80817, n80818, n80819, n80820, n80821,
         n80822, n80823, n80824, n80825, n80826, n80827, n80828, n80829,
         n80830, n80831, n80832, n80833, n80834, n80835, n80836, n80837,
         n80838, n80839, n80840, n80841, n80842, n80843, n80844, n80845,
         n80846, n80847, n80848, n80849, n80850, n80851, n80852, n80853,
         n80854, n80855, n80856, n80857, n80858, n80859, n80860, n80861,
         n80862, n80863, n80864, n80865, n80866, n80867, n80868, n80869,
         n80870, n80871, n80872, n80873, n80874, n80875, n80876, n80877,
         n80878, n80879, n80880, n80881, n80882, n80883, n80884, n80885,
         n80886, n80887, n80888, n80889, n80890, n80891, n80892, n80893,
         n80894, n80895, n80896, n80897, n80898, n80899, n80900, n80901,
         n80902, n80903, n80904, n80905, n80906, n80907, n80908, n80909,
         n80910, n80911, n80912, n80913, n80914, n80915, n80916, n80917,
         n80918, n80919, n80920, n80921, n80922, n80923, n80924, n80925,
         n80926, n80927, n80928, n80929, n80930, n80931, n80932, n80933,
         n80934, n80935, n80936, n80937, n80938, n80939, n80940, n80941,
         n80942, n80943, n80944, n80945, n80946, n80947, n80948, n80949,
         n80950, n80951, n80952, n80953, n80954, n80955, n80956, n80957,
         n80958, n80959, n80960, n80961, n80962, n80963, n80964, n80965,
         n80966, n80967, n80968, n80969, n80970, n80971, n80972, n80973,
         n80974, n80975, n80976, n80977, n80978, n80979, n80980, n80981,
         n80982, n80983, n80984, n80985, n80986, n80987, n80988, n80989,
         n80990, n80991, n80992, n80993, n80994, n80995, n80996, n80997,
         n80998, n80999, n81000, n81001, n81002, n81003, n81004, n81005,
         n81006, n81007, n81008, n81009, n81010, n81011, n81012, n81013,
         n81014, n81015, n81016, n81017, n81018, n81019, n81020, n81021,
         n81022, n81023, n81024, n81025, n81026, n81027, n81028, n81029,
         n81030, n81031, n81032, n81033, n81034, n81035, n81036, n81037,
         n81038, n81039, n81040, n81041, n81042, n81043, n81044, n81045,
         n81046, n81047, n81048, n81049, n81050, n81051, n81052, n81053,
         n81054, n81055, n81056, n81057, n81058, n81059, n81060, n81061,
         n81062, n81063, n81064, n81065, n81066, n81067, n81068, n81069,
         n81070, n81071, n81072, n81073, n81074, n81075, n81076, n81077,
         n81078, n81079, n81080, n81081, n81082, n81083, n81084, n81085,
         n81086, n81087, n81088, n81089, n81090, n81091, n81092, n81093,
         n81094, n81095, n81096, n81097, n81098, n81099, n81100, n81101,
         n81102, n81103, n81104, n81105, n81106, n81107, n81108, n81109,
         n81110, n81111, n81112, n81113, n81114, n81115, n81116, n81117,
         n81118, n81119, n81120, n81121, n81122, n81123, n81124, n81125,
         n81126, n81127, n81128, n81129, n81130, n81131, n81132, n81133,
         n81134, n81135, n81136, n81137, n81138, n81139, n81140, n81141,
         n81142, n81143, n81144, n81145, n81146, n81147, n81148, n81149,
         n81150, n81151, n81152, n81153, n81154, n81155, n81156, n81157,
         n81158, n81159, n81160, n81161, n81162, n81163, n81164, n81165,
         n81166, n81167, n81168, n81169, n81170, n81171, n81172, n81173,
         n81174, n81175, n81176, n81177, n81178, n81179, n81180, n81181,
         n81182, n81183, n81184, n81185, n81186, n81187, n81188, n81189,
         n81190, n81191, n81192, n81193, n81194, n81195, n81196, n81197,
         n81198, n81199, n81200, n81201, n81202, n81203, n81204, n81205,
         n81206, n81207, n81208, n81209, n81210, n81211, n81212, n81213,
         n81214, n81215, n81216, n81217, n81218, n81219, n81220, n81221,
         n81222, n81223, n81224, n81225, n81226, n81227, n81228, n81229,
         n81230, n81231, n81232, n81233, n81234, n81235, n81236, n81238,
         n81239, n81240, n81241, n81242, n81243, n81244, n81247, n81248,
         n81249, n81250, n81251, n81252, n81253, n81254, n81255, n81256,
         n81257, n81258, n81259, n81260, n81261, n81262, n81263, n81264,
         n81265, n81266, n81267, n81268, n81269, n81270, n81271, n81272,
         n81273, n81274, n81275, n81276, n81277, n81278, n81279, n81280,
         n81281, n81282, n81283, n81284, n81285, n81286, n81287, n81289,
         n81290, n81291, n81292, n81293, n81294, n81295, n81296, n81297,
         n81299, n81300, n81301, n81302, n81303, n81304, n81305, n81306,
         n81307, n81308, n81309, n81310, n81311, n81312, n81313, n81314,
         n81315, n81316, n81317, n81318, n81319, n81320, n81321, n81322,
         n81323, n81324, n81325, n81326, n81327, n81328, n81329, n81330,
         n81331, n81332, n81333, n81334, n81335, n81336, n81337, n81338,
         n81339, n81340, n81341, n81342, n81343, n81344, n81345, n81346,
         n81347, n81348, n81349, n81350, n81351, n81352, n81353, n81354,
         n81355, n81356, n81357, n81358, n81359, n81360, n81361, n81362,
         n81363, n81364, n81365, n81366, n81367, n81368, n81369, n81370,
         n81371, n81372, n81373, n81374, n81375, n81376, n81377, n81378,
         n81379, n81380, n81381, n81382, n81383, n81384, n81385, n81386,
         n81387, n81388, n81389, n81390, n81391, n81392, n81393, n81394,
         n81395, n81396, n81397, n81398, n81399, n81400, n81401, n81402,
         n81403, n81404, n81405, n81406, n81407, n81408, n81409, n81410,
         n81411, n81412, n81413, n81414, n81415, n81416, n81417, n81418,
         n81419, n81420, n81421, n81422, n81423, n81424, n81425, n81426,
         n81427, n81428, n81429, n81430, n81431, n81432, n81433, n81434,
         n81435, n81436, n81437, n81438, n81439, n81440, n81441, n81442,
         n81443, n81444, n81445, n81446, n81447, n81448, n81449, n81450,
         n81451, n81452, n81453, n81454, n81455, n81456, n81457, n81458,
         n81459, n81460, n81461, n81462, n81463, n81464, n81465, n81466,
         n81467, n81468, n81469, n81470, n81471, n81472, n81473, n81474,
         n81475, n81476, n81477, n81478, n81479, n81480, n81481, n81482,
         n81483, n81484, n81485, n81486, n81487, n81488, n81489, n81490,
         n81491, n81492, n81493, n81494, n81495, n81496, n81497, n81498,
         n81499, n81500, n81501, n81502, n81503, n81504, n81505, n81506,
         n81507, n81508, n81509, n81510, n81511, n81512, n81513, n81514,
         n81515, n81516, n81517, n81518, n81519, n81520, n81521, n81522,
         n81523, n81524, n81525, n81526, n81527, n81528, n81529, n81530,
         n81531, n81532, n81533, n81534, n81535, n81536, n81537, n81538,
         n81539, n81540, n81541, n81543, n81544, n81545, n81546, n81547,
         n81548, n81549, n81550, n81551, n81552, n81553, n81554, n81555,
         n81556, n81557, n81558, n81559, n81560, n81561, n81562, n81563,
         n81564, n81565, n81566, n81567, n81568, n81569, n81570, n81571,
         n81572, n81573, n81574, n81575, n81576, n81577, n81578, n81579,
         n81580, n81581, n81582, n81583, n81584, n81585, n81586, n81587,
         n81588, n81589, n81590, n81591, n81592, n81593, n81594, n81595,
         n81596, n81597, n81598, n81599, n81600, n81601, n81602, n81603,
         n81604, n81605, n81606, n81607, n81608, n81609, n81610, n81611,
         n81612, n81613, n81614, n81615, n81616, n81617, n81618, n81619,
         n81620, n81623, n81624, n81625, n81626, n81627, n81628, n81629,
         n81630, n81632, n81634, n81635, n81638, n81639, n81640, n81641,
         n81642, n81643, n81644, n81645, n81646, n81647, n81648, n81649,
         n81651, n81652, n81653, n81654, n81655, n81656, n81657, n81658,
         n81659, n81660, n81661, n81662, n81663, n81664, n81665, n81666,
         n81667, n81668, n81669, n81670, n81671, n81672, n81673, n81674,
         n81675, n81676, n81677, n81678, n81679, n81680, n81681, n81682,
         n81683, n81684, n81685, n81686, n81687, n81688, n81689, n81690,
         n81691, n81692, n81693, n81694, n81695, n81696, n81697, n81698,
         n81699, n81700, n81701, n81702, n81703, n81704, n81705, n81706,
         n81707, n81708, n81709, n81710, n81711, n81712, n81713, n81714,
         n81715, n81716, n81717, n81718, n81719, n81720, n81721, n81722,
         n81723, n81724, n81725, n81726, n81727, n81728, n81729, n81730,
         n81731, n81732, n81733, n81734, n81735, n81737, n81738, n81739,
         n81740, n81741, n81742, n81743, n81744, n81745, n81746, n81749,
         n81750, n81751, n81752, n81753, n81754, n81755, n81756, n81757,
         n81758, n81759, n81760, n81761, n81762, n81763, n81764, n81765,
         n81766, n81767, n81768, n81769, n81770, n81771, n81772, n81773,
         n81774, n81775, n81776, n81777, n81778, n81779, n81780, n81781,
         n81782, n81783, n81784, n81785, n81786, n81788, n81789, n81790,
         n81791, n81792, n81793, n81794, n81795, n81796, n81797, n81798,
         n81799, n81800, n81801, n81802, n81803, n81804, n81805, n81806,
         n81807, n81808, n81809, n81810, n81811, n81812, n81813, n81814,
         n81815, n81816, n81817, n81818, n81819, n81820, n81821, n81822,
         n81823, n81824, n81825, n81826, n81827, n81828, n81829, n81830,
         n81831, n81832, n81833, n81834, n81835, n81836, n81837, n81838,
         n81839, n81840, n81841, n81842, n81843, n81844, n81845, n81846,
         n81847, n81848, n81849, n81850, n81851, n81852, n81853, n81854,
         n81855, n81856, n81857, n81858, n81859, n81860, n81861, n81862,
         n81863, n81864, n81865, n81866, n81867, n81868, n81869, n81870,
         n81871, n81872, n81873, n81874, n81875, n81876, n81877, n81878,
         n81879, n81880, n81881, n81882, n81883, n81884, n81885, n81886,
         n81887, n81888, n81889, n81890, n81891, n81892, n81893, n81894,
         n81895, n81896, n81897, n81898, n81899, n81900, n81901, n81902,
         n81903, n81904, n81905, n81906, n81907, n81908, n81909, n81910,
         n81911, n81912, n81913, n81914, n81915, n81916, n81917, n81918,
         n81919, n81920, n81921, n81922, n81923, n81924, n81925, n81926,
         n81927, n81928, n81929, n81930, n81931, n81932, n81933, n81934,
         n81935, n81936, n81937, n81938, n81939, n81940, n81941, n81942,
         n81943, n81944, n81945, n81946, n81947, n81948, n81949, n81950,
         n81951, n81952, n81953, n81954, n81955, n81956, n81957, n81958,
         n81959, n81960, n81961, n81962, n81963, n81964, n81965, n81966,
         n81967, n81968, n81969, n81970, n81971, n81972, n81973, n81974,
         n81975, n81976, n81977, n81978, n81979, n81980, n81981, n81982,
         n81983, n81984, n81985, n81986, n81987, n81988, n81989, n81990,
         n81991, n81992, n81993, n81994, n81995, n81996, n81998, n82000,
         n82001, n82002, n82003, n82004, n82005, n82006, n82007, n82008,
         n82009, n82010, n82011, n82012, n82014, n82015, n82016, n82017,
         n82018, n82019, n82020, n82021, n82022, n82023, n82024, n82025,
         n82026, n82027, n82028, n82029, n82030, n82031, n82033, n82034,
         n82035, n82036, n82037, n82038, n82039, n82040, n82041, n82042,
         n82043, n82044, n82045, n82046, n82047, n82048, n82049, n82050,
         n82051, n82052, n82053, n82054, n82055, n82056, n82057, n82058,
         n82059, n82060, n82061, n82062, n82063, n82064, n82065, n82066,
         n82067, n82068, n82070, n82071, n82072, n82073, n82074, n82075,
         n82076, n82077, n82078, n82079, n82080, n82081, n82082, n82083,
         n82084, n82085, n82086, n82087, n82088, n82089, n82090, n82092,
         n82093, n82094, n82095, n82096, n82097, n82099, n82100, n82101,
         n82102, n82103, n82104, n82105, n82106, n82107, n82108, n82109,
         n82111, n82112, n82113, n82114, n82115, n82116, n82117, n82118,
         n82119, n82120, n82121, n82122, n82123, n82124, n82125, n82126,
         n82127, n82128, n82129, n82130, n82131, n82132, n82133, n82134,
         n82135, n82136, n82137, n82138, n82139, n82140, n82141, n82142,
         n82143, n82144, n82145, n82146, n82147, n82148, n82149, n82150,
         n82151, n82152, n82153, n82154, n82155, n82156, n82157, n82158,
         n82159, n82160, n82161, n82162, n82163, n82164, n82165, n82166,
         n82167, n82168, n82169, n82170, n82171, n82172, n82173, n82174,
         n82175, n82176, n82177, n82178, n82179, n82180, n82183, n82184,
         n82185, n82186, n82187, n82188, n82189, n82190, n82191, n82192,
         n82193, n82194, n82195, n82196, n82197, n82198, n82199, n82200,
         n82202, n82203, n82204, n82205, n82206, n82207, n82208, n82211,
         n82212, n82213, n82214, n82215, n82216, n82217, n82218, n82219,
         n82220, n82223, n82224, n82225, n82226, n82227, n82228, n82229,
         n82230, n82231, n82232, n82233, n82234, n82235, n82236, n82237,
         n82238, n82239, n82240, n82241, n82243, n82244, n82245, n82246,
         n82248, n82249, n82250, n82251, n82252, n82253, n82254, n82255,
         n82256, n82258, n82259, n82260, n82261, n82263, n82264, n82265,
         n82266, n82267, n82268, n82269, n82271, n82272, n82274, n82275,
         n82276, n82277, n82278, n82280, n82281, n82282, n82283, n82284,
         n82286, n82287, n82289, n82290, n82291, n82292, n82293, n82294,
         n82295, n82296, n82297, n82298, n82299, n82300, n82301, n82302,
         n82303, n82304, n82306, n82308, n82309, n82311, n82312, n82313,
         n82314, n82315, n82316, n82317, n82318, n82319, n82320, n82321,
         n82322, n82323, n82324, n82325, n82326, n82327, n82328, n82329,
         n82330, n82331, n82332, n82333, n82334, n82335, n82336, n82337,
         n82338, n82339, n82340, n82341, n82342, n82343, n82344, n82345,
         n82346, n82347, n82348, n82349, n82350, n82351, n82352, n82353,
         n82354, n82355, n82356, n82357, n82358, n82359, n82360, n82361,
         n82362, n82363, n82364, n82365, n82366, n82367, n82368, n82369,
         n82371, n82372, n82373, n82374, n82375, n82376, n82377, n82378,
         n82380, n82381, n82382, n82384, n82385, n82386, n82387, n82388,
         n82389, n82390, n82391, n82392, n82393, n82394, n82395, n82396,
         n82397, n82398, n82399, n82400, n82401, n82402, n82403, n82404,
         n82405, n82406, n82407, n82408, n82409, n82410, n82411, n82412,
         n82413, n82420, n82426, n82427, n82428, n82429, n82430, n82431,
         n82432, n82433, n82434, n82435, n82436, n82437, n82438, n82439,
         n82440, n82441, n82442, n82443, n82444, n82445, n82446, n82447,
         n82448, n82449, n82450, n82451, n82452, n82453, n82454, n82455,
         n82456, n82457, n82458, n82459, n82461, n82463, n82464, n82465,
         n82466, n82468, n82469, n82471, n82473, n82474, n82475, n82476,
         n82478, n82479, n82480, n82481, n82482, n82483, n82484, n82485,
         n82486, n82487, n82488, n82490, n82491, n82493, n82494, n82495,
         n82496, n82497, n82498, n82500, n82502, n82503, n82504, n82505,
         n82506, n82507, n82508, n82509, n82510, n82511, n82512, n82513,
         n82514, n82515, n82516, n82517, n82518, n82519, n82520, n82521,
         n82522, n82523, n82524, n82525, n82526, n82527, n82528, n82529,
         n82530, n82531, n82532, n82533, n82534, n82536, n82537, n82538,
         n82539, n82540, n82541, n82542, n82543, n82544, n82545, n82546,
         n82547, n82548, n82549, n82550, n82551, n82552, n82553, n82554,
         n82555, n82556, n82557, n82558, n82559, n82560, n82561, n82562,
         n82563, n82564, n82565, n82566, n82567, n82568, n82569, n82570,
         n82571, n82572, n82573, n82574, n82575, n82576, n82577, n82578,
         n82579, n82580, n82581, n82582, n82583, n82584, n82585, n82586,
         n82587, n82588, n82589, n82590, n82591, n82592, n82593, n82594,
         n82595, n82596, n82597, n82598, n82599, n82600, n82601, n82602,
         n82603, n82604, n82605, n82606, n82607, n82608, n82609, n82610,
         n82611, n82612, n82613, n82614, n82615, n82616, n82617, n82618,
         n82619, n82620, n82621, n82622, n82623, n82624, n82625, n82626,
         n82627, n82628, n82629, n82630, n82631, n82632, n82633, n82634,
         n82635, n82636, n82637, n82638, n82639, n82640, n82641, n82642,
         n82643, n82645, n82646, n82647, n82648, n82649, n82650, n82651,
         n82652, n82653, n82654, n82655, n82656, n82657, n82659, n82660,
         n82661, n82662, n82663, n82664, n82665, n82666, n82667, n82668,
         n82669, n82670, n82671, n82672, n82673, n82674, n82675, n82676,
         n82677, n82678, n82679, n82680, n82681, n82682, n82686, n82687,
         n82688, n82689, n82690, n82691, n82692, n82693, n82694, n82695,
         n82696, n82697, n82698, n82699, n82700, n82701, n82702, n82703,
         n82704, n82705, n82706, n82707, n82708, n82709, n82710, n82711,
         n82712, n82713, n82714, n82715, n82716, n82717, n82718, n82719,
         n82720, n82721, n82722, n82723, n82724, n82725, n82726, n82727,
         n82728, n82729, n82730, n82731, n82732, n82733, n82734, n82735,
         n82736, n82737, n82738, n82739, n82740, n82741, n82742, n82743,
         n82744, n82745, n82746, n82747, n82748, n82749, n82750, n82751,
         n82752, n82753, n82754, n82755, n82756, n82757, n82758, n82759,
         n82760, n82761, n82762, n82763, n82764, n82765, n82766, n82767,
         n82768, n82769, n82770, n82771, n82772, n82774, n82775, n82776,
         n82777, n82778, n82780, n82781, n82782, n82783, n82784, n82785,
         n82786, n82787, n82788, n82789, n82790, n82791, n82792, n82793,
         n82794, n82795, n82796, n82797, n82798, n82799, n82800, n82801,
         n82802, n82803, n82804, n82805, n82806, n82807, n82808, n82809,
         n82810, n82811, n82812, n82813, n82814, n82815, n82816, n82817,
         n82818, n82819, n82820, n82821, n82822, n82823, n82824, n82825,
         n82826, n82827, n82828, n82829, n82830, n82831, n82832, n82833,
         n82834, n82835, n82836, n82837, n82838, n82839, n82840, n82841,
         n82842, n82843, n82844, n82845, n82846, n82847, n82848, n82849,
         n82850, n82851, n82852, n82853, n82854, n82855, n82856, n82857,
         n82858, n82859, n82860, n82861, n82862, n82863, n82864, n82865,
         n82866, n82867, n82868, n82869, n82870, n82871, n82872, n82873,
         n82874, n82875, n82876, n82877, n82878, n82879, n82880, n82881,
         n82882, n82883, n82884, n82885, n82886, n82887, n82888, n82889,
         n82890, n82891, n82892, n82893, n82894, n82895, n82896, n82897,
         n82898, n82899, n82900, n82901, n82902, n82903, n82904, n82905,
         n82906, n82907, n82908, n82909, n82910, n82911, n82912, n82913,
         n82914, n82915, n82916, n82917, n82918, n82919, n82920, n82921,
         n82922, n82923, n82924, n82925, n82926, n82927, n82928, n82929,
         n82930, n82931, n82932, n82933, n82934, n82935, n82936, n82937,
         n82938, n82939, n82940, n82941, n82942, n82943, n82944, n82945,
         n82946, n82947, n82948, n82949, n82950, n82951, n82952, n82953,
         n82954, n82955, n82956, n82957, n82958, n82959, n82960, n82961,
         n82962, n82963, n82964, n82965, n82966, n82967, n82968, n82969,
         n82970, n82971, n82972, n82973, n82974, n82975, n82976, n82977,
         n82978, n82979, n82980, n82981, n82982, n82983, n82984, n82985,
         n82986, n82987, n82988, n82989, n82990, n82991, n82992, n82993,
         n82994, n82995, n82996, n82997, n82998, n82999, n83000, n83001,
         n83002, n83003, n83004, n83005, n83006, n83007, n83008, n83009,
         n83010, n83011, n83012, n83013, n83014, n83015, n83016, n83017,
         n83018, n83019, n83020, n83021, n83022, n83023, n83024, n83025,
         n83026, n83027, n83028, n83029, n83030, n83031, n83032, n83033,
         n83034, n83035, n83036, n83037, n83038, n83039, n83040, n83041,
         n83042, n83043, n83044, n83045, n83046, n83047, n83048, n83049,
         n83050, n83051, n83052, n83053, n83054, n83055, n83056, n83057,
         n83058, n83059, n83060, n83061, n83062, n83063, n83064, n83065,
         n83066, n83067, n83068, n83069, n83070, n83071, n83072, n83073,
         n83074, n83075, n83076, n83077, n83078, n83079, n83080, n83081,
         n83082, n83083, n83084, n83085, n83086, n83087, n83088, n83089,
         n83090, n83091, n83092, n83093, n83094, n83095, n83096, n83097,
         n83098, n83099, n83101, n83102, n83103, n83104, n83105, n83106,
         n83107, n83108, n83109, n83110, n83111, n83112, n83113, n83114,
         n83115, n83116, n83117, n83118, n83119, n83120, n83121, n83122,
         n83123, n83124, n83125, n83126, n83127, n83128, n83129, n83130,
         n83131, n83132, n83133, n83134, n83135, n83136, n83137, n83138,
         n83139, n83140, n83141, n83142, n83143, n83144, n83145, n83147,
         n83148, n83149, n83150, n83151, n83152, n83153, n83154, n83155,
         n83156, n83157, n83158, n83159, n83160, n83161, n83162, n83163,
         n83164, n83165, n83166, n83167, n83168, n83169, n83170, n83171,
         n83172, n83173, n83174, n83175, n83176, n83177, n83178, n83179,
         n83180, n83181, n83182, n83183, n83184, n83185, n83186, n83187,
         n83188, n83189, n83190, n83191, n83192, n83193, n83194, n83195,
         n83196, n83197, n83198, n83199, n83200, n83201, n83202, n83203,
         n83204, n83205, n83206, n83207, n83208, n83209, n83210, n83211,
         n83212, n83213, n83214, n83215, n83216, n83217, n83218, n83219,
         n83220, n83221, n83222, n83223, n83224, n83225, n83226, n83227,
         n83228, n83229, n83230, n83231, n83232, n83233, n83234, n83235,
         n83236, n83237, n83238, n83239, n83240, n83241, n83242, n83243,
         n83244, n83245, n83246, n83247, n83248, n83249, n83250, n83251,
         n83252, n83253, n83254, n83255, n83256, n83257, n83258, n83259,
         n83260, n83261, n83262, n83263, n83264, n83265, n83266, n83267,
         n83268, n83269, n83270, n83271, n83272, n83273, n83274, n83275,
         n83276, n83277, n83278, n83279, n83280, n83281, n83282, n83283,
         n83284, n83285, n83286, n83287, n83288, n83289, n83290, n83291,
         n83292, n83293, n83294, n83295, n83296, n83297, n83298, n83299,
         n83300, n83301, n83302, n83303, n83304, n83305, n83306, n83307,
         n83308, n83309, n83310, n83311, n83312, n83313, n83314, n83315,
         n83316, n83317, n83318, n83319, n83320, n83321, n83322, n83323,
         n83324, n83325, n83326, n83327, n83328, n83329, n83330, n83331,
         n83332, n83333, n83334, n83335, n83336, n83337, n83338, n83339,
         n83340, n83341, n83342, n83343, n83344, n83345, n83346, n83347,
         n83348, n83349, n83350, n83351, n83352, n83353, n83354, n83355,
         n83356, n83357, n83358, n83359, n83360, n83361, n83362, n83363,
         n83364, n83365, n83366, n83367, n83368, n83369, n83370, n83371,
         n83372, n83373, n83374, n83375, n83376, n83377, n83378, n83379,
         n83380, n83381, n83382, n83383, n83384, n83385, n83386, n83387,
         n83388, n83389, n83390, n83391, n83392, n83393, n83394, n83395,
         n83396, n83397, n83398, n83399, n83400, n83401, n83402, n83403,
         n83404, n83405, n83406, n83407, n83408, n83409, n83410, n83411,
         n83412, n83413, n83414, n83415, n83416, n83417, n83418, n83419,
         n83420, n83421, n83422, n83423, n83424, n83425, n83426, n83427,
         n83428, n83429, n83430, n83431, n83432, n83433, n83434, n83435,
         n83436, n83437, n83438, n83439, n83440, n83441, n83442, n83443,
         n83444, n83445, n83446, n83447, n83448, n83449, n83450, n83451,
         n83452, n83453, n83454, n83455, n83456, n83457, n83458, n83459,
         n83460, n83461, n83462, n83463, n83464, n83465, n83466, n83467,
         n83468, n83469, n83470, n83471, n83472, n83473, n83474, n83475,
         n83476, n83477, n83478, n83479, n83480, n83481, n83482, n83483,
         n83484, n83485, n83486, n83487, n83488, n83489, n83490, n83491,
         n83492, n83493, n83494, n83495, n83496, n83497, n83498, n83499,
         n83500, n83501, n83502, n83503, n83504, n83505, n83506, n83507,
         n83508, n83509, n83510, n83511, n83512, n83513, n83514, n83515,
         n83516, n83517, n83518, n83519, n83520, n83521, n83522, n83523,
         n83524, n83525, n83526, n83527, n83528, n83529, n83530, n83531,
         n83532, n83533, n83534, n83535, n83536, n83537, n83538, n83539,
         n83540, n83541, n83542, n83543, n83544, n83545, n83546, n83547,
         n83548, n83549, n83550, n83551, n83552, n83553, n83554, n83555,
         n83556, n83557, n83558, n83559, n83560, n83561, n83562, n83563,
         n83564, n83565, n83566, n83567, n83568, n83569, n83570, n83571,
         n83572, n83573, n83574, n83575, n83576, n83577, n83578, n83579,
         n83580, n83581, n83582, n83583, n83584, n83585, n83586, n83587,
         n83588, n83589, n83590, n83591, n83592, n83593, n83594, n83595,
         n83596, n83597, n83598, n83599, n83600, n83601, n83602, n83603,
         n83604, n83605, n83606, n83607, n83608, n83609, n83610, n83611,
         n83612, n83613, n83614, n83615, n83616, n83617, n83618, n83619,
         n83620, n83621, n83622, n83623, n83624, n83625, n83626, n83627,
         n83628, n83629, n83630, n83631, n83632, n83633, n83634, n83635,
         n83636, n83637, n83638, n83639, n83640, n83641, n83642, n83643,
         n83644, n83645, n83646, n83647, n83648, n83649, n83650, n83651,
         n83652, n83653, n83654, n83655, n83656, n83657, n83658, n83659,
         n83660, n83661, n83662, n83663, n83664, n83665, n83666, n83667,
         n83668, n83669, n83670, n83671, n83672, n83673, n83674, n83675,
         n83676, n83677, n83678, n83679, n83680, n83681, n83682, n83683,
         n83684, n83685, n83686, n83687, n83688, n83689, n83690, n83691,
         n83692, n83693, n83694, n83695, n83696, n83697, n83698, n83699,
         n83700, n83701, n83702, n83703, n83704, n83705, n83706, n83707,
         n83708, n83709, n83710, n83711, n83712, n83713, n83714, n83715,
         n83716, n83717, n83718, n83719, n83720, n83721, n83722, n83723,
         n83724, n83725, n83726, n83727, n83728, n83729, n83730, n83731,
         n83732, n83733, n83734, n83735, n83736, n83737, n83738, n83739,
         n83740, n83741, n83742, n83743, n83744, n83745, n83746, n83747,
         n83748, n83749, n83750, n83751, n83752, n83753, n83754, n83755,
         n83756, n83757, n83758, n83759, n83760, n83761, n83762, n83763,
         n83764, n83765, n83766, n83767, n83768, n83769, n83770, n83771,
         n83772, n83773, n83774, n83775, n83776, n83777, n83778, n83779,
         n83780, n83781, n83782, n83783, n83784, n83785, n83786, n83787,
         n83788, n83789, n83790, n83791, n83792, n83793, n83794, n83795,
         n83796, n83797, n83798, n83799, n83800, n83801, n83802, n83803,
         n83804, n83805, n83806, n83807, n83808, n83809, n83810, n83811,
         n83812, n83813, n83814, n83815, n83816, n83817, n83818, n83819,
         n83820, n83821, n83822, n83823, n83824, n83825, n83826, n83827,
         n83828, n83829, n83830, n83831, n83832, n83833, n83834, n83835,
         n83836, n83837, n83838, n83839, n83840, n83841, n83842, n83843,
         n83844, n83845, n83846, n83847, n83848, n83849, n83850, n83851,
         n83852, n83853, n83854, n83855, n83856, n83857, n83858, n83859,
         n83860, n83861, n83862, n83863, n83864, n83865, n83866, n83867,
         n83868, n83869, n83870, n83871, n83872, n83873, n83874, n83875,
         n83876, n83877, n83878, n83879, n83880, n83881, n83882, n83883,
         n83884, n83885, n83886, n83887, n83888, n83889, n83890, n83891,
         n83892, n83893, n83894, n83895, n83896, n83897, n83898, n83899,
         n83900, n83901, n83902, n83903, n83904, n83905, n83906, n83907,
         n83908, n83909, n83910, n83911, n83912, n83913, n83914, n83915,
         n83916, n83917, n83918, n83919, n83920, n83921, n83922, n83923,
         n83924, n83925, n83926, n83927, n83928, n83929, n83930, n83931,
         n83932, n83933, n83934, n83935, n83936, n83937, n83938, n83939,
         n83940, n83941, n83942, n83943, n83944, n83945, n83946, n83947,
         n83948, n83949, n83950, n83951, n83952, n83953, n83954, n83955,
         n83956, n83957, n83958, n83959, n83960, n83961, n83962, n83963,
         n83964, n83965, n83966, n83967, n83968, n83969, n83970, n83971,
         n83972, n83973, n83974, n83975, n83976, n83977, n83978, n83979,
         n83980, n83981, n83982, n83983, n83984, n83985, n83986, n83987,
         n83988, n83989, n83990, n83991, n83992, n83993, n83994, n83995,
         n83996, n83997, n83998, n83999, n84000, n84001, n84002, n84003,
         n84004, n84005, n84006, n84007, n84008, n84009, n84010, n84011,
         n84012, n84013, n84014, n84015, n84016, n84017, n84018, n84019,
         n84020, n84021, n84022, n84023, n84024, n84025, n84026, n84027,
         n84028, n84029, n84030, n84031, n84032, n84033, n84034, n84035,
         n84036, n84037, n84038, n84039, n84040, n84041, n84042, n84043,
         n84044, n84045, n84046, n84047, n84048, n84049, n84050, n84051,
         n84052, n84053, n84054, n84055, n84056, n84057, n84058, n84059,
         n84060, n84061, n84062, n84063, n84064, n84066, n84067, n84068,
         n84069, n84070, n84071, n84072, n84073, n84074, n84075, n84076,
         n84077, n84078, n84080, n84081, n84082, n84083, n84084, n84085,
         n84086, n84087, n84088, n84090, n84091, n84092, n84093, n84094,
         n84095, n84096, n84097, n84098, n84099, n84100, n84101, n84102,
         n84103, n84104, n84105, n84106, n84107, n84108, n84109, n84110,
         n84111, n84112, n84113, n84114, n84115, n84116, n84117, n84118,
         n84119, n84120, n84121, n84122, n84123, n84124, n84125, n84126,
         n84127, n84128, n84129, n84130, n84131, n84132, n84133, n84134,
         n84135, n84136, n84137, n84138, n84139, n84140, n84141, n84142,
         n84143, n84144, n84145, n84146, n84147, n84148, n84149, n84150,
         n84151, n84152, n84153, n84154, n84155, n84156, n84157, n84158,
         n84159, n84160, n84161, n84162, n84163, n84164, n84165, n84166,
         n84167, n84168, n84169, n84170, n84171, n84172, n84173, n84174,
         n84175, n84176, n84177, n84178, n84179, n84180, n84181, n84182,
         n84183, n84184, n84185, n84186, n84187, n84188, n84189, n84190,
         n84191, n84192, n84193, n84194, n84195, n84196, n84197, n84198,
         n84199, n84200, n84201, n84202, n84203, n84204, n84205, n84206,
         n84207, n84208, n84209, n84210, n84211, n84212, n84213, n84214,
         n84215, n84216, n84217, n84218, n84219, n84220, n84221, n84222,
         n84223, n84224, n84225, n84226, n84227, n84228, n84229, n84230,
         n84231, n84232, n84233, n84234, n84235, n84236, n84237, n84238,
         n84239, n84240, n84241, n84242, n84243, n84244, n84245, n84246,
         n84247, n84248, n84249, n84250, n84251, n84252, n84253, n84254,
         n84255, n84256, n84257, n84258, n84259, n84260, n84261, n84262,
         n84263, n84264, n84265, n84266, n84267, n84268, n84269, n84270,
         n84271, n84272, n84273, n84274, n84275, n84276, n84277, n84278,
         n84279, n84280, n84281, n84282, n84283, n84284, n84285, n84286,
         n84287, n84288, n84289, n84290, n84291, n84292, n84293, n84294,
         n84295, n84296, n84297, n84298, n84299, n84300, n84301, n84302,
         n84303, n84304, n84305, n84306, n84307, n84308, n84309, n84310,
         n84311, n84312, n84313, n84314, n84315, n84316, n84317, n84318,
         n84319, n84320, n84321, n84322, n84323, n84324, n84325, n84326,
         n84327, n84328, n84329, n84330, n84331, n84332, n84333, n84334,
         n84335, n84336, n84337, n84338, n84339, n84340, n84341, n84342,
         n84343, n84344, n84345, n84346, n84347, n84348, n84349, n84350,
         n84351, n84352, n84353, n84354, n84355, n84356, n84357, n84358,
         n84359, n84360, n84361, n84362, n84363, n84364, n84365, n84366,
         n84367, n84368, n84369, n84370, n84371, n84372, n84373, n84374,
         n84375, n84376, n84377, n84378, n84379, n84380, n84381, n84382,
         n84383, n84384, n84385, n84386, n84387, n84388, n84389, n84390,
         n84391, n84392, n84393, n84394, n84395, n84396, n84397, n84398,
         n84399, n84400, n84401, n84402, n84403, n84404, n84405, n84406,
         n84407, n84408, n84409, n84410, n84411, n84412, n84413, n84414,
         n84415, n84416, n84417, n84418, n84419, n84420, n84421, n84422,
         n84423, n84424, n84425, n84426, n84427, n84428, n84429, n84430,
         n84431, n84432, n84433, n84434, n84435, n84436, n84437, n84438,
         n84439, n84440, n84441, n84442, n84443, n84444, n84445, n84446,
         n84447, n84448, n84449, n84450, n84451, n84452, n84453, n84454,
         n84455, n84456, n84457, n84458, n84459, n84460, n84461, n84462,
         n84463, n84464, n84465, n84466, n84467, n84468, n84469, n84470,
         n84471, n84472, n84473, n84474, n84475, n84476, n84477, n84478,
         n84479, n84480, n84481, n84482, n84483, n84484, n84485, n84486,
         n84487, n84488, n84489, n84490, n84491, n84492, n84493, n84494,
         n84495, n84496, n84497, n84498, n84499, n84500, n84501, n84502,
         n84503, n84504, n84505, n84506, n84507, n84508, n84509, n84510,
         n84511, n84512, n84513, n84514, n84515, n84516, n84517, n84518,
         n84519, n84520, n84521, n84522, n84523, n84524, n84525, n84526,
         n84527, n84528, n84529, n84530, n84531, n84532, n84533, n84534,
         n84535, n84536, n84537, n84538, n84539, n84540, n84541, n84542,
         n84543, n84544, n84545, n84546, n84547, n84548, n84549, n84550,
         n84551, n84552, n84553, n84554, n84555, n84556, n84557, n84558,
         n84559, n84560, n84561, n84562, n84563, n84564, n84565, n84566,
         n84567, n84568, n84569, n84570, n84571, n84572, n84573, n84574,
         n84575, n84576, n84577, n84578, n84579, n84580, n84581, n84582,
         n84583, n84584, n84585, n84586, n84587, n84588, n84589, n84590,
         n84591, n84592, n84593, n84594, n84595, n84596, n84597, n84598,
         n84599, n84600, n84601, n84602, n84603, n84604, n84605, n84606,
         n84607, n84608, n84609, n84610, n84611, n84612, n84613, n84614,
         n84615, n84616, n84617, n84618, n84619, n84620, n84621, n84622,
         n84623, n84624, n84625, n84626, n84627, n84628, n84629, n84630,
         n84631, n84632, n84633, n84634, n84635, n84636, n84637, n84638,
         n84639, n84640, n84641, n84642, n84643, n84644, n84645, n84646,
         n84647, n84648, n84649, n84650, n84651, n84652, n84653, n84654,
         n84655, n84656, n84657, n84658, n84659, n84660, n84661, n84662,
         n84663, n84664, n84665, n84666, n84667, n84668, n84669, n84670,
         n84671, n84672, n84673, n84674, n84675, n84676, n84677, n84678,
         n84679, n84680, n84681, n84682, n84683, n84684, n84685, n84686,
         n84687, n84688, n84689, n84690, n84691, n84692, n84693, n84694,
         n84695, n84696, n84697, n84698, n84699, n84700, n84701, n84702,
         n84703, n84704, n84705, n84706, n84707, n84708, n84709, n84710,
         n84711, n84712, n84713, n84714, n84715, n84716, n84717, n84718,
         n84719, n84720, n84721, n84722, n84723, n84724, n84725, n84726,
         n84727, n84728, n84729, n84730, n84731, n84732, n84733, n84734,
         n84735, n84736, n84737, n84738, n84739, n84740, n84741, n84742,
         n84743, n84744, n84745, n84746, n84747, n84748, n84749, n84750,
         n84751, n84752, n84753, n84754, n84755, n84756, n84757, n84758,
         n84759, n84760, n84761, n84762, n84763, n84764, n84765, n84766,
         n84767, n84768, n84769, n84770, n84771, n84772, n84773, n84774,
         n84775, n84776, n84777, n84778, n84779, n84780, n84781, n84782,
         n84783, n84784, n84785, n84786, n84787, n84788, n84789, n84790,
         n84791, n84792, n84793, n84794, n84795, n84796, n84797, n84798,
         n84799, n84800, n84801, n84802, n84803, n84804, n84805, n84806,
         n84807, n84808, n84809, n84810, n84811, n84812, n84813, n84814,
         n84815, n84816, n84817, n84818, n84819, n84820, n84821, n84822,
         n84823, n84824, n84825, n84826, n84827, n84828, n84829, n84830,
         n84831, n84832, n84833, n84834, n84835, n84836, n84837, n84838,
         n84839, n84840, n84841, n84842, n84843, n84844, n84845, n84846,
         n84847, n84848, n84849, n84850, n84851, n84852, n84853, n84854,
         n84855, n84856, n84857, n84858, n84859, n84860, n84861, n84862,
         n84863, n84864, n84865, n84866, n84867, n84868, n84869, n84870,
         n84871, n84872, n84873, n84874, n84875, n84876, n84877, n84878,
         n84879, n84880, n84881, n84882, n84883, n84884, n84885, n84886,
         n84887, n84888, n84889, n84890, n84891, n84892, n84893, n84894,
         n84895, n84896, n84897, n84898, n84899, n84900, n84901, n84902,
         n84903, n84904, n84905, n84906, n84907, n84908, n84909, n84910,
         n84911, n84912, n84913, n84914, n84915, n84916, n84917, n84918,
         n84919, n84920, n84921, n84922, n84923, n84924, n84925, n84926,
         n84927, n84928, n84929, n84930, n84931, n84932, n84933, n84934,
         n84935, n84936, n84937, n84938, n84939, n84940, n84941, n84942,
         n84943, n84944, n84945, n84946, n84947, n84948, n84949, n84950,
         n84951, n84952, n84953, n84954, n84955, n84956, n84957, n84958,
         n84959, n84960, n84961, n84962, n84963, n84964, n84965, n84966,
         n84967, n84968, n84969, n84970, n84971, n84972, n84973, n84974,
         n84975, n84976, n84977, n84978, n84979, n84980, n84981, n84982,
         n84983, n84984, n84985, n84986, n84987, n84988, n84989, n84990,
         n84991, n84992, n84993, n84994, n84995, n84996, n84997, n84998,
         n84999, n85000, n85001, n85002, n85003, n85004, n85005, n85006,
         n85007, n85008, n85009, n85010, n85011, n85012, n85013, n85014,
         n85015, n85016, n85017, n85018, n85019, n85020, n85021, n85022,
         n85023, n85024, n85025, n85026, n85027, n85028, n85029, n85030,
         n85031, n85032, n85033, n85034, n85035, n85036, n85037, n85038,
         n85039, n85040, n85041, n85042, n85043, n85044, n85045, n85046,
         n85047, n85048, n85049, n85050, n85051, n85052, n85053, n85054,
         n85055, n85056, n85057, n85058, n85059, n85060, n85061, n85062,
         n85063, n85064, n85065, n85066, n85067, n85068, n85069, n85070,
         n85071, n85072, n85073, n85074, n85075, n85076, n85077, n85078,
         n85079, n85080, n85081, n85082, n85083, n85084, n85085, n85086,
         n85087, n85088, n85089, n85090, n85091, n85092, n85093, n85094,
         n85095, n85096, n85097, n85098, n85099, n85100, n85101, n85102,
         n85103, n85104, n85105, n85106, n85107, n85108, n85109, n85110,
         n85111, n85112, n85113, n85114, n85115, n85116, n85117, n85118,
         n85119, n85120, n85121, n85122, n85123, n85124, n85125, n85126,
         n85127, n85128, n85129, n85130, n85131, n85132, n85133, n85134,
         n85135, n85136, n85137, n85138, n85139, n85140, n85141, n85142,
         n85143, n85144, n85145, n85146, n85147, n85148, n85149, n85150,
         n85151, n85152, n85153, n85154, n85155, n85156, n85157, n85158,
         n85159, n85160, n85161, n85162, n85163, n85164, n85165, n85166,
         n85167, n85168, n85169, n85170, n85171, n85172, n85173, n85174,
         n85175, n85176, n85177, n85178, n85179, n85180, n85181, n85182,
         n85183, n85184, n85185, n85186, n85187, n85188, n85189, n85190,
         n85191, n85192, n85193, n85194, n85195, n85196, n85197, n85198,
         n85199, n85200, n85201, n85202, n85205, n85206, n85207, n85208,
         n85210, n85211, n85212, n85213, n85214, n85215, n85216, n85217,
         n85218, n85219, n85220, n85221, n85222, n85223, n85224, n85225,
         n85226, n85227, n85228, n85229, n85230, n85231, n85232, n85233,
         n85234, n85235, n85236, n85237, n85238, n85239, n85240, n85241,
         n85242, n85243, n85244, n85245, n85246, n85247, n85248, n85249,
         n85250, n85251, n85252, n85253, n85254, n85255, n85256, n85257,
         n85258, n85259, n85260, n85261, n85262, n85263, n85264, n85265,
         n85266, n85267, n85268, n85269, n85270, n85271, n85272, n85273,
         n85274, n85275, n85276, n85277, n85278, n85279, n85280, n85281,
         n85282, n85283, n85284, n85285, n85286, n85287, n85288, n85289,
         n85290, n85291, n85292, n85293, n85294, n85295, n85296, n85297,
         n85298, n85299, n85300, n85301, n85302, n85303, n85304, n85305,
         n85306, n85307, n85308, n85309, n85310, n85311, n85312, n85313,
         n85314, n85315, n85316, n85317, n85318, n85319, n85320, n85321,
         n85322, n85323, n85324, n85325, n85326, n85327, n85328, n85329,
         n85330, n85331, n85332, n85333, n85334, n85335, n85336, n85337,
         n85338, n85339, n85340, n85341, n85342, n85343, n85344, n85345,
         n85346, n85347, n85348, n85349, n85350, n85351, n85352, n85353,
         n85354, n85355, n85356, n85357, n85358, n85359, n85360, n85361,
         n85362, n85363, n85364, n85365, n85366, n85367, n85368, n85369,
         n85370, n85371, n85372, n85373, n85374, n85375, n85376, n85377,
         n85378, n85379, n85380, n85381, n85382, n85383, n85384, n85385,
         n85386, n85387, n85388, n85389, n85390, n85391, n85392, n85393,
         n85394, n85395, n85396, n85397, n85398, n85399, n85400, n85401,
         n85402, n85403, n85404, n85405, n85406, n85407, n85408, n85409,
         n85410, n85411, n85412, n85413, n85414, n85415, n85416, n85417,
         n85418, n85419, n85420, n85421, n85422, n85423, n85424, n85425,
         n85426, n85427, n85428, n85429, n85430, n85431, n85432, n85433,
         n85434, n85435, n85436, n85437, n85438, n85439, n85440, n85441,
         n85442, n85443, n85444, n85445, n85446, n85447, n85448, n85449,
         n85450, n85451, n85452, n85453, n85454, n85455, n85456, n85457,
         n85458, n85459, n85460, n85461, n85462, n85463, n85464, n85465,
         n85466, n85467, n85468, n85469, n85470, n85471, n85472, n85473,
         n85474, n85475, n85476, n85477, n85478, n85479, n85480, n85481,
         n85482, n85483, n85484, n85485, n85486, n85487, n85488, n85489,
         n85490, n85491, n85492, n85493, n85494, n85495, n85496, n85497,
         n85498, n85499, n85500, n85501, n85502, n85503, n85504, n85505,
         n85506, n85507, n85508, n85509, n85510, n85511, n85512, n85513,
         n85514, n85515, n85516, n85517, n85518, n85519, n85520, n85521,
         n85522, n85523, n85524, n85525, n85526, n85527, n85528, n85529,
         n85530, n85531, n85532, n85533, n85534, n85535, n85536, n85537,
         n85538, n85539, n85540, n85541, n85542, n85543, n85544, n85545,
         n85546, n85547, n85548, n85549, n85550, n85551, n85552, n85553,
         n85554, n85555, n85556, n85557, n85558, n85559, n85560, n85561,
         n85562, n85563, n85564, n85565, n85566, n85567, n85568, n85569,
         n85570, n85571, n85572, n85573, n85574, n85575, n85576, n85577,
         n85578, n85579, n85580, n85581, n85582, n85583, n85584, n85585,
         n85586, n85587, n85588, n85589, n85590, n85591, n85592, n85593,
         n85594, n85595, n85596, n85597, n85598, n85599, n85600, n85601,
         n85602, n85603, n85604, n85605, n85606, n85607, n85608, n85609,
         n85610, n85611, n85612, n85613, n85614, n85615, n85616, n85617,
         n85618, n85619, n85620, n85621, n85622, n85623, n85624, n85625,
         n85626, n85627, n85628, n85629, n85630, n85631, n85632, n85633,
         n85634, n85635, n85636, n85637, n85638, n85639, n85640, n85641,
         n85642, n85643, n85644, n85645, n85646, n85647, n85648, n85649,
         n85650, n85651, n85652, n85653, n85654, n85655, n85656, n85657,
         n85658, n85659, n85660, n85661, n85662, n85663, n85664, n85665,
         n85666, n85667, n85668, n85669, n85670, n85671, n85672, n85673,
         n85674, n85675, n85676, n85677, n85678, n85679, n85680, n85681,
         n85682, n85683, n85684, n85685, n85686, n85687, n85688, n85689,
         n85690, n85691, n85692, n85693, n85694, n85695, n85696, n85697,
         n85698, n85699, n85700, n85701, n85702, n85703, n85704, n85705,
         n85706, n85707, n85708, n85709, n85710, n85711, n85712, n85713,
         n85714, n85715, n85716, n85717, n85718, n85719, n85720, n85721,
         n85722, n85723, n85724, n85725, n85726, n85727, n85728, n85729,
         n85730, n85731, n85732, n85733, n85734, n85735, n85736, n85737,
         n85738, n85739, n85740, n85741, n85742, n85743, n85744, n85745,
         n85746, n85747, n85748, n85749, n85750, n85751, n85752, n85753,
         n85754, n85755, n85756, n85757, n85758, n85759, n85760, n85761,
         n85762, n85763, n85764, n85765, n85766, n85767, n85768, n85769,
         n85770, n85771, n85772, n85773, n85774, n85775, n85776, n85777,
         n85778, n85779, n85780, n85781, n85782, n85783, n85784, n85785,
         n85786, n85787, n85788, n85789, n85790, n85791, n85792, n85793,
         n85794, n85795, n85796, n85797, n85798, n85799, n85800, n85801,
         n85802, n85803, n85804, n85805, n85806, n85807, n85808, n85809,
         n85810, n85811, n85812, n85813, n85814, n85815, n85816, n85817,
         n85818, n85819, n85820, n85821, n85822, n85823, n85824, n85825,
         n85826, n85827, n85828, n85829, n85830, n85831, n85832, n85833,
         n85834, n85835, n85836, n85837, n85838, n85839, n85840, n85841,
         n85842, n85843, n85844, n85845, n85846, n85847, n85848, n85849,
         n85850, n85851, n85852, n85853, n85854, n85855, n85856, n85857,
         n85858, n85859, n85860, n85861, n85862, n85863, n85864, n85865,
         n85866, n85867, n85868, n85869, n85870, n85871, n85872, n85873,
         n85874, n85875, n85876, n85877, n85878, n85879, n85880, n85881,
         n85882, n85883, n85884, n85885, n85886, n85887, n85888, n85889,
         n85890, n85891, n85892, n85893, n85894, n85895, n85896, n85897,
         n85898, n85899, n85900, n85901, n85902, n85903, n85904, n85905,
         n85906, n85907, n85908, n85909, n85910, n85911, n85912, n85913,
         n85914, n85915, n85916, n85917, n85918, n85919, n85920, n85921,
         n85922, n85923, n85924, n85925, n85926, n85927, n85928, n85929,
         n85930, n85931, n85932, n85933, n85934, n85935, n85936, n85937,
         n85938, n85939, n85940, n85941, n85942, n85943, n85944, n85945,
         n85946, n85947, n85948, n85949, n85950, n85951, n85952, n85953,
         n85954, n85955, n85956, n85957, n85958, n85959, n85960, n85961,
         n85962, n85963, n85964, n85965, n85966, n85967, n85968, n85969,
         n85970, n85971, n85972, n85973, n85974, n85975, n85976, n85977,
         n85978, n85979, n85980, n85981, n85982, n85983, n85984, n85985,
         n85986, n85987, n85988, n85989, n85990, n85991, n85992, n85993,
         n85994, n85995, n85996, n85997, n85998, n85999, n86000, n86001,
         n86002, n86003, n86004, n86005, n86006, n86007, n86008, n86009,
         n86010, n86011, n86012, n86013, n86014, n86015, n86016, n86017,
         n86018, n86019, n86020, n86021, n86022, n86023, n86024, n86025,
         n86026, n86027, n86028, n86029, n86030, n86031, n86032, n86033,
         n86034, n86035, n86036, n86037, n86038, n86039, n86040, n86041,
         n86042, n86043, n86044, n86045, n86046, n86047, n86048, n86049,
         n86050, n86051, n86052, n86053, n86054, n86055, n86056, n86057,
         n86058, n86059, n86060, n86061, n86062, n86063, n86064, n86065,
         n86066, n86067, n86068, n86069, n86070, n86071, n86072, n86073,
         n86074, n86075, n86076, n86077, n86078, n86079, n86080, n86081,
         n86082, n86083, n86084, n86085, n86086, n86087, n86088, n86089,
         n86090, n86091, n86092, n86093, n86094, n86095, n86096, n86097,
         n86098, n86099, n86100, n86101, n86102, n86103, n86104, n86105,
         n86106, n86107, n86108, n86109, n86110, n86111, n86112, n86113,
         n86114, n86115, n86116, n86117, n86118, n86119, n86120, n86121,
         n86122, n86123, n86124, n86125, n86126, n86127, n86128, n86129,
         n86130, n86131, n86132, n86133, n86134, n86135, n86136, n86137,
         n86138, n86139, n86140, n86141, n86142, n86143, n86144, n86145,
         n86146, n86147, n86148, n86149, n86150, n86151, n86152, n86153,
         n86154, n86155, n86156, n86157, n86158, n86159, n86160, n86161,
         n86162, n86163, n86164, n86165, n86166, n86167, n86168, n86169,
         n86170, n86171, n86172, n86173, n86174, n86175, n86176, n86177,
         n86178, n86179, n86180, n86181, n86182, n86183, n86184, n86185,
         n86186, n86187, n86188, n86189, n86190, n86191, n86192, n86193,
         n86194, n86196, n86197, n86198, n86199, n86200, n86201, n86202,
         n86203, n86204, n86205, n86206, n86207, n86208, n86209, n86210,
         n86211, n86212, n86213, n86214, n86215, n86216, n86217, n86218,
         n86219, n86220, n86221, n86222, n86223, n86224, n86225, n86226,
         n86228, n86229, n86230, n86231, n86232, n86233, n86234, n86235,
         n86236, n86237, n86238, n86239, n86240, n86241, n86242, n86243,
         n86244, n86245, n86246, n86247, n86248, n86249, n86250, n86251,
         n86252, n86253, n86254, n86255, n86256, n86257, n86258, n86259,
         n86260, n86261, n86262, n86263, n86264, n86265, n86266, n86267,
         n86268, n86269, n86270, n86271, n86272, n86273, n86274, n86275,
         n86276, n86277, n86278, n86279, n86280, n86281, n86282, n86283,
         n86284, n86285, n86286, n86287, n86288, n86289, n86290, n86291,
         n86292, n86293, n86294, n86295, n86296, n86297, n86298, n86299,
         n86300, n86301, n86302, n86303, n86304, n86305, n86306, n86307,
         n86308, n86309, n86310, n86311, n86312, n86313, n86314, n86315,
         n86316, n86317, n86318, n86319, n86320, n86321, n86322, n86323,
         n86324, n86325, n86326, n86327, n86328, n86329, n86330, n86331,
         n86332, n86333, n86334, n86335, n86336, n86337, n86338, n86339,
         n86340, n86341, n86342, n86343, n86344, n86345, n86346, n86347,
         n86348, n86349, n86350, n86351, n86352, n86353, n86354, n86355,
         n86356, n86357, n86358, n86359, n86360, n86361, n86362, n86363,
         n86364, n86365, n86366, n86367, n86368, n86369, n86370, n86371,
         n86372, n86373, n86374, n86375, n86376, n86377, n86378, n86379,
         n86380, n86381, n86382, n86383, n86384, n86385, n86386, n86387,
         n86388, n86389, n86390, n86391, n86392, n86393, n86394, n86395,
         n86396, n86397, n86398, n86399, n86400, n86401, n86402, n86403,
         n86404, n86405, n86406, n86407, n86408, n86409, n86410, n86411,
         n86412, n86413, n86414, n86415, n86416, n86417, n86418, n86419,
         n86420, n86421, n86422, n86423, n86424, n86425, n86426, n86427,
         n86428, n86429, n86430, n86431, n86432, n86433, n86434, n86435,
         n86436, n86437, n86438, n86439, n86440, n86441, n86442, n86443,
         n86444, n86445, n86446, n86447, n86448, n86449, n86450, n86451,
         n86452, n86453, n86454, n86455, n86456, n86457, n86458, n86459,
         n86460, n86461, n86462, n86463, n86464, n86465, n86466, n86467,
         n86468, n86469, n86470, n86471, n86472, n86473, n86474, n86475,
         n86476, n86477, n86478, n86479, n86480, n86481, n86482, n86483,
         n86484, n86485, n86486, n86487, n86488, n86489, n86490, n86491,
         n86492, n86493, n86494, n86495, n86496, n86497, n86498, n86499,
         n86500, n86501, n86502, n86503, n86504, n86505, n86506, n86507,
         n86508, n86509, n86510, n86511, n86512, n86513, n86514, n86515,
         n86516, n86517, n86518, n86519, n86520, n86521, n86522, n86523,
         n86524, n86525, n86526, n86527, n86528, n86529, n86530, n86531,
         n86532, n86533, n86534, n86535, n86536, n86537, n86538, n86539,
         n86540, n86541, n86542, n86543, n86544, n86545, n86546, n86547,
         n86548, n86549, n86550, n86551, n86552, n86553, n86554, n86555,
         n86556, n86557, n86558, n86559, n86560, n86561, n86562, n86563,
         n86564, n86565, n86566, n86567, n86568, n86569, n86570, n86571,
         n86572, n86573, n86574, n86575, n86576, n86577, n86578, n86579,
         n86580, n86581, n86582, n86583, n86584, n86585, n86586, n86587,
         n86588, n86589, n86590, n86591, n86592, n86593, n86594, n86595,
         n86596, n86597, n86598, n86599, n86600, n86601, n86602, n86603,
         n86604, n86605, n86606, n86607, n86608, n86609, n86610, n86611,
         n86612, n86613, n86614, n86615, n86616, n86617, n86618, n86619,
         n86620, n86621, n86622, n86623, n86624, n86625, n86626, n86627,
         n86628, n86629, n86630, n86631, n86632, n86633, n86634, n86635,
         n86636, n86637, n86638, n86639, n86640, n86641, n86642, n86643,
         n86644, n86645, n86646, n86647, n86648, n86649, n86650, n86651,
         n86652, n86653, n86654, n86655, n86656, n86657, n86658, n86659,
         n86660, n86661, n86662, n86663, n86664, n86665, n86666, n86667,
         n86668, n86669, n86670, n86671, n86672, n86673, n86674, n86675,
         n86676, n86677, n86678, n86679, n86680, n86681, n86682, n86683,
         n86684, n86685, n86686, n86687, n86688, n86689, n86690, n86691,
         n86692, n86693, n86694, n86695, n86696, n86697, n86698, n86699,
         n86700, n86701, n86702, n86703, n86704, n86705, n86706, n86707,
         n86708, n86709, n86710, n86711, n86712, n86713, n86714, n86715,
         n86716, n86717, n86718, n86719, n86720, n86721, n86722, n86723,
         n86724, n86725, n86726, n86727, n86728, n86729, n86730, n86731,
         n86732, n86733, n86734, n86735, n86736, n86737, n86738, n86739,
         n86740, n86741, n86742, n86743, n86744, n86745, n86746, n86747,
         n86748, n86749, n86750, n86751, n86752, n86753, n86754, n86755,
         n86756, n86757, n86758, n86759, n86760, n86761, n86762, n86763,
         n86764, n86765, n86766, n86767, n86768, n86769, n86770, n86771,
         n86772, n86773, n86774, n86775, n86776, n86777, n86778, n86779,
         n86780, n86781, n86782, n86783, n86784, n86785, n86786, n86787,
         n86788, n86789, n86790, n86791, n86792, n86793, n86794, n86795,
         n86796, n86797, n86798, n86799, n86800, n86801, n86802, n86803,
         n86804, n86805, n86806, n86807, n86808, n86809, n86810, n86811,
         n86812, n86813, n86814, n86815, n86816, n86817, n86818, n86819,
         n86820, n86821, n86822, n86823, n86824, n86825, n86826, n86827,
         n86828, n86829, n86830, n86831, n86832, n86833, n86834, n86835,
         n86836, n86837, n86838, n86839, n86840, n86841, n86842, n86843,
         n86844, n86845, n86846, n86847, n86848, n86849, n86850, n86851,
         n86852, n86853, n86854, n86855, n86856, n86857, n86858, n86859,
         n86860, n86861, n86862, n86863, n86864, n86865, n86866, n86867,
         n86868, n86869, n86870, n86871, n86872, n86873, n86874, n86875,
         n86876, n86877, n86878, n86879, n86880, n86881, n86882, n86883,
         n86884, n86885, n86886, n86887, n86888, n86889, n86890, n86891,
         n86892, n86893, n86894, n86895, n86896, n86897, n86898, n86899,
         n86900, n86901, n86902, n86903, n86904, n86905, n86906, n86907,
         n86908, n86909, n86910, n86911, n86912, n86913, n86914, n86915,
         n86916, n86917, n86918, n86919, n86920, n86921, n86922, n86923,
         n86924, n86925, n86926, n86927, n86928, n86929, n86930, n86931,
         n86932, n86933, n86934, n86935, n86936, n86937, n86938, n86939,
         n86940, n86941, n86942, n86943, n86944, n86945, n86946, n86947,
         n86948, n86949, n86950, n86951, n86952, n86953, n86954, n86955,
         n86956, n86957, n86958, n86959, n86960, n86961, n86962, n86963,
         n86964, n86965, n86966, n86967, n86968, n86969, n86970, n86971,
         n86972, n86973, n86974, n86975, n86976, n86977, n86978, n86979,
         n86980, n86981, n86982, n86983, n86984, n86985, n86986, n86987,
         n86988, n86989, n86990, n86991, n86992, n86993, n86994, n86995,
         n86996, n86997, n86998, n86999, n87000, n87001, n87002, n87003,
         n87004, n87005, n87006, n87007, n87008, n87009, n87010, n87011,
         n87012, n87013, n87014, n87015, n87016, n87017, n87018, n87019,
         n87020, n87021, n87022, n87023, n87024, n87025, n87026, n87027,
         n87028, n87029, n87030, n87031, n87032, n87033, n87034, n87035,
         n87036, n87037, n87038, n87039, n87040, n87041, n87042, n87043,
         n87044, n87045, n87046, n87047, n87048, n87049, n87050, n87051,
         n87052, n87053, n87054, n87055, n87056, n87057, n87058, n87059,
         n87060, n87061, n87062, n87063, n87064, n87065, n87066, n87067,
         n87068, n87069, n87070, n87071, n87072, n87073, n87074, n87075,
         n87076, n87077, n87078, n87079, n87080, n87081, n87082, n87083,
         n87084, n87085, n87086, n87087, n87088, n87089, n87090, n87091,
         n87092, n87093, n87094, n87095, n87096, n87097, n87098, n87099,
         n87100, n87101, n87102, n87103, n87104, n87105, n87106, n87107,
         n87108, n87109, n87110, n87111, n87112, n87113, n87114, n87115,
         n87116, n87117, n87118, n87119, n87120, n87121, n87122, n87123,
         n87124, n87125, n87126, n87127, n87128, n87129, n87130, n87131,
         n87132, n87133, n87134, n87135, n87136, n87137, n87138, n87139,
         n87140, n87141, n87142, n87143, n87144, n87145, n87146, n87147,
         n87148, n87149, n87150, n87151, n87152, n87153, n87154, n87155,
         n87156, n87157, n87158, n87159, n87160, n87161, n87162, n87163,
         n87164, n87165, n87166, n87167, n87168, n87169, n87170, n87171,
         n87172, n87173, n87174, n87175, n87176, n87177, n87178, n87179,
         n87180, n87181, n87182, n87183, n87184, n87185, n87186, n87187,
         n87188, n87189, n87190, n87191, n87192, n87193, n87194, n87195,
         n87196, n87197, n87198, n87199, n87200, n87201, n87202, n87203,
         n87204, n87205, n87206, n87207, n87208, n87209, n87210, n87211,
         n87212, n87213, n87214, n87215, n87216, n87217, n87218, n87219,
         n87220, n87221, n87222, n87223, n87224, n87225, n87226, n87227,
         n87228, n87229, n87230, n87231, n87232, n87233, n87234, n87235,
         n87236, n87237, n87238, n87239, n87240, n87241, n87242, n87243,
         n87244, n87245, n87246, n87247, n87248, n87249, n87250, n87251,
         n87252, n87253, n87254, n87255, n87256, n87257, n87258, n87259,
         n87260, n87261, n87262, n87263, n87264, n87265, n87266, n87267,
         n87268, n87269, n87270, n87271, n87272, n87273, n87274, n87275,
         n87276, n87277, n87278, n87279, n87280, n87281, n87282, n87283,
         n87284, n87285, n87286, n87287, n87288, n87289, n87290, n87291,
         n87292, n87293, n87294, n87295, n87296, n87297, n87298, n87299,
         n87300, n87301, n87302, n87303, n87304, n87305, n87306, n87307,
         n87308, n87309, n87310, n87311, n87312, n87313, n87314, n87315,
         n87316, n87317, n87318, n87319, n87320, n87321, n87322, n87323,
         n87324, n87325, n87326, n87327, n87328, n87329, n87330, n87331,
         n87332, n87333, n87334, n87335, n87336, n87337, n87338, n87339,
         n87340, n87341, n87342, n87343, n87344, n87345, n87346, n87347,
         n87348, n87349, n87350, n87351, n87352, n87353, n87354, n87355,
         n87356, n87357, n87358, n87359, n87360, n87361, n87362, n87363,
         n87364, n87365, n87366, n87367, n87368, n87369, n87370, n87371,
         n87372, n87373, n87374, n87375, n87376, n87377, n87378, n87379,
         n87380, n87381, n87382, n87383, n87384, n87385, n87386, n87387,
         n87388, n87389, n87390, n87391, n87392, n87393, n87394, n87395,
         n87396, n87397, n87398, n87399, n87400, n87401, n87402, n87403,
         n87404, n87405, n87406, n87407, n87408, n87409, n87410, n87411,
         n87412, n87413, n87414, n87415, n87416, n87417, n87418, n87419,
         n87420, n87421, n87422, n87423, n87424, n87425, n87426, n87427,
         n87428, n87429, n87430, n87431, n87432, n87433, n87434, n87435,
         n87436, n87437, n87438, n87439, n87440, n87441, n87442, n87443,
         n87444, n87445, n87446, n87447, n87448, n87449, n87450, n87451,
         n87452, n87453, n87454, n87455, n87456, n87457, n87458, n87459,
         n87460, n87461, n87462, n87463, n87464, n87465, n87466, n87467,
         n87468, n87469, n87470, n87471, n87472, n87473, n87474, n87475,
         n87476, n87477, n87478, n87479, n87480, n87481, n87482, n87483,
         n87484, n87485, n87486, n87487, n87488, n87489, n87490, n87491,
         n87492, n87493, n87494, n87495, n87496, n87497, n87498, n87499,
         n87500, n87501, n87502, n87503, n87504, n87505, n87506, n87507,
         n87508, n87509, n87510, n87511, n87512, n87513, n87514, n87515,
         n87516, n87517, n87518, n87519, n87520, n87521, n87522, n87523,
         n87524, n87525, n87526, n87527, n87528, n87529, n87530, n87531,
         n87532, n87533, n87534, n87535, n87536, n87537, n87538, n87539,
         n87540, n87541, n87542, n87543, n87544, n87545, n87546, n87547,
         n87548, n87549, n87550, n87551, n87552, n87553, n87554, n87555,
         n87556, n87557, n87558, n87559, n87560, n87561, n87562, n87563,
         n87564, n87565, n87566, n87567, n87568, n87569, n87570, n87571,
         n87572, n87573, n87574, n87575, n87576, n87577, n87578, n87579,
         n87580, n87581, n87582, n87583, n87584, n87585, n87586, n87587,
         n87588, n87589, n87590, n87591, n87592, n87593, n87594, n87595,
         n87596, n87597, n87598, n87599, n87600, n87601, n87602, n87603,
         n87604, n87605, n87606, n87607, n87608, n87609, n87610, n87611,
         n87612, n87613, n87614, n87615, n87616, n87617, n87618, n87619,
         n87620, n87621, n87622, n87623, n87624, n87625, n87626, n87627,
         n87628, n87629, n87630, n87631, n87632, n87633, n87634, n87635,
         n87636, n87637, n87638, n87639, n87640, n87641, n87642, n87643,
         n87644, n87645, n87646, n87647, n87648, n87649, n87650, n87651,
         n87652, n87653, n87654, n87655, n87656, n87657, n87658, n87659,
         n87660, n87661, n87662, n87663, n87664, n87665, n87666, n87667,
         n87668, n87669, n87670, n87671, n87672, n87673, n87674, n87675,
         n87676, n87677, n87678, n87679, n87680, n87681, n87682, n87683,
         n87684, n87685, n87686, n87687, n87688, n87689, n87690, n87691,
         n87692, n87693, n87694, n87695, n87696, n87697, n87698, n87699,
         n87700, n87701, n87702, n87703, n87704, n87705, n87706, n87707,
         n87708, n87709, n87710, n87711, n87712, n87713, n87714, n87715,
         n87716, n87717, n87718, n87719, n87720, n87721, n87722, n87723,
         n87724, n87725, n87726, n87727, n87728, n87729, n87730, n87731,
         n87732, n87733, n87734, n87735, n87736, n87737, n87738, n87739,
         n87740, n87741, n87742, n87743, n87744, n87745, n87746, n87747,
         n87748, n87749, n87750, n87751, n87752, n87753, n87754, n87755,
         n87756, n87757, n87758, n87759, n87760, n87761, n87762, n87763,
         n87764, n87765, n87766, n87767, n87768, n87769, n87770, n87771,
         n87772, n87773, n87774, n87775, n87776, n87777, n87778, n87779,
         n87780, n87781, n87782, n87783, n87784, n87785, n87786, n87787,
         n87788, n87789, n87790, n87791, n87792, n87793, n87794, n87795,
         n87796, n87797, n87798, n87799, n87800, n87801, n87802, n87803,
         n87804, n87805, n87806, n87807, n87808, n87809, n87810, n87811,
         n87812, n87813, n87814, n87815, n87816, n87817, n87818, n87819,
         n87820, n87821, n87822, n87823, n87824, n87825, n87826, n87827,
         n87828, n87829, n87830, n87831, n87832, n87833, n87834, n87835,
         n87836, n87837, n87838, n87839, n87840, n87841, n87842, n87843,
         n87844, n87845, n87846, n87847, n87848, n87849, n87850, n87851,
         n87852, n87853, n87854, n87855, n87856, n87857, n87858, n87859,
         n87860, n87861, n87862, n87863, n87864, n87865, n87866, n87867,
         n87868, n87869, n87870, n87871, n87872, n87873, n87874, n87875,
         n87876, n87877, n87878, n87879, n87880, n87881, n87882, n87883,
         n87884, n87885, n87886, n87887, n87888, n87889, n87890, n87891,
         n87892, n87893, n87894, n87895, n87896, n87897, n87898, n87899,
         n87900, n87901, n87902, n87903, n87904, n87905, n87906, n87907,
         n87908, n87909, n87910, n87911, n87912, n87913, n87914, n87915,
         n87916, n87917, n87918, n87919, n87920, n87921, n87922, n87923,
         n87924, n87925, n87926, n87927, n87928, n87929, n87930, n87931,
         n87932, n87933, n87934, n87935, n87936, n87937, n87938, n87939,
         n87940, n87941, n87942, n87943, n87944, n87945, n87946, n87947,
         n87948, n87949, n87950, n87951, n87952, n87953, n87954, n87955,
         n87956, n87957, n87958, n87959, n87960, n87961, n87962, n87963,
         n87964, n87965, n87966, n87967, n87968, n87969, n87970, n87971,
         n87972, n87973, n87974, n87975, n87976, n87977, n87978, n87979,
         n87980, n87981, n87982, n87983, n87984, n87985, n87986, n87987,
         n87988, n87989, n87990, n87991, n87992, n87993, n87994, n87995,
         n87996, n87997, n87998, n87999, n88000, n88001, n88002, n88003,
         n88004, n88005, n88006, n88007, n88008, n88009, n88010, n88011,
         n88012, n88013, n88014, n88015, n88016, n88017, n88018, n88019,
         n88020, n88021, n88022, n88023, n88024, n88025, n88026, n88027,
         n88028, n88029, n88030, n88031, n88032, n88033, n88034, n88035,
         n88036, n88037, n88038, n88039, n88040, n88041, n88042, n88043,
         n88044, n88045, n88046, n88047, n88048, n88049, n88050, n88051,
         n88052, n88053, n88054, n88055, n88056, n88057, n88058, n88059,
         n88060, n88061, n88062, n88063, n88064, n88065, n88066, n88067,
         n88068, n88069, n88070, n88071, n88072, n88073, n88074, n88075,
         n88076, n88077, n88078, n88079, n88080, n88081, n88082, n88083,
         n88084, n88085, n88086, n88087, n88088, n88089, n88090, n88091,
         n88092, n88093, n88094, n88095, n88096, n88097, n88098, n88099,
         n88100, n88101, n88102, n88103, n88104, n88105, n88106, n88107,
         n88108, n88109, n88110, n88111, n88112, n88113, n88114, n88115,
         n88116, n88117, n88118, n88119, n88120, n88121, n88122, n88123,
         n88124, n88125, n88126, n88127, n88128, n88129, n88130, n88131,
         n88132, n88133, n88134, n88135, n88136, n88137, n88138, n88139,
         n88140, n88141, n88142, n88143, n88144, n88145, n88146, n88147,
         n88148, n88149, n88150, n88151, n88152, n88153, n88154, n88155,
         n88156, n88157, n88158, n88159, n88160, n88161, n88162, n88163,
         n88164, n88165, n88166, n88167, n88168, n88169, n88170, n88171,
         n88172, n88173, n88174, n88175, n88176, n88177, n88178, n88179,
         n88180, n88181, n88182, n88183, n88184, n88185, n88186, n88187,
         n88188, n88189, n88190, n88191, n88192, n88193, n88194, n88195,
         n88196, n88197, n88198, n88199, n88200, n88201, n88202, n88203,
         n88204, n88205, n88206, n88207, n88208, n88209, n88210, n88211,
         n88212, n88213, n88214, n88215, n88216, n88217, n88218, n88219,
         n88220, n88221, n88222, n88223, n88224, n88225, n88226, n88227,
         n88228, n88229, n88230, n88231, n88232, n88233, n88234, n88235,
         n88236, n88237, n88238, n88239, n88240, n88241, n88242, n88243,
         n88244, n88245, n88246, n88247, n88248, n88249, n88250, n88251,
         n88252, n88253, n88254, n88255, n88256, n88257, n88258, n88259,
         n88260, n88261, n88262, n88263, n88264, n88265, n88266, n88267,
         n88268, n88269, n88270, n88271, n88272, n88273, n88274, n88275,
         n88276, n88277, n88278, n88279, n88280, n88281, n88282, n88283,
         n88284, n88285, n88286, n88287, n88288, n88289, n88290, n88291,
         n88292, n88293, n88294, n88295, n88296, n88297, n88298, n88299,
         n88300, n88301, n88302, n88303, n88304, n88305, n88306, n88307,
         n88308, n88309, n88310, n88311, n88312, n88313, n88314, n88315,
         n88316, n88317, n88318, n88319, n88320, n88321, n88322, n88323,
         n88324, n88325, n88326, n88327, n88328, n88329, n88330, n88331,
         n88332, n88333, n88334, n88335, n88336, n88337, n88338, n88339,
         n88340, n88341, n88342, n88343, n88344, n88345, n88346, n88347,
         n88348, n88349, n88350, n88351, n88352, n88353, n88354, n88355,
         n88356, n88357, n88358, n88359, n88360, n88361, n88362, n88363,
         n88364, n88365, n88366, n88367, n88368, n88369, n88370, n88371,
         n88372, n88373, n88374, n88375, n88376, n88377, n88378, n88379,
         n88380, n88381, n88382, n88383, n88384, n88385, n88386, n88387,
         n88388, n88389, n88390, n88391, n88392, n88393, n88394, n88395,
         n88396, n88397, n88398, n88399, n88400, n88401, n88402, n88403,
         n88404, n88405, n88406, n88407, n88408, n88409, n88410, n88411,
         n88412, n88413, n88414, n88415, n88416, n88417, n88418, n88419,
         n88420, n88421, n88422, n88423, n88424, n88425, n88426, n88427,
         n88428, n88429, n88430, n88431, n88432, n88433, n88434, n88435,
         n88436, n88437, n88438, n88439, n88440, n88441, n88442, n88443,
         n88444, n88445, n88446, n88447, n88448, n88449, n88450, n88451,
         n88452, n88453, n88454, n88455, n88456, n88457, n88458, n88459,
         n88460, n88461, n88462, n88463, n88464, n88465, n88466, n88467,
         n88468, n88469, n88470, n88471, n88472, n88473, n88474, n88475,
         n88476, n88477, n88478, n88479, n88480, n88481, n88482, n88483,
         n88484, n88485, n88486, n88487, n88488, n88489, n88490, n88491,
         n88492, n88493, n88494, n88495, n88496, n88497, n88498, n88499,
         n88500, n88501, n88502, n88503, n88504, n88505, n88506, n88507,
         n88508, n88509, n88510, n88511, n88512, n88513, n88514, n88515,
         n88516, n88517, n88518, n88519, n88520, n88521, n88522, n88523,
         n88524, n88525, n88526, n88527, n88528, n88529, n88530, n88531,
         n88532, n88533, n88534, n88535, n88536, n88537, n88538, n88539,
         n88540, n88541, n88542, n88543, n88544, n88545, n88546, n88547,
         n88548, n88549, n88550, n88551, n88552, n88553, n88554, n88555,
         n88556, n88557, n88558, n88559, n88560, n88561, n88562, n88563,
         n88564, n88565, n88566, n88567, n88568, n88569, n88570, n88571,
         n88572, n88573, n88574, n88575, n88576, n88577, n88578, n88579,
         n88580, n88581, n88582, n88583, n88584, n88585, n88586, n88587,
         n88588, n88589, n88590, n88591, n88592, n88593, n88594, n88595,
         n88596, n88597, n88598, n88599, n88600, n88601, n88602, n88603,
         n88604, n88605, n88606, n88607, n88608, n88609, n88610, n88611,
         n88612, n88613, n88614, n88615, n88616, n88617, n88618, n88619,
         n88620, n88621, n88622, n88623, n88624, n88625, n88626, n88627,
         n88628, n88629, n88630, n88631, n88632, n88633, n88634, n88635,
         n88636, n88637, n88638, n88639, n88640, n88641, n88642, n88643,
         n88644, n88645, n88646, n88647, n88648, n88649, n88650, n88651,
         n88652, n88653, n88654, n88655, n88656, n88657, n88658, n88659,
         n88660, n88661, n88662, n88663, n88664, n88665, n88666, n88667,
         n88668, n88669, n88670, n88671, n88672, n88673, n88674, n88675,
         n88676, n88677, n88678, n88679, n88680, n88681, n88682, n88683,
         n88684, n88685, n88686, n88687, n88688, n88689, n88690, n88691,
         n88692, n88693, n88694, n88695, n88696, n88697, n88698, n88699,
         n88700, n88701, n88702, n88703, n88704, n88705, n88706, n88707,
         n88708, n88709, n88710, n88711, n88712, n88713, n88714, n88715,
         n88716, n88717, n88718, n88719, n88720, n88721, n88722, n88723,
         n88724, n88725, n88726, n88727, n88728, n88729, n88730, n88731,
         n88732, n88733, n88734, n88735, n88736, n88737, n88738, n88739,
         n88740, n88741, n88742, n88743, n88744, n88745, n88746, n88747,
         n88748, n88749, n88750, n88751, n88752, n88753, n88754, n88755,
         n88756, n88757, n88758, n88759, n88760, n88761, n88762, n88763,
         n88764, n88765, n88766, n88767, n88768, n88769, n88770, n88771,
         n88772, n88773, n88774, n88775, n88776, n88777, n88778, n88779,
         n88780, n88781, n88782, n88783, n88784, n88785, n88786, n88787,
         n88788, n88789, n88790, n88791, n88792, n88793, n88794, n88795,
         n88796, n88797, n88798, n88799, n88800, n88801, n88802, n88803,
         n88804, n88805, n88806, n88807, n88808, n88809, n88810, n88811,
         n88812, n88813, n88814, n88815, n88816, n88817, n88818, n88819,
         n88820, n88821, n88822, n88823, n88824, n88825, n88826, n88827,
         n88828, n88829, n88830, n88831, n88832, n88833, n88834, n88835,
         n88836, n88837, n88838, n88839, n88840, n88841, n88842, n88843,
         n88844, n88845, n88846, n88847, n88848, n88849, n88850, n88851,
         n88852, n88853, n88854, n88855, n88856, n88857, n88858, n88859,
         n88860, n88861, n88862, n88863, n88864, n88865, n88866, n88867,
         n88868, n88869, n88870, n88871, n88872, n88873, n88874, n88875,
         n88876, n88877, n88878, n88879, n88880, n88881, n88882, n88883,
         n88884, n88885, n88886, n88887, n88888, n88889, n88890, n88891,
         n88892, n88893, n88894, n88895, n88896, n88897, n88898, n88899,
         n88900, n88901, n88902, n88903, n88904, n88905, n88906, n88907,
         n88908, n88909, n88910, n88911, n88912, n88913, n88914, n88915,
         n88916, n88917, n88918, n88919, n88920, n88921, n88922, n88923,
         n88924, n88925, n88926, n88927, n88928, n88929, n88930, n88931,
         n88932, n88933, n88934, n88935, n88936, n88937, n88938, n88939,
         n88940, n88941, n88942, n88943, n88944, n88945, n88946, n88947,
         n88948, n88949, n88950, n88951, n88952, n88953, n88954, n88955,
         n88956, n88957, n88958, n88959, n88960, n88961, n88962, n88963,
         n88964, n88965, n88966, n88967, n88968, n88969, n88970, n88971,
         n88972, n88973, n88974, n88975, n88976, n88977, n88978, n88979,
         n88980, n88981, n88982, n88983, n88984, n88985, n88986, n88987,
         n88988, n88989, n88990, n88991, n88992, n88993, n88994, n88995,
         n88996, n88997, n88998, n88999, n89000, n89001, n89002, n89003,
         n89004, n89005, n89006, n89007, n89008, n89009, n89010, n89011,
         n89012, n89013, n89014, n89015, n89016, n89017, n89018, n89019,
         n89020, n89021, n89022, n89023, n89024, n89025, n89026, n89027,
         n89028, n89029, n89030, n89031, n89032, n89033, n89034, n89035,
         n89036, n89037, n89038, n89039, n89040, n89041, n89042, n89043,
         n89044, n89045, n89046, n89047, n89048, n89049, n89050, n89051,
         n89052, n89053, n89054, n89055, n89056, n89057, n89058, n89059,
         n89060, n89061, n89062, n89063, n89064, n89065, n89066, n89067,
         n89068, n89069, n89070, n89071, n89072, n89073, n89074, n89075,
         n89076, n89077, n89078, n89079, n89080, n89081, n89082, n89083,
         n89084, n89085, n89086, n89087, n89088, n89089, n89090, n89091,
         n89092, n89093, n89094, n89095, n89096, n89097, n89098, n89099,
         n89100, n89101, n89102, n89103, n89104, n89105, n89106, n89107,
         n89108, n89109, n89110, n89111, n89112, n89113, n89114, n89115,
         n89116, n89117, n89118, n89119, n89120, n89121, n89122, n89123,
         n89124, n89125, n89126, n89127, n89128, n89129, n89130, n89131,
         n89132, n89133, n89134, n89135, n89136, n89137, n89138, n89139,
         n89140, n89141, n89142, n89143, n89144, n89145, n89146, n89147,
         n89148, n89149, n89150, n89151, n89152, n89153, n89154, n89155,
         n89156, n89157, n89158, n89159, n89160, n89161, n89162, n89163,
         n89164, n89165, n89166, n89167, n89168, n89169, n89170, n89171,
         n89172, n89173, n89174, n89175, n89176, n89177, n89178, n89179,
         n89180, n89181, n89182, n89183, n89184, n89185, n89186, n89187,
         n89188, n89189, n89190, n89191, n89192, n89193, n89194, n89195,
         n89196, n89197, n89198, n89199, n89200, n89201, n89202, n89203,
         n89204, n89205, n89206, n89207, n89208, n89209, n89210, n89211,
         n89212, n89213, n89214, n89215, n89216, n89217, n89218, n89219,
         n89220, n89221, n89222, n89223, n89224, n89225, n89226, n89227,
         n89228, n89229, n89230, n89231, n89232, n89233, n89234, n89235,
         n89236, n89237, n89238, n89239, n89240, n89241, n89242, n89243,
         n89244, n89245, n89246, n89247, n89248, n89249, n89250, n89251,
         n89252, n89253, n89254, n89255, n89256, n89257, n89258, n89259,
         n89260, n89261, n89262, n89263, n89264, n89265, n89266, n89267,
         n89268, n89269, n89270, n89271, n89272, n89273, n89274, n89275,
         n89276, n89277, n89278, n89279, n89280, n89281, n89282, n89283,
         n89284, n89285, n89286, n89287, n89288, n89289, n89290, n89291,
         n89292, n89293, n89294, n89295, n89296, n89297, n89298, n89299,
         n89300, n89301, n89302, n89303, n89304, n89305, n89306, n89307,
         n89308, n89309, n89310, n89311, n89312, n89313, n89314, n89315,
         n89316, n89317, n89318, n89319, n89320, n89321, n89322, n89323,
         n89324, n89325, n89326, n89327, n89328, n89329, n89330, n89331,
         n89332, n89333, n89334, n89335, n89336, n89337, n89338, n89339,
         n89340, n89341, n89342, n89343, n89344, n89345, n89346, n89347,
         n89348, n89349, n89350, n89351, n89352, n89353, n89354, n89355,
         n89356, n89357, n89358, n89359, n89360, n89361, n89362, n89363,
         n89364, n89365, n89366, n89367, n89368, n89369, n89370, n89371,
         n89372, n89373, n89374, n89375, n89376, n89377, n89378, n89379,
         n89380, n89381, n89382, n89383, n89384, n89385, n89386, n89387,
         n89388, n89389, n89390, n89391, n89392, n89393, n89394, n89395,
         n89396, n89397, n89398, n89399, n89400, n89401, n89402, n89403,
         n89404, n89405, n89406, n89407, n89408, n89409, n89410, n89411,
         n89412, n89413, n89414, n89415, n89416, n89417, n89418, n89419,
         n89420, n89421, n89422, n89423, n89424, n89425, n89426, n89427,
         n89428, n89429, n89430, n89431, n89432, n89433, n89434, n89435,
         n89436, n89437, n89438, n89439, n89440, n89441, n89442, n89443,
         n89444, n89445, n89446, n89447, n89448, n89449, n89450, n89451,
         n89452, n89453, n89454, n89455, n89456, n89457, n89458, n89459,
         n89460, n89461, n89462, n89463, n89464, n89465, n89466, n89467,
         n89468, n89469, n89470, n89471, n89472, n89473, n89474, n89475,
         n89476, n89477, n89478, n89479, n89480, n89481, n89482, n89483,
         n89484, n89485, n89486, n89487, n89488, n89489, n89490, n89491,
         n89492, n89493, n89494, n89495, n89496, n89497, n89498, n89499,
         n89500, n89501, n89502, n89503, n89504, n89505, n89506, n89507,
         n89508, n89509, n89510, n89511, n89512, n89513, n89514, n89515,
         n89516, n89517, n89518, n89519, n89520, n89521, n89522, n89523,
         n89524, n89525, n89526, n89527, n89528, n89529, n89530, n89531,
         n89532, n89533, n89534, n89535, n89536, n89537, n89538, n89539,
         n89540, n89541, n89542, n89543, n89544, n89545, n89546, n89547,
         n89548, n89549, n89550, n89551, n89552, n89553, n89554, n89555,
         n89556, n89557, n89558, n89559, n89560, n89561, n89562, n89563,
         n89564, n89565, n89566, n89567, n89568, n89569, n89570, n89571,
         n89572, n89573, n89574, n89575, n89576, n89577, n89578, n89579,
         n89580, n89581, n89582, n89583, n89584, n89585, n89586, n89587,
         n89588, n89589, n89590, n89591, n89592, n89593, n89594, n89595,
         n89596, n89597, n89598, n89599, n89600, n89601, n89602, n89603,
         n89604, n89605, n89606, n89607, n89608, n89609, n89610, n89611,
         n89612, n89613, n89614, n89615, n89616, n89617, n89618, n89619,
         n89620, n89621, n89622, n89623, n89624, n89625, n89626, n89627,
         n89628, n89629, n89630, n89631, n89632, n89633, n89634, n89635,
         n89636, n89637, n89638, n89639, n89640, n89641, n89642, n89643,
         n89644, n89645, n89646, n89647, n89648, n89649, n89650, n89651,
         n89652, n89653, n89654, n89655, n89656, n89657, n89658, n89659,
         n89660, n89661, n89662, n89663, n89664, n89665, n89666, n89667,
         n89668, n89669, n89670, n89671, n89672, n89673, n89674, n89675,
         n89676, n89677, n89678, n89679, n89680, n89681, n89682, n89683,
         n89684, n89685, n89686, n89687, n89688, n89689, n89690, n89691,
         n89692, n89693, n89694, n89695, n89696, n89697, n89698, n89699,
         n89700, n89701, n89702, n89703, n89704, n89705, n89706, n89707,
         n89708, n89709, n89710, n89711, n89712, n89713, n89714, n89715,
         n89716, n89717, n89718, n89719, n89720, n89721, n89722, n89723,
         n89724, n89725, n89726, n89727, n89728, n89729, n89730, n89731,
         n89732, n89733, n89734, n89735, n89736, n89737, n89738, n89739,
         n89740, n89741, n89742, n89743, n89744, n89745, n89746, n89747,
         n89748, n89749, n89750, n89751, n89752, n89753, n89754, n89755,
         n89756, n89757, n89758, n89759, n89760, n89761, n89762, n89763,
         n89764, n89765, n89766, n89767, n89768, n89769, n89770, n89771,
         n89772, n89773, n89774, n89775, n89776, n89777, n89778, n89779,
         n89780, n89781, n89782, n89783, n89784, n89785, n89786, n89787,
         n89788, n89789, n89790, n89791, n89792, n89793, n89794, n89795,
         n89796, n89797, n89798, n89799, n89800, n89801, n89802, n89803,
         n89804, n89805, n89806, n89807, n89808, n89809, n89810, n89811,
         n89812, n89813, n89814, n89815, n89816, n89817, n89818, n89819,
         n89820, n89821, n89822, n89823, n89824, n89825, n89826, n89827,
         n89828, n89829, n89830, n89831, n89832, n89833, n89834, n89835,
         n89836, n89837, n89838, n89839, n89840, n89841, n89842, n89843,
         n89844, n89845, n89846, n89847, n89848, n89849, n89850, n89851,
         n89852, n89853, n89854, n89855, n89856, n89857, n89858, n89859,
         n89860, n89861, n89862, n89863, n89864, n89865, n89866, n89867,
         n89868, n89869, n89870, n89871, n89872, n89873, n89874, n89875,
         n89876, n89877, n89878, n89879, n89880, n89881, n89882, n89883,
         n89884, n89885, n89886, n89887, n89888, n89889, n89890, n89891,
         n89892, n89893, n89894, n89895, n89896, n89897, n89898, n89899,
         n89900, n89901, n89902, n89903, n89904, n89905, n89906, n89907,
         n89908, n89909, n89910, n89911, n89912, n89913, n89914, n89915,
         n89916, n89917, n89918, n89919, n89920, n89921, n89922, n89923,
         n89924, n89925, n89926, n89927, n89928, n89929, n89930, n89931,
         n89932, n89933, n89934, n89935, n89936, n89937, n89938, n89939,
         n89940, n89941, n89942, n89943, n89944, n89945, n89946, n89947,
         n89948, n89949, n89950, n89951, n89952, n89953, n89954, n89955,
         n89956, n89957, n89958, n89959, n89960, n89961, n89962, n89963,
         n89964, n89965, n89966, n89967, n89968, n89969, n89970, n89971,
         n89972, n89973, n89974, n89975, n89976, n89977, n89978, n89979,
         n89980, n89981, n89982, n89983, n89984, n89985, n89986, n89987,
         n89988, n89989, n89990, n89991, n89992, n89993, n89994, n89995,
         n89996, n89997, n89998, n89999, n90000, n90001, n90002, n90003,
         n90004, n90005, n90006, n90007, n90008, n90009, n90010, n90011,
         n90012, n90013, n90014, n90015, n90016, n90017, n90018, n90019,
         n90020, n90021, n90022, n90023, n90024, n90025, n90026, n90027,
         n90028, n90029, n90030, n90031, n90032, n90033, n90034, n90035,
         n90036, n90037, n90038, n90039, n90040, n90041, n90042, n90043,
         n90044, n90045, n90046, n90047, n90048, n90049, n90050, n90051,
         n90052, n90053, n90054, n90055, n90056, n90057, n90058, n90059,
         n90060, n90061, n90062, n90063, n90064, n90065, n90066, n90067,
         n90068, n90069, n90070, n90071, n90072, n90073, n90074, n90075,
         n90076, n90077, n90078, n90079, n90080, n90081, n90082, n90083,
         n90084, n90085, n90086, n90087, n90088, n90089, n90090, n90091,
         n90092, n90093, n90094, n90095, n90096, n90097, n90098, n90099,
         n90100, n90101, n90102, n90103, n90104, n90105, n90106, n90107,
         n90108, n90109, n90110, n90111, n90112, n90113, n90114, n90115,
         n90116, n90117, n90118, n90119, n90120, n90121, n90122, n90123,
         n90124, n90125, n90126, n90127, n90128, n90129, n90130, n90131,
         n90132, n90133, n90134, n90135, n90136, n90137, n90138, n90139,
         n90140, n90141, n90142, n90143, n90144, n90145, n90146, n90147,
         n90148, n90149, n90150, n90151, n90152, n90153, n90154, n90155,
         n90156, n90157, n90158, n90159, n90160, n90161, n90162, n90163,
         n90164, n90165, n90166, n90167, n90168, n90169, n90170, n90171,
         n90172, n90173, n90174, n90175, n90176, n90177, n90178, n90179,
         n90180, n90181, n90182, n90183, n90184, n90185, n90186, n90187,
         n90188, n90189, n90190, n90191, n90192, n90193, n90194, n90195,
         n90196, n90197, n90198, n90199, n90200, n90201, n90202, n90203,
         n90204, n90205, n90206, n90207, n90208, n90209, n90210, n90211,
         n90212, n90213, n90214, n90215, n90216, n90217, n90218, n90219,
         n90220, n90221, n90222, n90223, n90224, n90225, n90226, n90227,
         n90228, n90229, n90230, n90231, n90232, n90233, n90234, n90235,
         n90236, n90237, n90238, n90239, n90240, n90241, n90242, n90243,
         n90244, n90245, n90246, n90247, n90248, n90249, n90250, n90251,
         n90252, n90253, n90254, n90255, n90256, n90257, n90258, n90259,
         n90260, n90261, n90262, n90263, n90264, n90265, n90266, n90267,
         n90268, n90269, n90270, n90271, n90272, n90273, n90274, n90275,
         n90276, n90277, n90278, n90279, n90280, n90282, n90283, n90284,
         n90285, n90286, n90290, n90291, n90292, n90293, n90294, n90295,
         n90296, n90297, n90298, n90299, n90300, n90301, n90302, n90303,
         n90304, n90305, n90306, n90307, n90308, n90309, n90310, n90311,
         n90312, n90313, n90314, n90315, n90316, n90317, n90318, n90319,
         n90320, n90321, n90322, n90323, n90324, n90325, n90326, n90327,
         n90328, n90329, n90330, n90331, n90332, n90333, n90334, n90335,
         n90336, n90337, n90338, n90339, n90340, n90341, n90342, n90343,
         n90344, n90345, n90346, n90347, n90348, n90349, n90350, n90351,
         n90352, n90353, n90354, n90355, n90356, n90357, n90358, n90359,
         n90360, n90361, n90362, n90363, n90364, n90365, n90366, n90367,
         n90368, n90369, n90370, n90371, n90372, n90373, n90374, n90375,
         n90376, n90377, n90378, n90379, n90380, n90381, n90382, n90383,
         n90384, n90385, n90386, n90387, n90388, n90389, n90390, n90391,
         n90392, n90393, n90394, n90395, n90396, n90397, n90398, n90399,
         n90400, n90401, n90402, n90403, n90404, n90405, n90406, n90407,
         n90408, n90409, n90410, n90411, n90412, n90413, n90414, n90415,
         n90416, n90417, n90418, n90419, n90420, n90421, n90422, n90423,
         n90424, n90425, n90426, n90427, n90428, n90429, n90430, n90431,
         n90432, n90433, n90434, n90435, n90436, n90437, n90438, n90439,
         n90440, n90441, n90442, n90443, n90444, n90445, n90446, n90447,
         n90448, n90449, n90450, n90451, n90452, n90453, n90454, n90455,
         n90456, n90457, n90458, n90459, n90460, n90461, n90462, n90463,
         n90464, n90465, n90466, n90467, n90468, n90469, n90470, n90471,
         n90472, n90473, n90474, n90475, n90476, n90477, n90478, n90479,
         n90480, n90481, n90482, n90483, n90484, n90485, n90486, n90487,
         n90488, n90489, n90490, n90491, n90492, n90493, n90494, n90495,
         n90496, n90497, n90498, n90499, n90500, n90501, n90502, n90503,
         n90504, n90505, n90506, n90507, n90508, n90509, n90510, n90511,
         n90512, n90513, n90514, n90515, n90516, n90517, n90518, n90519,
         n90520, n90521, n90522, n90523, n90524, n90525, n90526, n90527,
         n90528, n90529, n90530, n90531, n90532, n90533, n90534, n90535,
         n90536, n90537, n90538, n90539, n90540, n90541, n90542, n90543,
         n90544, n90545, n90546, n90547, n90548, n90549, n90550, n90551,
         n90552, n90553, n90554, n90555, n90556, n90557, n90558, n90559,
         n90560, n90561, n90562, n90563, n90564, n90565, n90566, n90567,
         n90568, n90569, n90570, n90571, n90572, n90573, n90574, n90575,
         n90576, n90577, n90578, n90579, n90580, n90581, n90582, n90583,
         n90584, n90585, n90586, n90587, n90588, n90589, n90590, n90591,
         n90592, n90593, n90594, n90595, n90596, n90597, n90598, n90599,
         n90600, n90601, n90602, n90603, n90604, n90605, n90606, n90607,
         n90608, n90609, n90610, n90611, n90612, n90613, n90614, n90615,
         n90616, n90617, n90618, n90619, n90620, n90621, n90622, n90623,
         n90624, n90625, n90626, n90627, n90628, n90629, n90630, n90631,
         n90632, n90633, n90634, n90635, n90636, n90637, n90638, n90639,
         n90640, n90641, n90642, n90643, n90644, n90645, n90646, n90647,
         n90648, n90649, n90650, n90651, n90652, n90653, n90654, n90655,
         n90656, n90657, n90658, n90659, n90660, n90661, n90662, n90663,
         n90664, n90665, n90666, n90667, n90668, n90669, n90670, n90671,
         n90672, n90673, n90674, n90675, n90676, n90677, n90678, n90679,
         n90680, n90681, n90682, n90683, n90684, n90685, n90686, n90687,
         n90688, n90689, n90690, n90691, n90692, n90693, n90694, n90695,
         n90696, n90697, n90698, n90699, n90700, n90701, n90702, n90703,
         n90704, n90705, n90706, n90707, n90708, n90709, n90710, n90711,
         n90712, n90713, n90714, n90715, n90716, n90717, n90718, n90719,
         n90720, n90721, n90722, n90723, n90724, n90725, n90726, n90727,
         n90728, n90729, n90730, n90731, n90732, n90733, n90734, n90735,
         n90736, n90737, n90738, n90739, n90740, n90741, n90742, n90743,
         n90744, n90745, n90746, n90747, n90748, n90749, n90750, n90751,
         n90752, n90753, n90754, n90755, n90756, n90757, n90758, n90759,
         n90760, n90761, n90762, n90763, n90764, n90765, n90766, n90767,
         n90768, n90769, n90770, n90771, n90772, n90773, n90774, n90775,
         n90776, n90777, n90778, n90779, n90780, n90781, n90782, n90783,
         n90784, n90785, n90786, n90787, n90788, n90789, n90790, n90791,
         n90792, n90793, n90794, n90795, n90796, n90797, n90798, n90799,
         n90800, n90801, n90802, n90803, n90804, n90805, n90806, n90807,
         n90808, n90809, n90810, n90811, n90812, n90813, n90814, n90815,
         n90816, n90817, n90818, n90819, n90820, n90821, n90822, n90823,
         n90824, n90825, n90826, n90827, n90828, n90829, n90830, n90831,
         n90832, n90833, n90834, n90835, n90836, n90837, n90838, n90839,
         n90840, n90841, n90842, n90843, n90844, n90845, n90846, n90847,
         n90848, n90849, n90850, n90851, n90852, n90853, n90854, n90855,
         n90856, n90857, n90858, n90859, n90860, n90861, n90862, n90863,
         n90864, n90865, n90866, n90867, n90868, n90869, n90870, n90871,
         n90872, n90873, n90874, n90875, n90876, n90877, n90878, n90879,
         n90880, n90881, n90882, n90883, n90884, n90885, n90886, n90887,
         n90888, n90889, n90890, n90891, n90892, n90893, n90894, n90895,
         n90896, n90897, n90898, n90899, n90900, n90901, n90902, n90903,
         n90904, n90905, n90906, n90907, n90908, n90909, n90910, n90911,
         n90912, n90913, n90914, n90915, n90916, n90917, n90918, n90919,
         n90920, n90921, n90922, n90923, n90924, n90925, n90926, n90927,
         n90928, n90929, n90930, n90931, n90932, n90933, n90934, n90935,
         n90936, n90937, n90938, n90939, n90940, n90941, n90942, n90943,
         n90944, n90945, n90946, n90947, n90948, n90949, n90950, n90951,
         n90952, n90953, n90954, n90955, n90956, n90957, n90958, n90959,
         n90960, n90961, n90962, n90963, n90964, n90965, n90966, n90967,
         n90968, n90969, n90970, n90971, n90972, n90973, n90974, n90975,
         n90976, n90977, n90978, n90979, n90980, n90981, n90982, n90983,
         n90984, n90985, n90986, n90987, n90988, n90989, n90990, n90991,
         n90992, n90993, n90994, n90995, n90996, n90997, n90998, n90999,
         n91000, n91001, n91002, n91003, n91004, n91005, n91006, n91007,
         n91008, n91009, n91010, n91011, n91012, n91013, n91014, n91015,
         n91016, n91017, n91018, n91019, n91020, n91021, n91022, n91023,
         n91024, n91025, n91026, n91027, n91028, n91029, n91030, n91031,
         n91032, n91033, n91034, n91035, n91036, n91037, n91038, n91039,
         n91040, n91041, n91042, n91043, n91044, n91045, n91046, n91047,
         n91048, n91049, n91050, n91051, n91052, n91053, n91054, n91055,
         n91056, n91057, n91058, n91059, n91060, n91061, n91062, n91063,
         n91064, n91065, n91066, n91067, n91068, n91069, n91070, n91071,
         n91072, n91073, n91074, n91075, n91076, n91077, n91078, n91079,
         n91080, n91081, n91082, n91083, n91084, n91085, n91086, n91087,
         n91088, n91089, n91090, n91091, n91092, n91093, n91094, n91095,
         n91096, n91097, n91098, n91099, n91100, n91101, n91102, n91103,
         n91104, n91105, n91106, n91107, n91108, n91109, n91110, n91111,
         n91112, n91113, n91114, n91115, n91116, n91117, n91118, n91119,
         n91120, n91121, n91122, n91123, n91124, n91125, n91126, n91127,
         n91128, n91129, n91130, n91131, n91132, n91133, n91134, n91135,
         n91136, n91137, n91138, n91139, n91140, n91141, n91142, n91143,
         n91144, n91145, n91146, n91147, n91148, n91149, n91150, n91151,
         n91152, n91153, n91154, n91155, n91156, n91157, n91158, n91159,
         n91160, n91161, n91162, n91163, n91164, n91165, n91166, n91167,
         n91168, n91169, n91170, n91171, n91172, n91173, n91174, n91175,
         n91176, n91177, n91178, n91179, n91180, n91181, n91182, n91183,
         n91184, n91185, n91186, n91187, n91188, n91189, n91190, n91191,
         n91192, n91193, n91194, n91195, n91196, n91197, n91198, n91199,
         n91200, n91201, n91202, n91203, n91204, n91205, n91206, n91207,
         n91208, n91209, n91210, n91211, n91212, n91213, n91214, n91215,
         n91216, n91217, n91218, n91219, n91220, n91221, n91222, n91223,
         n91224, n91225, n91226, n91227, n91228, n91229, n91230, n91231,
         n91232, n91233, n91234, n91235, n91236, n91237, n91238, n91239,
         n91240, n91241, n91242, n91243, n91244, n91245, n91246, n91247,
         n91248, n91249, n91250, n91251, n91252, n91253, n91254, n91255,
         n91256, n91257, n91258, n91259, n91260, n91261, n91262, n91263,
         n91264, n91265, n91266, n91267, n91268, n91269, n91270, n91271,
         n91272, n91273, n91274, n91275, n91276, n91277, n91278, n91279,
         n91280, n91281, n91282, n91283, n91284, n91285, n91286, n91287,
         n91288, n91289, n91290, n91291, n91292, n91293, n91294, n91295,
         n91296, n91297, n91298, n91299, n91300, n91301, n91302, n91303,
         n91304, n91305, n91306, n91307, n91308, n91309, n91310, n91311,
         n91312, n91313, n91314, n91315, n91316, n91317, n91318, n91319,
         n91320, n91321, n91322, n91323, n91324, n91325, n91326, n91327,
         n91328, n91329, n91330, n91331, n91332, n91333, n91334, n91335,
         n91336, n91337, n91338, n91339, n91340, n91341, n91342, n91343,
         n91344, n91345, n91346, n91347, n91348, n91349, n91350, n91351,
         n91352, n91353, n91354, n91355, n91356, n91357, n91358, n91359,
         n91360, n91361, n91362, n91363, n91364, n91365, n91366, n91367,
         n91368, n91369, n91370, n91371, n91372, n91373, n91374, n91375,
         n91376, n91377, n91378, n91379, n91380, n91381, n91382, n91383,
         n91384, n91385, n91386, n91387, n91388, n91389, n91390, n91391,
         n91392, n91393, n91394, n91395, n91396, n91397, n91398, n91399,
         n91400, n91401, n91402, n91403, n91404, n91405, n91406, n91407,
         n91408, n91409, n91410, n91411, n91412, n91413, n91414, n91415,
         n91416, n91417, n91418, n91419, n91420, n91421, n91422, n91423,
         n91424, n91425, n91426, n91427, n91428, n91429, n91430, n91431,
         n91432, n91433, n91434, n91435, n91436, n91437, n91438, n91439,
         n91440, n91441, n91442, n91443, n91444, n91445, n91446, n91447,
         n91448, n91449, n91450, n91451, n91452, n91453, n91454, n91455,
         n91456, n91457, n91458, n91459, n91460, n91461, n91462, n91463,
         n91464, n91465, n91466, n91467, n91468, n91469, n91470, n91471,
         n91472, n91473, n91474, n91475, n91476, n91477, n91478, n91479,
         n91480, n91481, n91482, n91483, n91484, n91485, n91486, n91487,
         n91488, n91489, n91490, n91491, n91492, n91493, n91494, n91495,
         n91496, n91497, n91498, n91499, n91500, n91501, n91502, n91503,
         n91504, n91505, n91506, n91507, n91508, n91509, n91510, n91511,
         n91512, n91513, n91514, n91515, n91516, n91517, n91518, n91519,
         n91520, n91521, n91522, n91523, n91524, n91525, n91526, n91527,
         n91528, n91529, n91530, n91531, n91532, n91533, n91534, n91535,
         n91536, n91537, n91538, n91539, n91540, n91541, n91542, n91543,
         n91544, n91545, n91546, n91547, n91548, n91549, n91550, n91551,
         n91552, n91553, n91554, n91555, n91556, n91557, n91558, n91559,
         n91560, n91561, n91562, n91563, n91564, n91565, n91566, n91567,
         n91568, n91569, n91570, n91571, n91572, n91573, n91574, n91575,
         n91576, n91577, n91578, n91579, n91580, n91581, n91582, n91583,
         n91584, n91585, n91586, n91587, n91588, n91589, n91590, n91591,
         n91592, n91593, n91594, n91595, n91596, n91597, n91598, n91599,
         n91600, n91601, n91602, n91603, n91604, n91605, n91606, n91607,
         n91608, n91609, n91610, n91611, n91612, n91613, n91614, n91615,
         n91616, n91617, n91618, n91619, n91620, n91621, n91622, n91623,
         n91624, n91625, n91626, n91627, n91628, n91629, n91630, n91631,
         n91632, n91633, n91634, n91635, n91636, n91637, n91638, n91639,
         n91640, n91641, n91642, n91643, n91644, n91645, n91646, n91647,
         n91648, n91649, n91650, n91651, n91652, n91653, n91654, n91655,
         n91656, n91657, n91658, n91659, n91660, n91661, n91662, n91663,
         n91664, n91665, n91666, n91667, n91668, n91669, n91670, n91671,
         n91672, n91673, n91674, n91675, n91676, n91677, n91678, n91679,
         n91680, n91681, n91682, n91683, n91684, n91685, n91686, n91687,
         n91688, n91689, n91690, n91691, n91692, n91693, n91694, n91695,
         n91696, n91697, n91698, n91699, n91700, n91701, n91702, n91703,
         n91704, n91705, n91706, n91707, n91708, n91709, n91710, n91711,
         n91712, n91713, n91714, n91715, n91716, n91717, n91718, n91719,
         n91720, n91721, n91722, n91723, n91724, n91725, n91726, n91727,
         n91728, n91729, n91730, n91731, n91732, n91733, n91734, n91735,
         n91736, n91737, n91738, n91739, n91740, n91741, n91742, n91743,
         n91744, n91745, n91746, n91747, n91748, n91749, n91750, n91751,
         n91752, n91753, n91754, n91755, n91756, n91757, n91758, n91759,
         n91760, n91761, n91762, n91763, n91764, n91765, n91766, n91767,
         n91768, n91769, n91770, n91771, n91772, n91773, n91774, n91775,
         n91776, n91777, n91778, n91779, n91780, n91781, n91782, n91783,
         n91784, n91785, n91786, n91787, n91788, n91789, n91790, n91791,
         n91792, n91793, n91794, n91795, n91796, n91797, n91798, n91799,
         n91800, n91801, n91802, n91803, n91804, n91805, n91806, n91807,
         n91808, n91809, n91810, n91811, n91812, n91813, n91814, n91815,
         n91816, n91817, n91818, n91819, n91820, n91821, n91822, n91823,
         n91824, n91825, n91826, n91827, n91828, n91829, n91830, n91831,
         n91832, n91833, n91834, n91835, n91836, n91837, n91838, n91839,
         n91840, n91841, n91842, n91843, n91844, n91845, n91846, n91847,
         n91848, n91849, n91850, n91851, n91852, n91853, n91854, n91855,
         n91856, n91857, n91858, n91859, n91860, n91861, n91862, n91863,
         n91864, n91865, n91866, n91867, n91868, n91869, n91870, n91871,
         n91872, n91873, n91874, n91875, n91876, n91877, n91878, n91879,
         n91880, n91881, n91882, n91883, n91884, n91885, n91886, n91887,
         n91888, n91889, n91890, n91891, n91892, n91893, n91894, n91895,
         n91896, n91897, n91898, n91899, n91900, n91901, n91902, n91903,
         n91904, n91905, n91906, n91907, n91908, n91909, n91910, n91911,
         n91912, n91913, n91914, n91915, n91916, n91917, n91918, n91919,
         n91920, n91921, n91922, n91923, n91924, n91925, n91926, n91927,
         n91928, n91929, n91930, n91931, n91932, n91933, n91934, n91935,
         n91936, n91937, n91938, n91939, n91940, n91941, n91942, n91943,
         n91944, n91945, n91946, n91947, n91948, n91949, n91950, n91951,
         n91952, n91953, n91954, n91955, n91956, n91957, n91958, n91959,
         n91960, n91961, n91962, n91963, n91964, n91965, n91966, n91967,
         n91968, n91969, n91970, n91971, n91972, n91973, n91974, n91975,
         n91976, n91977, n91978, n91979, n91980, n91981, n91982, n91983,
         n91984, n91985, n91986, n91987, n91988, n91989, n91990, n91991,
         n91992, n91993, n91994, n91995, n91996, n91997, n91998, n91999,
         n92000, n92001, n92002, n92003, n92004, n92005, n92006, n92007,
         n92008, n92009, n92010, n92011, n92012, n92013, n92014, n92015,
         n92016, n92017, n92018, n92019, n92020, n92021, n92022, n92023,
         n92024, n92025, n92026, n92027, n92028, n92029, n92030, n92031,
         n92032, n92033, n92034, n92035, n92036, n92037, n92038, n92039,
         n92040, n92041, n92042, n92043, n92044, n92045, n92046, n92047,
         n92048, n92049, n92050, n92051, n92052, n92053, n92054, n92055,
         n92056, n92057, n92058, n92059, n92060, n92061, n92062, n92063,
         n92064, n92065, n92066, n92067, n92068, n92069, n92070, n92071,
         n92072, n92073, n92074, n92075, n92076, n92077, n92078, n92079,
         n92080, n92081, n92082, n92083, n92084, n92085, n92086, n92087,
         n92088, n92089, n92090, n92091, n92092, n92093, n92094, n92095,
         n92096, n92097, n92098, n92099, n92100, n92101, n92102, n92103,
         n92104, n92105, n92106, n92107, n92108, n92109, n92110, n92111,
         n92112, n92113, n92114, n92115, n92116, n92117, n92118, n92119,
         n92120, n92121, n92122, n92123, n92124, n92125, n92126, n92127,
         n92128, n92129, n92130, n92131, n92132, n92133, n92134, n92135,
         n92136, n92137, n92138, n92139, n92140, n92141, n92142, n92143,
         n92144, n92145, n92146, n92147, n92148, n92149, n92150, n92151,
         n92152, n92153, n92154, n92155, n92156, n92157, n92158, n92159,
         n92160, n92161, n92162, n92163, n92164, n92165, n92166, n92167,
         n92168, n92169, n92170, n92171, n92172, n92173, n92174, n92175,
         n92176, n92177, n92178, n92179, n92180, n92181, n92182, n92183,
         n92184, n92185, n92186, n92187, n92188, n92189, n92190, n92191,
         n92192, n92193, n92194, n92195, n92196, n92197, n92198, n92199,
         n92200, n92201, n92202, n92203, n92204, n92205, n92206, n92207,
         n92208, n92209, n92210, n92211, n92212, n92213, n92214, n92215,
         n92216, n92217, n92218, n92219, n92220, n92221, n92222, n92223,
         n92224, n92225, n92226, n92227, n92228, n92229, n92230, n92231,
         n92232, n92233, n92234, n92235, n92236, n92237, n92238, n92239,
         n92240, n92241, n92242, n92243, n92244, n92245, n92246, n92247,
         n92248, n92249, n92250, n92251, n92252, n92253, n92254, n92255,
         n92256, n92257, n92258, n92259, n92260, n92261, n92262, n92263,
         n92264, n92265, n92266, n92267, n92268, n92269, n92270, n92271,
         n92272, n92273, n92274, n92275, n92276, n92277, n92278, n92279,
         n92280, n92281, n92282, n92283, n92284, n92285, n92286, n92287,
         n92288, n92289, n92290, n92291, n92292, n92293, n92294, n92295,
         n92296, n92297, n92298, n92299, n92300, n92301, n92302, n92303,
         n92304, n92305, n92306, n92307, n92308, n92309, n92310, n92311,
         n92312, n92313, n92314, n92315, n92316, n92317, n92318, n92319,
         n92320, n92321, n92322, n92323, n92324, n92325, n92326, n92327,
         n92328, n92329, n92330, n92331, n92332, n92333, n92334, n92335,
         n92336, n92337, n92338, n92339, n92340, n92341, n92342, n92343,
         n92344, n92345, n92346, n92347, n92348, n92349, n92350, n92351,
         n92352, n92353, n92354, n92355, n92356, n92357, n92358, n92359,
         n92360, n92361, n92362, n92363, n92364, n92365, n92366, n92367,
         n92368, n92369, n92370, n92371, n92372, n92373, n92374, n92375,
         n92376, n92377, n92378, n92379, n92380, n92381, n92382, n92383,
         n92384, n92385, n92386, n92387, n92388, n92389, n92390, n92391,
         n92392, n92393, n92394, n92395, n92396, n92397, n92398, n92399,
         n92400, n92401, n92402, n92403, n92404, n92405, n92406, n92407,
         n92408, n92409, n92410, n92411, n92412, n92413, n92414, n92415,
         n92416, n92417, n92418, n92419, n92420, n92421, n92422, n92423,
         n92424, n92425, n92426, n92427, n92428, n92429, n92430, n92431,
         n92432, n92433, n92434, n92435, n92436, n92437, n92438, n92439,
         n92440, n92441, n92442, n92443, n92444, n92445, n92446, n92447,
         n92448, n92449, n92450, n92451, n92452, n92453, n92454, n92455,
         n92456, n92457, n92458, n92459, n92460, n92461, n92462, n92463,
         n92464, n92465, n92466, n92467, n92468, n92469, n92470, n92471,
         n92472, n92473, n92474, n92475, n92476, n92477, n92478, n92479,
         n92480, n92481, n92482, n92483, n92484, n92485, n92486, n92487,
         n92488, n92489, n92490, n92491, n92492, n92493, n92494, n92495,
         n92496, n92497, n92498, n92499, n92500, n92501, n92502, n92503,
         n92504, n92505, n92506, n92507, n92508, n92509, n92510, n92511,
         n92512, n92513, n92514, n92515, n92516, n92517, n92518, n92519,
         n92520, n92521, n92522, n92523, n92524, n92525, n92526, n92527,
         n92528, n92529, n92530, n92531, n92532, n92533, n92534, n92535,
         n92536, n92537, n92538, n92539, n92540, n92541, n92542, n92543,
         n92544, n92545, n92546, n92547, n92548, n92549, n92550, n92551,
         n92552, n92553, n92554, n92555, n92556, n92557, n92558, n92559,
         n92560, n92561, n92562, n92563, n92564, n92565, n92566, n92567,
         n92568, n92569, n92570, n92571, n92572, n92573, n92574, n92575,
         n92576, n92577, n92578, n92579, n92580, n92581, n92582, n92583,
         n92584, n92585, n92586, n92587, n92588, n92589, n92590, n92591,
         n92592, n92593, n92594, n92595, n92596, n92597, n92598, n92599,
         n92600, n92601, n92602, n92603, n92604, n92605, n92606, n92607,
         n92608, n92609, n92610, n92611, n92612, n92613, n92614, n92615,
         n92616, n92617, n92618, n92619, n92620, n92621, n92622, n92623,
         n92624, n92625, n92626, n92627, n92628, n92629, n92630, n92631,
         n92632, n92633, n92634, n92635, n92636, n92637, n92638, n92639,
         n92640, n92641, n92642, n92643, n92644, n92645, n92646, n92647,
         n92648, n92649, n92650, n92651, n92652, n92653, n92654, n92655,
         n92656, n92657, n92658, n92659, n92660, n92661, n92662, n92663,
         n92664, n92665, n92666, n92667, n92668, n92669, n92670, n92671,
         n92672, n92673, n92674, n92675, n92676, n92677, n92678, n92679,
         n92680, n92681, n92682, n92683, n92684, n92685, n92686, n92687,
         n92688, n92689, n92690, n92691, n92692, n92693, n92694, n92695,
         n92696, n92697, n92698, n92699, n92700, n92701, n92702, n92703,
         n92704, n92705, n92706, n92707, n92708, n92709, n92710, n92711,
         n92712, n92713, n92714, n92715, n92716, n92717, n92718, n92719,
         n92720, n92721, n92722, n92723, n92724, n92725, n92726, n92727,
         n92728, n92729, n92730, n92731, n92732, n92733, n92734, n92735,
         n92736, n92737, n92738, n92739, n92740, n92741, n92742, n92743,
         n92744, n92745, n92746, n92747, n92748, n92749, n92750, n92751,
         n92752, n92753, n92754, n92755, n92756, n92757, n92758, n92759,
         n92760, n92761, n92762, n92763, n92764, n92765, n92766, n92767,
         n92768, n92769, n92770, n92771, n92772, n92773, n92774, n92775,
         n92776, n92777, n92778, n92779, n92780, n92781, n92782, n92783,
         n92784, n92785, n92786, n92787, n92788, n92789, n92790, n92791,
         n92792, n92793, n92794, n92795, n92796, n92797, n92798, n92799,
         n92800, n92801, n92802, n92803, n92804, n92805, n92806, n92807,
         n92808, n92809, n92810, n92811, n92812, n92813, n92814, n92815,
         n92816, n92817, n92818, n92819, n92820, n92821, n92822, n92823,
         n92824, n92825, n92826, n92827, n92828, n92829, n92830, n92831,
         n92832, n92833, n92834, n92835, n92836, n92837, n92838, n92839,
         n92840, n92841, n92842, n92843, n92844, n92845, n92846, n92847,
         n92848, n92849, n92850, n92851, n92852, n92853, n92854, n92855,
         n92856, n92857, n92858, n92859, n92860, n92861, n92862, n92863,
         n92864, n92865, n92866, n92867, n92868, n92869, n92870, n92871,
         n92872, n92873, n92874, n92875, n92876, n92877, n92878, n92879,
         n92880, n92881, n92882, n92883, n92884, n92885, n92886, n92887,
         n92888, n92889, n92890, n92891, n92892, n92893, n92894, n92895,
         n92896, n92897, n92898, n92899, n92900, n92901, n92902, n92903,
         n92904, n92905, n92906, n92907, n92908, n92909, n92910, n92911,
         n92912, n92913, n92914, n92915, n92916, n92917, n92918, n92919,
         n92920, n92921, n92922, n92923, n92924, n92925, n92926, n92927,
         n92928, n92929, n92930, n92931, n92932, n92933, n92934, n92935,
         n92936, n92937, n92938, n92939, n92940, n92941, n92942, n92943,
         n92944, n92945, n92946, n92947, n92948, n92949, n92950, n92951,
         n92952, n92953, n92954, n92955, n92956, n92957, n92958, n92959,
         n92960, n92961, n92962, n92963, n92964, n92965, n92966, n92967,
         n92968, n92969, n92970, n92971, n92972, n92973, n92974, n92975,
         n92976, n92977, n92978, n92979, n92980, n92981, n92982, n92983,
         n92984, n92985, n92986, n92987, n92988, n92989, n92990, n92991,
         n92992, n92993, n92994, n92995, n92996, n92997, n92998, n92999,
         n93000, n93001, n93002, n93003, n93004, n93005, n93006, n93007,
         n93008, n93009, n93010, n93011, n93012, n93013, n93014, n93015,
         n93016, n93017, n93018, n93019, n93020, n93021, n93022, n93023,
         n93024, n93025, n93026, n93027, n93028, n93029, n93030, n93031,
         n93032, n93033, n93034, n93035, n93036, n93037, n93038, n93039,
         n93040, n93041, n93042, n93043, n93044, n93045, n93046, n93047,
         n93048, n93049, n93050, n93051, n93052, n93053, n93054, n93055,
         n93056, n93057, n93058, n93059, n93060, n93061, n93062, n93063,
         n93064, n93065, n93066, n93067, n93068, n93069, n93070, n93071,
         n93072, n93073, n93074, n93075, n93076, n93077, n93078, n93079,
         n93080, n93081, n93082, n93083, n93084, n93085, n93086, n93087,
         n93088, n93089, n93090, n93091, n93092, n93093, n93094, n93095,
         n93096, n93097, n93098, n93099, n93100, n93101, n93102, n93103,
         n93104, n93105, n93106, n93107, n93108, n93109, n93110, n93111,
         n93112, n93113, n93114, n93115, n93116, n93117, n93118, n93119,
         n93120, n93121, n93122, n93123, n93124, n93125, n93126, n93127,
         n93128, n93129, n93130, n93131, n93132, n93133, n93134, n93135,
         n93136, n93137, n93138, n93139, n93140, n93141, n93142, n93143,
         n93144, n93145, n93146, n93147, n93148, n93149, n93150, n93151,
         n93152, n93153, n93154, n93155, n93156, n93157, n93158, n93159,
         n93160, n93161, n93162, n93163, n93164, n93165, n93166, n93167,
         n93168, n93169, n93170, n93171, n93172, n93173, n93174, n93175,
         n93176, n93177, n93178, n93179, n93180, n93181, n93182, n93183,
         n93184, n93185, n93186, n93187, n93188, n93189, n93190, n93191,
         n93192, n93193, n93194, n93195, n93196, n93197, n93198, n93199,
         n93200, n93201, n93202, n93203, n93204, n93205, n93206, n93207,
         n93208, n93209, n93210, n93211, n93212, n93213, n93214, n93215,
         n93216, n93217, n93218, n93219, n93220, n93221, n93222, n93223,
         n93224, n93225, n93226, n93227, n93228, n93229, n93230, n93231,
         n93232, n93233, n93234, n93235, n93236, n93237, n93238, n93239,
         n93240, n93241, n93242, n93243, n93244, n93245, n93246, n93247,
         n93248, n93249, n93250, n93251, n93252, n93253, n93254, n93255,
         n93256, n93257, n93258, n93259, n93260, n93261, n93262, n93263,
         n93264, n93265, n93266, n93267, n93268, n93269, n93270, n93271,
         n93272, n93273, n93274, n93275, n93276, n93277, n93278, n93279,
         n93280, n93281, n93282, n93283, n93284, n93285, n93286, n93287,
         n93288, n93289, n93290, n93291, n93292, n93293, n93294, n93295,
         n93296, n93297, n93298, n93299, n93300, n93301, n93302, n93303,
         n93304, n93305, n93306, n93307, n93308, n93309, n93310, n93311,
         n93312, n93313, n93314, n93315, n93316, n93317, n93318, n93319,
         n93320, n93321, n93322, n93323, n93324, n93325, n93326, n93327,
         n93328, n93329, n93330, n93331, n93332, n93333, n93334, n93335,
         n93336, n93337, n93338, n93339, n93340, n93341, n93342, n93343,
         n93344, n93345, n93346, n93347, n93348, n93349, n93350, n93351,
         n93352, n93353, n93354, n93355, n93356, n93357, n93358, n93359,
         n93360, n93361, n93362, n93363, n93364, n93365, n93366, n93367,
         n93368, n93369, n93370, n93371, n93372, n93373, n93374, n93375,
         n93376, n93377, n93378, n93379, n93380, n93381, n93382, n93383,
         n93384, n93385, n93386, n93387, n93388, n93389, n93390, n93391,
         n93392, n93393, n93394, n93395, n93396, n93397, n93398, n93399,
         n93400, n93401, n93402, n93403, n93404, n93405, n93406, n93407,
         n93408, n93409, n93410, n93411, n93412, n93413, n93414, n93415,
         n93416, n93417, n93418, n93419, n93420, n93421, n93422, n93423,
         n93424, n93425, n93426, n93427, n93428, n93429, n93430, n93431,
         n93432, n93433, n93434, n93435, n93436, n93437, n93438, n93439,
         n93440, n93441, n93442, n93443, n93444, n93445, n93446, n93447,
         n93448, n93449, n93450, n93451, n93452, n93453, n93454, n93455,
         n93456, n93457, n93458, n93459, n93460, n93461, n93462, n93463,
         n93464, n93465, n93466, n93467, n93468, n93469, n93470, n93471,
         n93472, n93473, n93474, n93475, n93476, n93477, n93478, n93479,
         n93480, n93481, n93482, n93483, n93484, n93485, n93486, n93487,
         n93488, n93489, n93490, n93491, n93492, n93493, n93494, n93495,
         n93496, n93497, n93498, n93499, n93500, n93501, n93502, n93503,
         n93504, n93505, n93506, n93507, n93508, n93509, n93510, n93511,
         n93512, n93513, n93514, n93515, n93516, n93517, n93518, n93519,
         n93520, n93521, n93522, n93523, n93524, n93525, n93526, n93527,
         n93528, n93529, n93530, n93531, n93532, n93533, n93534, n93535,
         n93536, n93537, n93538, n93539, n93540, n93541, n93542, n93543,
         n93544, n93545, n93546, n93547, n93548, n93549, n93550, n93551,
         n93552, n93553, n93554, n93555, n93556, n93557, n93558, n93559,
         n93560, n93561, n93562, n93563, n93564, n93565, n93566, n93567,
         n93568, n93569, n93570, n93571, n93572, n93573, n93574, n93575,
         n93576, n93577, n93578, n93579, n93580, n93581, n93582, n93583,
         n93584, n93585, n93586, n93587, n93588, n93589, n93590, n93591,
         n93592, n93593, n93594, n93595, n93596, n93597, n93598, n93599,
         n93600, n93601, n93602, n93603, n93604, n93605, n93606, n93607,
         n93608, n93609, n93610, n93611, n93612, n93613, n93614, n93615,
         n93616, n93617, n93618, n93619, n93620, n93621, n93622, n93623,
         n93624, n93625, n93626, n93627, n93628, n93629, n93630, n93631,
         n93632, n93633, n93634, n93635, n93636, n93637, n93638, n93639,
         n93640, n93641, n93642, n93643, n93644, n93645, n93646, n93647,
         n93648, n93649, n93650, n93651, n93652, n93653, n93654, n93655,
         n93656, n93657, n93658, n93659, n93660, n93661, n93662, n93663,
         n93664, n93665, n93666, n93667, n93668, n93669, n93670, n93671,
         n93672, n93673, n93674, n93675, n93676, n93677, n93678, n93679,
         n93680, n93681, n93682, n93683, n93684, n93685, n93686, n93687,
         n93688, n93689, n93690, n93691, n93692, n93693, n93694, n93695,
         n93696, n93697, n93698, n93699, n93700, n93701, n93702, n93703,
         n93704, n93705, n93706, n93707, n93708, n93709, n93710, n93711,
         n93712, n93713, n93714, n93715, n93716, n93717, n93718, n93719,
         n93720, n93721, n93722, n93723, n93724, n93725, n93726, n93727,
         n93728, n93729, n93730, n93731, n93732, n93733, n93734, n93735,
         n93736, n93737, n93738, n93739, n93740, n93741, n93742, n93743,
         n93744, n93745, n93746, n93747, n93748, n93749, n93750, n93751,
         n93752, n93753, n93754, n93755, n93756, n93757, n93758, n93759,
         n93760, n93761, n93762, n93763, n93764, n93765, n93766, n93767,
         n93768, n93769, n93770, n93771, n93772, n93773, n93774, n93775,
         n93776, n93777, n93778, n93779, n93780, n93781, n93782, n93783,
         n93784, n93785, n93786, n93787, n93788, n93789, n93790, n93791,
         n93792, n93793, n93794, n93795, n93796, n93797, n93798, n93799,
         n93800, n93801, n93802, n93803, n93804, n93805, n93806, n93807,
         n93808, n93809, n93810, n93811, n93812, n93813, n93814, n93815,
         n93816, n93817, n93818, n93819, n93820, n93821, n93822, n93823,
         n93824, n93825, n93826, n93827, n93828, n93829, n93830, n93831,
         n93832, n93833, n93834, n93835, n93836, n93837, n93838, n93839,
         n93840, n93841, n93842, n93843, n93844, n93845, n93846, n93847,
         n93848, n93849, n93850, n93851, n93852, n93853, n93854, n93855,
         n93856, n93857, n93858, n93859, n93860, n93861, n93862, n93863,
         n93864, n93865, n93866, n93867, n93868, n93869, n93870, n93871,
         n93872, n93873, n93874, n93875, n93876, n93877, n93878, n93879,
         n93880, n93881, n93882, n93883, n93884, n93885, n93886, n93887,
         n93888, n93889, n93890, n93891, n93892, n93893, n93894, n93895,
         n93896, n93897, n93898, n93899, n93900, n93901, n93902, n93903,
         n93904, n93905, n93906, n93907, n93908, n93909, n93910, n93911,
         n93912, n93913, n93914, n93915, n93916, n93917, n93918, n93919,
         n93920, n93921, n93922, n93923, n93924, n93925, n93926, n93927,
         n93928, n93929, n93930, n93931, n93932, n93933, n93934, n93935,
         n93936, n93937, n93938, n93939, n93940, n93941, n93942, n93943,
         n93944, n93945, n93946, n93947, n93948, n93949, n93950, n93951,
         n93952, n93953, n93954, n93955, n93956, n93957, n93958, n93959,
         n93960, n93961, n93962, n93963, n93964, n93965, n93966, n93967,
         n93968, n93969, n93970, n93971, n93972, n93973, n93974, n93975,
         n93976, n93977, n93978, n93979, n93980, n93981, n93982, n93983,
         n93984, n93985, n93986, n93987, n93988, n93989, n93990, n93991,
         n93992, n93993, n93994, n93995, n93996, n93997, n93998, n93999,
         n94000, n94001, n94002, n94003, n94004, n94005, n94006, n94007,
         n94008, n94009, n94010, n94011, n94012, n94013, n94014, n94015,
         n94016, n94017, n94018, n94019, n94020, n94021, n94022, n94023,
         n94024, n94025, n94026, n94027, n94028, n94029, n94030, n94031,
         n94032, n94033, n94034, n94035, n94036, n94037, n94038, n94039,
         n94040, n94041, n94042, n94043, n94044, n94045, n94046, n94047,
         n94048, n94049, n94050, n94051, n94052, n94053, n94054, n94055,
         n94056, n94057, n94058, n94059, n94060, n94061, n94062, n94063,
         n94064, n94065, n94066, n94067, n94068, n94069, n94070, n94071,
         n94072, n94073, n94074, n94075, n94076, n94077, n94078, n94079,
         n94080, n94081, n94082, n94083, n94084, n94085, n94086, n94087,
         n94088, n94089, n94090, n94091, n94092, n94093, n94094, n94095,
         n94096, n94097, n94098, n94099, n94100, n94101, n94102, n94103,
         n94104, n94105, n94106, n94107, n94108, n94109, n94110, n94111,
         n94112, n94113, n94114, n94115, n94116, n94117, n94118, n94119,
         n94120, n94121, n94122, n94123, n94124, n94125, n94126, n94127,
         n94128, n94129, n94130, n94131, n94132, n94133, n94134, n94135,
         n94136, n94137, n94138, n94139, n94140, n94141, n94142, n94143,
         n94144, n94145, n94146, n94147, n94148, n94149, n94150, n94151,
         n94152, n94153, n94154, n94155, n94156, n94157, n94158, n94159,
         n94160, n94161, n94162, n94163, n94164, n94165, n94166, n94167,
         n94168, n94169, n94170, n94171, n94172, n94173, n94174, n94175,
         n94176, n94177, n94178, n94179, n94180, n94181, n94182, n94183,
         n94184, n94185, n94186, n94187, n94188, n94189, n94190, n94191,
         n94192, n94193, n94194, n94195, n94196, n94197, n94198, n94199,
         n94200, n94201, n94202, n94203, n94204, n94205, n94206, n94207,
         n94208, n94209, n94210, n94211, n94212, n94213, n94214, n94215,
         n94216, n94217, n94218, n94219, n94220, n94221, n94222, n94223,
         n94224, n94225, n94226, n94227, n94228, n94229, n94230, n94231,
         n94232, n94233, n94234, n94235, n94236, n94237, n94238, n94239,
         n94240, n94241, n94242, n94243, n94244, n94245, n94246, n94247,
         n94248, n94249, n94250, n94251, n94252, n94253, n94254, n94256,
         n94257, n94258, n94259, n94260, n94261, n94262, n94263, n94264,
         n94265, n94266, n94267, n94268, n94269, n94270, n94271, n94272,
         n94273, n94274, n94275, n94276, n94277, n94278, n94279, n94280,
         n94281, n94282, n94283, n94284, n94285, n94286, n94287, n94288,
         n94289, n94290, n94291, n94292, n94293, n94294, n94295, n94296,
         n94297, n94298, n94299, n94300, n94301, n94302, n94303, n94304,
         n94305, n94306, n94307, n94308, n94309, n94310, n94311, n94312,
         n94313, n94314, n94315, n94316, n94317, n94318, n94319, n94320,
         n94321, n94322, n94323, n94324, n94325, n94326, n94327, n94328,
         n94329, n94330, n94331, n94332, n94333, n94334, n94335, n94336,
         n94337, n94338, n94339, n94340, n94341, n94342, n94343, n94344,
         n94345, n94346, n94347, n94348, n94349, n94350, n94351, n94352,
         n94353, n94354, n94355, n94356, n94357, n94358, n94359, n94360,
         n94361, n94362, n94363, n94364, n94365, n94366, n94367, n94368,
         n94369, n94370, n94371, n94372, n94373, n94374, n94375, n94376,
         n94377, n94378, n94379, n94380, n94381, n94382, n94383, n94384,
         n94385, n94386, n94387, n94388, n94389, n94390, n94391, n94392,
         n94393, n94394, n94395, n94396, n94397, n94398, n94399, n94400,
         n94401, n94402, n94403, n94404, n94405, n94406, n94407, n94408,
         n94409, n94410, n94411, n94412, n94413, n94414, n94415, n94416,
         n94417, n94418, n94419, n94420, n94421, n94422, n94423, n94424,
         n94425, n94426, n94427, n94428, n94429, n94430, n94431, n94432,
         n94433, n94434, n94435, n94436, n94437, n94438, n94439, n94440,
         n94441, n94442, n94443, n94444, n94445, n94446, n94447, n94448,
         n94449, n94450, n94451, n94452, n94453, n94454, n94455, n94456,
         n94457, n94458, n94459, n94460, n94461, n94462, n94463, n94464,
         n94465, n94466, n94467, n94468, n94469, n94470, n94471, n94472,
         n94473, n94474, n94475, n94476, n94477, n94478, n94479, n94480,
         n94481, n94482, n94483, n94484, n94485, n94486, n94487, n94488,
         n94489, n94490, n94491, n94492, n94493, n94494, n94495, n94496,
         n94497, n94498, n94499, n94500, n94501, n94502, n94503, n94504,
         n94505, n94506, n94507, n94508, n94509, n94510, n94511, n94512,
         n94513, n94514, n94515, n94516, n94517, n94518, n94519, n94520,
         n94521, n94522, n94523, n94524, n94525, n94526, n94527, n94528,
         n94529, n94530, n94531, n94532, n94533, n94534, n94535, n94536,
         n94537, n94538, n94539, n94540, n94541, n94542, n94543, n94544,
         n94545, n94546, n94547, n94548, n94549, n94550, n94551, n94552,
         n94553, n94554, n94555, n94556, n94557, n94558, n94559, n94561,
         n94562, n94563, n94564, n94565, n94566, n94567, n94568, n94569,
         n94570, n94571, n94572, n94573, n94574, n94575, n94576, n94577,
         n94578, n94579, n94580, n94581, n94582, n94583, n94584, n94585,
         n94586, n94587, n94588, n94589, n94590, n94591, n94592, n94593,
         n94594, n94595, n94596, n94597, n94598, n94599, n94600, n94601,
         n94602, n94603, n94604, n94605, n94606, n94607, n94608, n94609,
         n94610, n94611, n94612, n94613, n94614, n94615, n94616, n94617,
         n94618, n94619, n94620, n94621, n94622, n94623, n94624, n94625,
         n94626, n94627, n94628, n94630, n94631, n94632, n94633, n94634,
         n94635, n94636, n94637, n94638, n94639, n94640, n94641, n94642,
         n94643, n94644, n94645, n94646, n94647, n94648, n94649, n94650,
         n94651, n94652, n94653, n94654, n94655, n94656, n94657, n94658,
         n94659, n94660, n94661, n94662, n94663, n94664, n94665, n94666,
         n94667, n94668, n94669, n94670, n94671, n94672, n94673, n94674,
         n94675, n94676, n94677, n94678, n94679, n94680, n94681, n94682,
         n94683, n94684, n94685, n94686, n94687, n94688, n94689, n94690,
         n94691, n94692, n94693, n94694, n94695, n94696, n94697, n94698,
         n94699, n94700, n94701, n94702, n94703, n94704, n94705, n94706,
         n94707, n94708, n94709, n94710, n94711, n94712, n94713, n94714,
         n94715, n94716, n94717, n94718, n94719, n94720, n94721, n94722,
         n94723, n94724, n94725, n94726, n94727, n94728, n94729, n94730,
         n94731, n94732, n94733, n94734, n94735, n94736, n94737, n94739,
         n94740, n94741, n94742, n94743, n94744, n94745, n94746, n94747,
         n94748, n94749, n94750, n94751, n94752, n94753, n94754, n94755,
         n94756, n94757, n94758, n94759, n94760, n94761, n94762, n94763,
         n94764, n94765, n94766, n94767, n94768, n94769, n94770, n94771,
         n94772, n94773, n94774, n94775, n94776, n94777, n94778, n94779,
         n94780, n94781, n94782, n94783, n94784, n94785, n94786, n94787,
         n94788, n94789, n94790, n94791, n94792, n94793, n94794, n94795,
         n94796, n94797, n94798, n94799, n94800, n94801, n94802, n94803,
         n94804, n94805, n94806, n94807, n94808, n94809, n94810, n94812,
         n94813, n94814, n94815, n94816, n94817, n94818, n94819, n94820,
         n94821, n94822, n94823, n94824, n94825, n94826, n94827, n94828,
         n94829, n94830, n94831, n94832, n94833, n94834, n94835, n94836,
         n94837, n94838, n94839, n94840, n94841, n94842, n94843, n94844,
         n94845, n94847, n94848, n94849, n94850, n94851, n94852, n94853,
         n94854, n94855, n94856, n94857, n94858, n94859, n94860, n94861,
         n94862, n94863, n94864, n94865, n94866, n94867, n94868, n94869,
         n94870, n94871, n94872, n94873, n94874, n94875, n94876, n94877,
         n94878, n94879, n94880, n94881, n94882, n94883, n94884, n94885,
         n94886, n94887, n94888, n94889, n94890, n94892, n94893, n94894,
         n94895, n94896, n94897, n94898, n94899, n94900, n94901, n94902,
         n94903, n94904, n94905, n94906, n94907, n94908, n94909, n94910,
         n94911, n94912, n94913, n94914, n94915, n94916, n94917, n94918,
         n94919, n94920, n94921, n94922, n94923, n94924, n94925, n94926,
         n94927, n94928, n94929, n94930, n94931, n94932, n94933, n94934,
         n94935, n94936, n94937, n94938, n94939, n94940, n94941, n94942,
         n94943, n94944, n94945, n94946, n94947, n94948, n94949, n94950,
         n94951, n94952, n94953, n94954, n94955, n94956, n94957, n94958,
         n94959, n94960, n94961, n94962, n94963, n94964, n94965, n94966,
         n94967, n94968, n94969, n94970, n94971, n94972, n94973, n94974,
         n94975, n94976, n94977, n94978, n94979, n94980, n94981, n94982,
         n94983, n94984, n94985, n94986, n94987, n94988, n94989, n94990,
         n94991, n94992, n94993, n94994, n94995, n94996, n94997, n94998,
         n94999, n95000, n95001, n95003, n95004, n95005, n95006, n95007,
         n95008, n95009, n95010, n95011, n95012, n95013, n95014, n95015,
         n95016, n95017, n95018, n95019, n95020, n95021, n95022, n95023,
         n95024, n95025, n95026, n95027, n95028, n95029, n95030, n95031,
         n95032, n95033, n95034, n95035, n95036, n95037, n95038, n95039,
         n95040, n95041, n95042, n95043, n95044, n95045, n95046, n95047,
         n95048, n95049, n95050, n95051, n95052, n95053, n95054, n95055,
         n95056, n95057, n95058, n95059, n95060, n95061, n95062, n95063,
         n95064, n95065, n95066, n95067, n95068, n95069, n95070, n95071,
         n95072, n95073, n95074, n95075, n95076, n95077, n95078, n95079,
         n95080, n95081, n95082, n95083, n95084, n95085, n95086, n95087,
         n95088, n95089, n95090, n95091, n95092, n95093, n95094, n95095,
         n95096, n95097, n95098, n95099, n95100, n95101, n95102, n95103,
         n95104, n95105, n95106, n95107, n95108, n95109, n95110, n95111,
         n95112, n95113, n95114, n95115, n95116, n95117, n95118, n95119,
         n95120, n95121, n95122, n95123, n95124, n95125, n95126, n95127,
         n95128, n95129, n95130, n95131, n95132, n95133, n95134, n95136,
         n95137, n95138, n95139, n95140, n95141, n95142, n95143, n95144,
         n95145, n95146, n95147, n95148, n95149, n95150, n95151, n95152,
         n95153, n95154, n95155, n95156, n95157, n95158, n95159, n95160,
         n95161, n95162, n95163, n95164, n95165, n95166, n95167, n95168,
         n95169, n95170, n95171, n95172, n95173, n95174, n95175, n95176,
         n95177, n95178, n95179, n95180, n95181, n95182, n95183, n95184,
         n95185, n95186, n95187, n95188, n95189, n95190, n95191, n95192,
         n95193, n95194, n95195, n95196, n95197, n95198, n95199, n95200,
         n95201, n95202, n95203, n95204, n95205, n95206, n95207, n95208,
         n95209, n95210, n95211, n95212, n95213, n95214, n95215, n95216,
         n95217, n95218, n95219, n95220, n95221, n95222, n95223, n95224,
         n95225, n95226, n95227, n95228, n95229, n95230, n95231, n95232,
         n95233, n95234, n95235, n95236, n95237, n95238, n95239, n95240,
         n95241, n95242, n95243, n95244, n95245, n95246, n95247, n95248,
         n95249, n95250, n95251, n95252, n95253, n95254, n95255, n95256,
         n95257, n95258, n95259, n95260, n95261, n95262, n95263, n95264,
         n95265, n95266, n95267, n95268, n95269, n95270, n95271, n95272,
         n95273, n95274, n95275, n95276, n95277, n95278, n95279, n95280,
         n95281, n95282, n95283, n95284, n95285, n95286, n95287, n95288,
         n95289, n95290, n95291, n95292, n95293, n95294, n95295, n95296,
         n95297, n95298, n95299, n95300, n95301, n95302, n95303, n95304,
         n95305, n95306, n95307, n95308, n95309, n95310, n95311, n95312,
         n95313, n95314, n95315, n95316, n95317, n95318, n95319, n95320,
         n95321, n95322, n95323, n95324, n95325, n95326, n95327, n95328,
         n95329, n95330, n95331, n95332, n95333, n95334, n95335, n95336,
         n95337, n95338, n95339, n95340, n95341, n95342, n95343, n95344,
         n95345, n95346, n95347, n95348, n95349, n95350, n95351, n95352,
         n95353, n95354, n95355, n95356, n95357, n95358, n95359, n95360,
         n95361, n95362, n95363, n95364, n95365, n95366, n95367, n95368,
         n95369, n95370, n95371, n95372, n95373, n95374, n95375, n95376,
         n95377, n95378, n95379, n95380, n95381, n95382, n95383, n95384,
         n95385, n95386, n95387, n95388, n95389, n95390, n95391, n95392,
         n95393, n95394, n95395, n95396, n95397, n95398, n95399, n95400,
         n95401, n95402, n95403, n95404, n95405, n95406, n95407, n95408,
         n95409, n95410, n95411, n95412, n95413, n95414, n95415, n95417,
         n95418, n95419, n95420, n95421, n95422, n95423, n95424, n95425,
         n95426, n95427, n95428, n95429, n95430, n95431, n95432, n95433,
         n95434, n95435, n95436, n95437, n95438, n95439, n95440, n95441,
         n95442, n95443, n95444, n95445, n95446, n95447, n95448, n95449,
         n95450, n95451, n95452, n95453, n95454, n95455, n95457, n95458,
         n95459, n95460, n95461, n95462, n95463, n95464, n95465, n95466,
         n95467, n95468, n95469, n95470, n95471, n95472, n95473, n95474,
         n95475, n95476, n95477, n95478, n95479, n95480, n95481, n95482,
         n95483, n95484, n95485, n95486, n95487, n95488, n95489, n95490,
         n95491, n95492, n95493, n95494, n95495, n95496, n95497, n95498,
         n95499, n95500, n95501, n95502, n95503, n95504, n95505, n95506,
         n95507, n95508, n95509, n95510, n95511, n95512, n95513, n95514,
         n95515, n95516, n95517, n95518, n95519, n95520, n95521, n95522,
         n95523, n95524, n95525, n95526, n95527, n95528, n95529, n95530,
         n95531, n95532, n95533, n95534, n95535, n95536, n95537, n95538,
         n95539, n95540, n95541, n95542, n95543, n95544, n95545, n95546,
         n95547, n95548, n95549, n95550, n95551, n95552, n95553, n95554,
         n95555, n95556, n95557, n95558, n95559, n95560, n95561, n95562,
         n95563, n95564, n95565, n95566, n95567, n95568, n95569, n95570,
         n95571, n95572, n95573, n95574, n95575, n95576, n95577, n95578,
         n95579, n95580, n95581, n95582, n95583, n95584, n95585, n95586,
         n95587, n95588, n95589, n95590, n95591, n95592, n95593, n95594,
         n95595, n95596, n95597, n95598, n95599, n95600, n95601, n95602,
         n95603, n95604, n95605, n95606, n95607, n95608, n95609, n95610,
         n95611, n95612, n95613, n95614, n95615, n95616, n95617, n95618,
         n95619, n95620, n95621, n95622, n95623, n95624, n95625, n95626,
         n95627, n95628, n95629, n95630, n95631, n95632, n95633, n95634,
         n95635, n95636, n95637, n95638, n95639, n95640, n95641, n95642,
         n95643, n95644, n95645, n95646, n95647, n95648, n95649, n95650,
         n95651, n95652, n95653, n95654, n95655, n95656, n95657, n95658,
         n95659, n95660, n95661, n95662, n95663, n95664, n95665, n95666,
         n95667, n95668, n95669, n95670, n95671, n95672, n95673, n95674,
         n95675, n95676, n95677, n95678, n95679, n95680, n95681, n95682,
         n95683, n95684, n95685, n95686, n95687, n95688, n95689, n95690,
         n95691, n95694, n95695, n95696, n95697, n95698, n95699, n95700,
         n95701, n95702, n95703, n95704, n95705, n95706, n95707, n95708,
         n95709, n95710, n95711, n95712, n95713, n95714, n95715, n95716,
         n95717, n95718, n95719, n95720, n95721, n95722, n95723, n95724,
         n95725, n95726, n95727, n95728, n95729, n95731, n95732, n95733,
         n95734, n95735, n95736, n95737, n95738, n95739, n95740, n95741,
         n95742, n95743, n95744, n95745, n95746, n95747, n95748, n95749,
         n95750, n95751, n95752, n95753, n95754, n95755, n95756, n95757,
         n95758, n95759, n95760, n95761, n95762, n95763, n95764, n95765,
         n95768, n95769, n95770, n95771, n95772, n95773, n95774, n95775,
         n95776, n95777, n95778, n95779, n95780, n95781, n95782, n95783,
         n95784, n95785, n95786, n95787, n95788, n95789, n95790, n95791,
         n95792, n95793, n95794, n95795, n95796, n95797, n95798, n95799,
         n95800, n95801, n95802, n95803, n95804, n95805, n95806, n95807,
         n95808, n95809, n95810, n95811, n95812, n95813, n95814, n95815,
         n95816, n95817, n95818, n95819, n95820, n95821, n95822, n95823,
         n95824, n95825, n95826, n95827, n95828, n95829, n95830, n95831,
         n95832, n95833, n95834, n95835, n95836, n95837, n95838, n95839,
         n95840, n95841, n95842, n95843, n95844, n95845, n95846, n95847,
         n95848, n95849, n95850, n95851, n95852, n95853, n95854, n95855,
         n95856, n95857, n95858, n95859, n95860, n95861, n95862, n95863,
         n95864, n95865, n95866, n95867, n95868, n95869, n95870, n95871,
         n95872, n95873, n95874, n95875, n95876, n95878, n95879, n95880,
         n95881, n95882, n95883, n95884, n95885, n95886, n95887, n95888,
         n95889, n95890, n95891, n95892, n95893, n95894, n95895, n95896,
         n95897, n95898, n95899, n95900, n95901, n95902, n95903, n95904,
         n95905, n95906, n95907, n95908, n95909, n95911, n95912, n95913,
         n95914, n95915, n95917, n95918, n95919, n95920, n95921, n95922,
         n95923, n95924, n95925, n95926, n95927, n95928, n95929, n95930,
         n95931, n95932, n95933, n95934, n95935, n95936, n95937, n95938,
         n95939, n95940, n95941, n95942, n95943, n95944, n95945, n95946,
         n95947, n95948, n95949, n95950, n95951, n95952, n95953, n95955,
         n95956, n95957, n95958, n95959, n95960, n95961, n95962, n95963,
         n95964, n95965, n95966, n95967, n95968, n95969, n95970, n95971,
         n95972, n95973, n95974, n95975, n95976, n95977, n95978, n95979,
         n95980, n95981, n95982, n95983, n95984, n95985, n95986, n95987,
         n95988, n95989, n95990, n95991, n95992, n95993, n95994, n95995,
         n95996, n95997, n95998, n95999, n96000, n96001, n96002, n96003,
         n96004, n96005, n96006, n96007, n96008, n96009, n96010, n96011,
         n96012, n96013, n96014, n96015, n96016, n96017, n96019, n96020,
         n96021, n96022, n96023, n96024, n96025, n96026, n96027, n96028,
         n96029, n96030, n96031, n96032, n96033, n96034, n96035, n96036,
         n96037, n96038, n96039, n96040, n96041, n96042, n96043, n96044,
         n96045, n96046, n96047, n96048, n96049, n96050, n96051, n96052,
         n96053, n96054, n96056, n96057, n96058, n96059, n96060, n96061,
         n96062, n96063, n96064, n96065, n96066, n96067, n96068, n96069,
         n96070, n96071, n96072, n96073, n96074, n96075, n96076, n96077,
         n96078, n96079, n96080, n96081, n96082, n96083, n96084, n96085,
         n96086, n96087, n96088, n96089, n96090, n96091, n96092, n96093,
         n96095, n96096, n96097, n96098, n96099, n96100, n96101, n96102,
         n96103, n96104, n96105, n96106, n96107, n96108, n96109, n96110,
         n96111, n96112, n96113, n96114, n96115, n96116, n96117, n96118,
         n96119, n96120, n96121, n96122, n96123, n96124, n96125, n96126,
         n96127, n96128, n96129, n96130, n96131, n96132, n96133, n96135,
         n96136, n96137, n96138, n96139, n96140, n96141, n96142, n96143,
         n96144, n96145, n96146, n96147, n96148, n96149, n96150, n96151,
         n96152, n96153, n96154, n96155, n96156, n96157, n96158, n96159,
         n96160, n96161, n96162, n96163, n96164, n96165, n96166, n96167,
         n96168, n96169, n96172, n96173, n96174, n96175, n96176, n96177,
         n96178, n96179, n96180, n96181, n96182, n96183, n96184, n96185,
         n96186, n96187, n96188, n96189, n96190, n96191, n96192, n96193,
         n96194, n96195, n96196, n96197, n96198, n96199, n96200, n96201,
         n96202, n96203, n96204, n96205, n96206, n96207, n96208, n96209,
         n96210, n96211, n96212, n96213, n96214, n96215, n96216, n96217,
         n96218, n96219, n96220, n96221, n96222, n96223, n96224, n96225,
         n96226, n96227, n96228, n96229, n96230, n96231, n96232, n96233,
         n96234, n96236, n96237, n96238, n96239, n96240, n96241, n96242,
         n96243, n96244, n96245, n96246, n96247, n96248, n96249, n96250,
         n96251, n96252, n96253, n96254, n96255, n96256, n96257, n96258,
         n96259, n96260, n96261, n96262, n96263, n96264, n96265, n96266,
         n96267, n96268, n96269, n96270, n96271, n96272, n96273, n96274,
         n96275, n96276, n96277, n96278, n96279, n96280, n96281, n96282,
         n96283, n96284, n96285, n96286, n96287, n96288, n96289, n96290,
         n96291, n96292, n96293, n96294, n96295, n96296, n96299, n96300,
         n96301, n96302, n96303, n96304, n96305, n96306, n96307, n96308,
         n96309, n96310, n96311, n96312, n96313, n96314, n96315, n96316,
         n96317, n96318, n96319, n96320, n96321, n96322, n96323, n96324,
         n96325, n96326, n96327, n96328, n96329, n96330, n96331, n96332,
         n96333, n96334, n96335, n96336, n96337, n96338, n96339, n96340,
         n96341, n96342, n96343, n96344, n96345, n96346, n96347, n96348,
         n96349, n96350, n96351, n96352, n96353, n96354, n96355, n96356,
         n96357, n96358, n96359, n96360, n96361, n96362, n96363, n96364,
         n96365, n96366, n96367, n96368, n96369, n96370, n96371, n96372,
         n96373, n96374, n96375, n96376, n96377, n96378, n96379, n96380,
         n96381, n96382, n96383, n96384, n96385, n96386, n96387, n96388,
         n96389, n96390, n96391, n96392, n96393, n96394, n96395, n96396,
         n96397, n96398, n96399, n96400, n96401, n96402, n96403, n96404,
         n96405, n96406, n96407, n96408, n96409, n96410, n96411, n96412,
         n96413, n96414, n96415, n96416, n96417, n96418, n96419, n96422,
         n96423, n96424, n96425, n96426, n96427, n96428, n96429, n96430,
         n96431, n96432, n96433, n96434, n96435, n96436, n96437, n96438,
         n96439, n96440, n96441, n96442, n96443, n96444, n96445, n96446,
         n96447, n96448, n96449, n96450, n96451, n96452, n96453, n96454,
         n96455, n96456, n96457, n96458, n96459, n96460, n96461, n96462,
         n96463, n96464, n96465, n96466, n96467, n96468, n96469, n96470,
         n96471, n96472, n96473, n96474, n96475, n96476, n96477, n96478,
         n96479, n96480, n96481, n96482, n96483, n96484, n96485, n96486,
         n96487, n96488, n96489, n96491, n96493, n96494, n96495, n96496,
         n96497, n96498, n96499, n96500, n96501, n96502, n96503, n96504,
         n96505, n96506, n96507, n96508, n96509, n96510, n96511, n96512,
         n96513, n96514, n96515, n96516, n96517, n96518, n96519, n96520,
         n96521, n96522, n96523, n96524, n96525, n96526, n96527, n96528,
         n96529, n96530, n96531, n96532, n96533, n96534, n96535, n96536,
         n96537, n96538, n96539, n96540, n96541, n96542, n96543, n96544,
         n96545, n96546, n96547, n96548, n96549, n96550, n96551, n96552,
         n96553, n96554, n96555, n96556, n96557, n96558, n96559, n96560,
         n96561, n96562, n96563, n96564, n96565, n96566, n96567, n96568,
         n96569, n96570, n96571, n96572, n96573, n96574, n96575, n96576,
         n96577, n96578, n96579, n96580, n96581, n96582, n96583, n96584,
         n96585, n96586, n96587, n96588, n96589, n96590, n96591, n96592,
         n96593, n96594, n96595, n96596, n96597, n96598, n96599, n96600,
         n96601, n96602, n96603, n96604, n96605, n96606, n96607, n96608,
         n96609, n96610, n96611, n96612, n96613, n96614, n96615, n96616,
         n96617, n96618, n96619, n96620, n96621, n96622, n96623, n96624,
         n96625, n96626, n96627, n96628, n96629, n96630, n96631, n96632,
         n96633, n96634, n96635, n96636, n96637, n96638, n96639, n96640,
         n96641, n96642, n96643, n96644, n96645, n96646, n96647, n96648,
         n96649, n96650, n96651, n96652, n96653, n96654, n96655, n96656,
         n96657, n96658, n96659, n96660, n96661, n96662, n96663, n96664,
         n96665, n96666, n96667, n96668, n96669, n96670, n96671, n96672,
         n96673, n96674, n96675, n96676, n96677, n96678, n96679, n96680,
         n96681, n96682, n96683, n96684, n96685, n96686, n96687, n96688,
         n96689, n96690, n96691, n96692, n96693, n96694, n96695, n96696,
         n96697, n96698, n96699, n96700, n96701, n96702, n96703, n96704,
         n96705, n96706, n96707, n96708, n96709, n96710, n96711, n96712,
         n96713, n96714, n96715, n96716, n96717, n96718, n96719, n96720,
         n96721, n96722, n96723, n96724, n96725, n96726, n96727, n96728,
         n96729, n96730, n96731, n96732, n96733, n96734, n96735, n96736,
         n96737, n96738, n96739, n96740, n96741, n96742, n96743, n96744,
         n96745, n96746, n96747, n96748, n96749, n96750, n96751, n96752,
         n96753, n96754, n96755, n96756, n96757, n96758, n96759, n96760,
         n96761, n96762, n96763, n96764, n96765, n96766, n96767, n96768,
         n96769, n96770, n96771, n96772, n96773, n96774, n96775, n96776,
         n96777, n96778, n96779, n96780, n96781, n96782, n96783, n96784,
         n96785, n96786, n96787, n96788, n96789, n96790, n96791, n96792,
         n96793, n96794, n96795, n96796, n96797, n96798, n96799, n96800,
         n96801, n96802, n96803, n96804, n96805, n96806, n96807, n96808,
         n96809, n96810, n96811, n96812, n96813, n96814, n96815, n96816,
         n96817, n96818, n96819, n96820, n96821, n96822, n96823, n96824,
         n96825, n96826, n96827, n96828, n96829, n96830, n96831, n96832,
         n96833, n96834, n96835, n96836, n96837, n96838, n96839, n96840,
         n96841, n96842, n96843, n96844, n96845, n96846, n96847, n96848,
         n96849, n96850, n96851, n96852, n96853, n96854, n96855, n96856,
         n96857, n96858, n96859, n96860, n96861, n96862, n96863, n96864,
         n96865, n96866, n96867, n96868, n96869, n96870, n96871, n96872,
         n96873, n96874, n96875, n96876, n96877, n96879, n96880, n96881,
         n96882, n96883, n96884, n96885, n96886, n96887, n96888, n96889,
         n96890, n96891, n96892, n96893, n96894, n96895, n96896, n96897,
         n96898, n96899, n96900, n96901, n96902, n96903, n96904, n96905,
         n96906, n96907, n96908, n96909, n96910, n96911, n96912, n96913,
         n96914, n96915, n96916, n96917, n96918, n96919, n96920, n96921,
         n96922, n96923, n96924, n96925, n96926, n96927, n96928, n96929,
         n96930, n96931, n96932, n96933, n96934, n96935, n96936, n96938,
         n96939, n96940, n96941, n96942, n96943, n96944, n96945, n96946,
         n96947, n96948, n96949, n96950, n96951, n96952, n96953, n96954,
         n96955, n96956, n96957, n96958, n96959, n96960, n96961, n96962,
         n96963, n96964, n96965, n96966, n96967, n96968, n96969, n96970,
         n96971, n96972, n96973, n96974, n96975, n96976, n96977, n96978,
         n96979, n96980, n96981, n96982, n96983, n96984, n96985, n96986,
         n96987, n96988, n96989, n96990, n96991, n96992, n96993, n96994,
         n96995, n96996, n96997, n96998, n96999, n97000, n97001, n97002,
         n97003, n97004, n97005, n97006, n97007, n97008, n97009, n97010,
         n97011, n97012, n97013, n97014, n97015, n97016, n97017, n97018,
         n97019, n97020, n97021, n97022, n97023, n97024, n97025, n97026,
         n97027, n97028, n97029, n97030, n97031, n97032, n97033, n97034,
         n97035, n97036, n97037, n97038, n97039, n97040, n97041, n97042,
         n97043, n97044, n97045, n97046, n97047, n97048, n97049, n97050,
         n97051, n97052, n97053, n97054, n97055, n97056, n97057, n97058,
         n97059, n97060, n97061, n97062, n97063, n97064, n97065, n97066,
         n97067, n97068, n97069, n97070, n97071, n97072, n97073, n97074,
         n97075, n97076, n97077, n97078, n97079, n97080, n97081, n97082,
         n97083, n97084, n97085, n97086, n97087, n97088, n97089, n97090,
         n97091, n97092, n97093, n97094, n97095, n97096, n97097, n97098,
         n97099, n97100, n97101, n97102, n97103, n97104, n97105, n97106,
         n97107, n97108, n97109, n97110, n97111, n97112, n97113, n97114,
         n97115, n97116, n97117, n97118, n97119, n97120, n97121, n97122,
         n97123, n97124, n97125, n97126, n97127, n97128, n97129, n97130,
         n97131, n97132, n97133, n97134, n97135, n97136, n97137, n97138,
         n97139, n97140, n97141, n97142, n97143, n97144, n97145, n97146,
         n97147, n97148, n97149, n97150, n97151, n97152, n97153, n97154,
         n97155, n97156, n97157, n97158, n97159, n97160, n97161, n97162,
         n97163, n97164, n97165, n97166, n97167, n97168, n97169, n97170,
         n97171, n97172, n97173, n97174, n97175, n97176, n97177, n97178,
         n97179, n97180, n97181, n97182, n97183, n97184, n97185, n97186,
         n97187, n97188, n97189, n97190, n97191, n97192, n97193, n97194,
         n97195, n97196, n97197, n97198, n97199, n97200, n97201, n97202,
         n97203, n97204, n97205, n97206, n97207, n97208, n97209, n97210,
         n97211, n97212, n97213, n97214, n97215, n97216, n97217, n97218,
         n97219, n97220, n97221, n97222, n97223, n97224, n97225, n97226,
         n97227, n97228, n97229, n97230, n97231, n97232, n97233, n97234,
         n97235, n97236, n97237, n97238, n97239, n97240, n97241, n97242,
         n97243, n97244, n97245, n97246, n97247, n97248, n97249, n97250,
         n97251, n97252, n97253, n97254, n97255, n97256, n97257, n97258,
         n97259, n97260, n97261, n97262, n97263, n97264, n97265, n97266,
         n97267, n97268, n97269, n97270, n97271, n97272, n97273, n97274,
         n97275, n97276, n97277, n97278, n97279, n97280, n97281, n97282,
         n97283, n97284, n97285, n97286, n97287, n97288, n97289, n97290,
         n97291, n97292, n97293, n97294, n97295, n97296, n97297, n97298,
         n97299, n97300, n97301, n97302, n97303, n97304, n97305, n97306,
         n97307, n97308, n97309, n97310, n97311, n97312, n97313, n97314,
         n97315, n97316, n97317, n97318, n97320, n97321, n97322, n97323,
         n97324, n97325, n97326, n97327, n97328, n97329, n97330, n97331,
         n97332, n97333, n97334, n97335, n97336, n97337, n97338, n97339,
         n97340, n97341, n97342, n97343, n97344, n97345, n97346, n97347,
         n97348, n97349, n97350, n97351, n97352, n97353, n97354, n97355,
         n97356, n97357, n97358, n97359, n97360, n97361, n97362, n97363,
         n97364, n97365, n97366, n97367, n97368, n97369, n97370, n97371,
         n97372, n97373, n97374, n97375, n97376, n97377, n97378, n97379,
         n97380, n97381, n97382, n97383, n97384, n97385, n97386, n97387,
         n97388, n97389, n97390, n97391, n97392, n97393, n97394, n97395,
         n97396, n97397, n97398, n97399, n97400, n97401, n97402, n97403,
         n97404, n97405, n97406, n97407, n97408, n97409, n97410, n97411,
         n97412, n97413, n97414, n97415, n97416, n97417, n97418, n97419,
         n97420, n97421, n97422, n97423, n97424, n97425, n97426, n97427,
         n97428, n97429, n97430, n97431, n97432, n97433, n97434, n97435,
         n97436, n97437, n97438, n97439, n97440, n97441, n97442, n97443,
         n97444, n97445, n97446, n97447, n97448, n97449, n97450, n97451,
         n97452, n97453, n97454, n97455, n97456, n97457, n97458, n97459,
         n97460, n97461, n97462, n97463, n97464, n97465, n97466, n97467,
         n97468, n97469, n97470, n97471, n97472, n97473, n97474, n97475,
         n97476, n97477, n97478, n97479, n97480, n97481, n97482, n97483,
         n97484, n97485, n97486, n97487, n97488, n97489, n97490, n97491,
         n97492, n97493, n97494, n97495, n97496, n97497, n97498, n97499,
         n97500, n97501, n97502, n97503, n97504, n97505, n97506, n97507,
         n97508, n97509, n97510, n97511, n97512, n97513, n97514, n97515,
         n97516, n97517, n97518, n97519, n97520, n97521, n97522, n97523,
         n97524, n97525, n97526, n97527, n97528, n97529, n97530, n97531,
         n97532, n97533, n97534, n97535, n97536, n97537, n97538, n97539,
         n97540, n97541, n97542, n97543, n97544, n97545, n97546, n97547,
         n97548, n97549, n97550, n97551, n97552, n97553, n97554, n97555,
         n97556, n97557, n97558, n97559, n97560, n97561, n97562, n97563,
         n97564, n97565, n97566, n97567, n97568, n97569, n97570, n97571,
         n97572, n97573, n97574, n97575, n97576, n97577, n97578, n97579,
         n97580, n97581, n97582, n97583, n97584, n97585, n97586, n97587,
         n97588, n97589, n97590, n97591, n97592, n97593, n97594, n97595,
         n97596, n97597, n97598, n97599, n97600, n97601, n97602, n97603,
         n97604, n97605, n97606, n97607, n97608, n97609, n97610, n97611,
         n97612, n97613, n97614, n97615, n97616, n97617, n97618, n97619,
         n97620, n97621, n97622, n97623, n97624, n97625, n97626, n97627,
         n97628, n97629, n97630, n97631, n97632, n97633, n97634, n97635,
         n97636, n97637, n97638, n97639, n97641, n97642, n97643, n97644,
         n97645, n97646, n97647, n97648, n97649, n97650, n97651, n97652,
         n97653, n97654, n97655, n97656, n97657, n97658, n97659, n97660,
         n97661, n97662, n97663, n97664, n97665, n97666, n97667, n97668,
         n97669, n97670, n97671, n97672, n97673, n97674, n97675, n97676,
         n97677, n97679, n97680, n97681, n97682, n97683, n97684, n97685,
         n97686, n97687, n97688, n97689, n97690, n97691, n97692, n97693,
         n97694, n97695, n97696, n97697, n97698, n97699, n97700, n97701,
         n97702, n97703, n97704, n97705, n97706, n97707, n97708, n97709,
         n97710, n97711, n97712, n97713, n97714, n97715, n97716, n97717,
         n97718, n97719, n97720, n97721, n97722, n97723, n97724, n97725,
         n97726, n97727, n97728, n97729, n97730, n97731, n97732, n97733,
         n97734, n97735, n97736, n97737, n97738, n97739, n97740, n97741,
         n97742, n97743, n97744, n97745, n97746, n97747, n97748, n97749,
         n97750, n97751, n97752, n97753, n97754, n97755, n97756, n97757,
         n97758, n97759, n97760, n97761, n97762, n97763, n97764, n97765,
         n97766, n97767, n97768, n97769, n97770, n97771, n97772, n97773,
         n97774, n97775, n97776, n97777, n97778, n97779, n97780, n97781,
         n97782, n97783, n97784, n97785, n97786, n97787, n97788, n97789,
         n97790, n97791, n97792, n97793, n97794, n97795, n97796, n97797,
         n97798, n97799, n97800, n97801, n97802, n97803, n97804, n97805,
         n97806, n97807, n97808, n97809, n97810, n97811, n97812, n97813,
         n97814, n97815, n97816, n97817, n97818, n97819, n97820, n97821,
         n97822, n97823, n97824, n97825, n97826, n97827, n97828, n97829,
         n97830, n97831, n97832, n97833, n97834, n97835, n97836, n97837,
         n97838, n97839, n97840, n97841, n97842, n97843, n97844, n97845,
         n97846, n97847, n97848, n97849, n97850, n97851, n97852, n97853,
         n97854, n97855, n97856, n97857, n97858, n97859, n97860, n97861,
         n97862, n97863, n97864, n97865, n97866, n97867, n97868, n97869,
         n97870, n97871, n97872, n97873, n97874, n97875, n97876, n97877,
         n97878, n97879, n97880, n97881, n97882, n97883, n97884, n97885,
         n97886, n97887, n97888, n97889, n97890, n97891, n97892, n97893,
         n97894, n97895, n97896, n97897, n97898, n97899, n97900, n97901,
         n97902, n97903, n97904, n97905, n97906, n97907, n97908, n97909,
         n97910, n97911, n97912, n97913, n97914, n97915, n97916, n97917,
         n97918, n97919, n97920, n97921, n97922, n97923, n97924, n97925,
         n97926, n97927, n97928, n97929, n97930, n97931, n97932, n97933,
         n97934, n97935, n97936, n97937, n97938, n97939, n97940, n97941,
         n97942, n97943, n97944, n97945, n97946, n97947, n97948, n97949,
         n97950, n97951, n97952, n97953, n97954, n97955, n97956, n97957,
         n97958, n97959, n97960, n97961, n97962, n97963, n97964, n97965,
         n97966, n97967, n97968, n97969, n97970, n97973, n97974, n97975,
         n97976, n97977, n97978, n97979, n97980, n97981, n97982, n97983,
         n97984, n97985, n97986, n97987, n97988, n97989, n97990, n97991,
         n97992, n97993, n97994, n97995, n97996, n97997, n97998, n97999,
         n98000, n98001, n98002, n98003, n98004, n98005, n98006, n98007,
         n98008, n98009, n98010, n98011, n98012, n98013, n98014, n98015,
         n98016, n98017, n98018, n98019, n98020, n98021, n98022, n98023,
         n98024, n98025, n98026, n98027, n98028, n98029, n98030, n98031,
         n98032, n98033, n98034, n98035, n98036, n98037, n98038, n98039,
         n98040, n98041, n98042, n98043, n98044, n98045, n98046, n98047,
         n98048, n98049, n98050, n98051, n98052, n98053, n98054, n98055,
         n98056, n98057, n98058, n98059, n98060, n98061, n98062, n98063,
         n98064, n98065, n98066, n98067, n98068, n98069, n98070, n98071,
         n98072, n98073, n98074, n98075, n98076, n98077, n98078, n98079,
         n98080, n98081, n98082, n98083, n98084, n98085, n98086, n98087,
         n98088, n98089, n98090, n98091, n98092, n98093, n98094, n98095,
         n98096, n98097, n98098, n98099, n98100, n98101, n98102, n98103,
         n98104, n98105, n98106, n98107, n98108, n98109, n98110, n98111,
         n98112, n98113, n98114, n98115, n98116, n98117, n98118, n98119,
         n98120, n98121, n98122, n98123, n98124, n98125, n98126, n98127,
         n98128, n98129, n98130, n98131, n98132, n98133, n98134, n98135,
         n98136, n98137, n98138, n98139, n98140, n98141, n98142, n98143,
         n98144, n98145, n98146, n98147, n98148, n98149, n98150, n98151,
         n98152, n98153, n98154, n98155, n98156, n98157, n98158, n98159,
         n98160, n98161, n98162, n98163, n98164, n98165, n98166, n98167,
         n98168, n98169, n98170, n98171, n98172, n98173, n98174, n98175,
         n98176, n98177, n98178, n98179, n98180, n98181, n98182, n98183,
         n98184, n98185, n98186, n98187, n98188, n98189, n98190, n98191,
         n98192, n98193, n98194, n98195, n98196, n98197, n98198, n98199,
         n98200, n98201, n98202, n98203, n98204, n98205, n98206, n98207,
         n98208, n98209, n98210, n98211, n98212, n98213, n98214, n98215,
         n98216, n98217, n98218, n98219, n98220, n98221, n98222, n98223,
         n98224, n98225, n98226, n98227, n98228, n98229, n98230, n98231,
         n98232, n98233, n98234, n98235, n98236, n98237, n98238, n98239,
         n98240, n98241, n98242, n98243, n98244, n98245, n98246, n98247,
         n98248, n98249, n98250, n98251, n98252, n98253, n98254, n98255,
         n98256, n98257, n98258, n98259, n98260, n98261, n98262, n98263,
         n98264, n98265, n98266, n98267, n98268, n98269, n98270, n98271,
         n98272, n98273, n98274, n98275, n98276, n98277, n98278, n98279,
         n98280, n98281, n98282, n98283, n98284, n98285, n98286, n98287,
         n98288, n98289, n98290, n98291, n98292, n98293, n98294, n98295,
         n98296, n98297, n98298, n98299, n98300, n98301, n98302, n98303,
         n98304, n98305, n98306, n98307, n98308, n98309, n98310, n98311,
         n98312, n98313, n98314, n98315, n98316, n98317, n98318, n98319,
         n98320, n98321, n98322, n98323, n98324, n98325, n98326, n98327,
         n98328, n98329, n98330, n98331, n98332, n98333, n98334, n98335,
         n98336, n98337, n98338, n98339, n98340, n98341, n98342, n98343,
         n98344, n98345, n98346, n98347, n98348, n98349, n98350, n98351,
         n98352, n98353, n98354, n98355, n98356, n98357, n98358, n98359,
         n98360, n98361, n98362, n98363, n98364, n98365, n98366, n98367,
         n98368, n98369, n98370, n98371, n98372, n98373, n98374, n98375,
         n98376, n98377, n98378, n98379, n98380, n98381, n98382, n98383,
         n98384, n98385, n98386, n98387, n98388, n98389, n98390, n98391,
         n98392, n98393, n98394, n98395, n98396, n98397, n98398, n98399,
         n98400, n98401, n98402, n98403, n98404, n98405, n98406, n98407,
         n98408, n98409, n98410, n98411, n98412, n98413, n98414, n98415,
         n98416, n98417, n98418, n98419, n98420, n98421, n98422, n98423,
         n98424, n98425, n98426, n98427, n98428, n98429, n98430, n98431,
         n98432, n98433, n98434, n98435, n98436, n98437, n98438, n98439,
         n98440, n98441, n98442, n98443, n98444, n98445, n98446, n98447,
         n98448, n98449, n98450, n98451, n98452, n98453, n98454, n98455,
         n98456, n98457, n98458, n98459, n98460, n98461, n98462, n98463,
         n98464, n98465, n98466, n98467, n98468, n98469, n98470, n98471,
         n98472, n98473, n98474, n98475, n98476, n98477, n98478, n98479,
         n98480, n98481, n98482, n98483, n98484, n98485, n98486, n98487,
         n98488, n98489, n98490, n98491, n98492, n98493, n98494, n98495,
         n98496, n98497, n98498, n98499, n98500, n98501, n98502, n98503,
         n98504, n98505, n98506, n98507, n98508, n98509, n98510, n98511,
         n98512, n98513, n98514, n98515, n98516, n98517, n98518, n98519,
         n98520, n98521, n98522, n98523, n98524, n98525, n98526, n98527,
         n98528, n98529, n98530, n98531, n98532, n98533, n98534, n98535,
         n98536, n98537, n98538, n98539, n98540, n98541, n98542, n98543,
         n98544, n98545, n98546, n98547, n98548, n98549, n98550, n98551,
         n98552, n98553, n98554, n98555, n98556, n98557, n98558, n98559,
         n98560, n98561, n98562, n98563, n98564, n98565, n98566, n98567,
         n98568, n98569, n98570, n98571, n98572, n98573, n98574, n98575,
         n98576, n98577, n98578, n98579, n98580, n98581, n98582, n98583,
         n98584, n98585, n98586, n98587, n98588, n98589, n98590, n98591,
         n98592, n98593, n98594, n98595, n98596, n98597, n98598, n98599,
         n98600, n98601, n98602, n98603, n98604, n98605, n98606, n98607,
         n98608, n98609, n98610, n98611, n98612, n98613, n98614, n98615,
         n98616, n98617, n98618, n98619, n98620, n98621, n98622, n98623,
         n98624, n98625, n98626, n98627, n98628, n98629, n98630, n98631,
         n98632, n98633, n98634, n98635, n98636, n98637, n98638, n98639,
         n98640, n98641, n98642, n98643, n98644, n98645, n98646, n98647,
         n98648, n98649, n98650, n98651, n98652, n98653, n98654, n98655,
         n98656, n98657, n98658, n98659, n98660, n98661, n98662, n98663,
         n98664, n98665, n98666, n98667, n98668, n98669, n98670, n98671,
         n98672, n98673, n98674, n98675, n98676, n98677, n98678, n98679,
         n98680, n98681, n98682, n98683, n98684, n98685, n98686, n98687,
         n98688, n98689, n98690, n98691, n98692, n98693, n98694, n98695,
         n98696, n98697, n98698, n98699, n98700, n98701, n98702, n98703,
         n98704, n98705, n98706, n98707, n98708, n98709, n98710, n98711,
         n98712, n98713, n98714, n98715, n98716, n98717, n98718, n98719,
         n98720, n98721, n98722, n98723, n98724, n98725, n98726, n98727,
         n98728, n98729, n98730, n98731, n98732, n98733, n98734, n98735,
         n98736, n98737, n98738, n98739, n98740, n98741, n98742, n98743,
         n98744, n98745, n98746, n98747, n98748, n98749, n98750, n98751,
         n98752, n98753, n98754, n98755, n98756, n98757, n98758, n98759,
         n98760, n98761, n98762, n98763, n98764, n98765, n98766, n98767,
         n98768, n98769, n98770, n98771, n98772, n98773, n98774, n98775,
         n98776, n98777, n98778, n98779, n98780, n98781, n98782, n98783,
         n98784, n98785, n98786, n98787, n98788, n98789, n98790, n98791,
         n98792, n98793, n98794, n98795, n98796, n98797, n98798, n98799,
         n98800, n98801, n98802, n98803, n98804, n98805, n98806, n98807,
         n98808, n98809, n98810, n98811, n98812, n98813, n98814, n98815,
         n98816, n98817, n98818, n98819, n98820, n98821, n98822, n98823,
         n98824, n98825, n98826, n98827, n98828, n98829, n98830, n98831,
         n98832, n98833, n98834, n98835, n98836, n98837, n98838, n98839,
         n98840, n98841, n98842, n98843, n98844, n98845, n98846, n98847,
         n98848, n98849, n98850, n98851, n98852, n98853, n98854, n98855,
         n98856, n98857, n98858, n98859, n98860, n98861, n98862, n98863,
         n98864, n98865, n98866, n98867, n98868, n98869, n98870, n98871,
         n98872, n98873, n98874, n98875, n98876, n98877, n98878, n98879,
         n98880, n98881, n98882, n98883, n98884, n98885, n98886, n98887,
         n98888, n98889, n98890, n98891, n98892, n98893, n98894, n98895,
         n98896, n98897, n98898, n98899, n98900, n98901, n98902, n98903,
         n98904, n98905, n98906, n98907, n98908, n98909, n98910, n98911,
         n98912, n98913, n98914, n98915, n98916, n98917, n98918, n98919,
         n98920, n98921, n98922, n98923, n98924, n98925, n98926, n98927,
         n98928, n98929, n98930, n98931, n98932, n98933, n98934, n98935,
         n98936, n98937, n98938, n98940, n98941, n98942, n98943, n98944,
         n98946, n98947, n98948, n98949, n98950, n98951, n98952, n98953,
         n98954, n98955, n98956, n98957, n98958, n98959, n98960, n98961,
         n98962, n98963, n98964, n98965, n98966, n98967, n98968, n98969,
         n98970, n98971, n98972, n98973, n98974, n98975, n98976, n98977,
         n98978, n98979, n98980, n98981, n98982, n98983, n98984, n98985,
         n98986, n98987, n98988, n98989, n98990, n98991, n98992, n98993,
         n98994, n98995, n98996, n98997, n98998, n98999, n99000, n99001,
         n99002, n99003, n99004, n99005, n99006, n99007, n99008, n99009,
         n99010, n99011, n99012, n99013, n99014, n99015, n99016, n99017,
         n99018, n99019, n99020, n99021, n99022, n99023, n99024, n99025,
         n99026, n99027, n99028, n99029, n99030, n99031, n99032, n99033,
         n99034, n99035, n99036, n99037, n99038, n99039, n99040, n99041,
         n99042, n99043, n99044, n99045, n99046, n99047, n99048, n99049,
         n99050, n99051, n99052, n99053, n99054, n99055, n99056, n99057,
         n99058, n99059, n99060, n99061, n99062, n99063, n99064, n99065,
         n99066, n99067, n99068, n99069, n99070, n99071, n99072, n99073,
         n99074, n99075, n99076, n99077, n99078, n99079, n99080, n99081,
         n99082, n99083, n99084, n99085, n99086, n99087, n99088, n99089,
         n99090, n99091, n99092, n99093, n99094, n99095, n99096, n99097,
         n99098, n99099, n99100, n99101, n99102, n99103, n99104, n99105,
         n99106, n99107, n99108, n99109, n99110, n99111, n99112, n99113,
         n99114, n99115, n99116, n99117, n99118, n99119, n99120, n99121,
         n99122, n99123, n99124, n99125, n99126, n99127, n99128, n99129,
         n99130, n99131, n99132, n99133, n99134, n99135, n99136, n99137,
         n99138, n99139, n99140, n99141, n99142, n99143, n99144, n99145,
         n99146, n99147, n99148, n99149, n99150, n99151, n99152, n99153,
         n99154, n99155, n99156, n99157, n99158, n99159, n99160, n99161,
         n99162, n99163, n99164, n99165, n99166, n99167, n99168, n99169,
         n99170, n99171, n99172, n99173, n99174, n99175, n99176, n99177,
         n99178, n99179, n99180, n99181, n99182, n99183, n99184, n99185,
         n99186, n99187, n99188, n99189, n99190, n99191, n99192, n99193,
         n99194, n99195, n99196, n99197, n99198, n99199, n99200, n99201,
         n99202, n99203, n99204, n99205, n99206, n99207, n99208, n99209,
         n99210, n99211, n99212, n99213, n99214, n99215, n99216, n99217,
         n99218, n99219, n99220, n99221, n99222, n99223, n99224, n99225,
         n99226, n99227, n99228, n99229, n99230, n99231, n99232, n99233,
         n99234, n99235, n99236, n99237, n99238, n99239, n99240, n99241,
         n99242, n99243, n99244, n99245, n99246, n99247, n99248, n99249,
         n99250, n99251, n99252, n99253, n99254, n99255, n99256, n99257,
         n99258, n99259, n99260, n99261, n99262, n99263, n99264, n99265,
         n99266, n99267, n99268, n99269, n99270, n99271, n99272, n99273,
         n99274, n99275, n99276, n99277, n99278, n99279, n99280, n99281,
         n99282, n99283, n99284, n99285, n99286, n99287, n99288, n99289,
         n99290, n99291, n99292, n99293, n99294, n99295, n99296, n99297,
         n99298, n99299, n99300, n99301, n99302, n99303, n99304, n99305,
         n99306, n99307, n99308, n99309, n99310, n99311, n99312, n99313,
         n99314, n99315, n99316, n99317, n99318, n99319, n99320, n99321,
         n99322, n99323, n99324, n99325, n99326, n99327, n99328, n99329,
         n99330, n99331, n99332, n99333, n99334, n99335, n99336, n99337,
         n99338, n99339, n99340, n99341, n99342, n99343, n99344, n99345,
         n99346, n99347, n99348, n99349, n99350, n99351, n99352, n99353,
         n99354, n99355, n99356, n99357, n99358, n99359, n99360, n99361,
         n99362, n99363, n99364, n99365, n99366, n99367, n99368, n99369,
         n99370, n99371, n99372, n99373, n99374, n99375, n99376, n99377,
         n99378, n99379, n99380, n99381, n99382, n99383, n99384, n99385,
         n99386, n99387, n99388, n99389, n99390, n99391, n99392, n99393,
         n99394, n99395, n99396, n99397, n99398, n99399, n99400, n99401,
         n99402, n99403, n99404, n99405, n99406, n99407, n99408, n99409,
         n99410, n99411, n99412, n99413, n99414, n99415, n99416, n99417,
         n99418, n99419, n99420, n99421, n99422, n99423, n99424, n99425,
         n99426, n99427, n99428, n99429, n99430, n99431, n99432, n99433,
         n99434, n99435, n99436, n99437, n99438, n99439, n99440, n99441,
         n99442, n99443, n99444, n99445, n99446, n99447, n99448, n99449,
         n99450, n99451, n99452, n99453, n99454, n99455, n99456, n99457,
         n99458, n99459, n99460, n99461, n99462, n99463, n99464, n99465,
         n99466, n99467, n99468, n99469, n99470, n99471, n99472, n99473,
         n99474, n99475, n99476, n99477, n99478, n99479, n99480, n99481,
         n99482, n99483, n99484, n99485, n99486, n99487, n99488, n99489,
         n99490, n99491, n99492, n99493, n99494, n99495, n99496, n99497,
         n99498, n99499, n99500, n99501, n99502, n99503, n99504, n99505,
         n99506, n99507, n99508, n99509, n99510, n99511, n99512, n99513,
         n99514, n99515, n99516, n99517, n99518, n99519, n99520, n99521,
         n99522, n99523, n99524, n99525, n99526, n99527, n99528, n99529,
         n99530, n99531, n99532, n99533, n99534, n99535, n99536, n99537,
         n99538, n99539, n99540, n99541, n99542, n99543, n99544, n99545,
         n99546, n99547, n99548, n99549, n99550, n99551, n99552, n99553,
         n99554, n99555, n99556, n99557, n99558, n99559, n99560, n99561,
         n99562, n99563, n99564, n99565, n99566, n99567, n99568, n99569,
         n99570, n99571, n99572, n99573, n99574, n99575, n99576, n99577,
         n99578, n99579, n99580, n99581, n99582, n99583, n99584, n99585,
         n99586, n99587, n99588, n99589, n99590, n99591, n99592, n99593,
         n99594, n99595, n99596, n99597, n99598, n99599, n99600, n99601,
         n99602, n99603, n99604, n99605, n99606, n99607, n99608, n99609,
         n99610, n99611, n99612, n99613, n99614, n99615, n99616, n99617,
         n99618, n99619, n99620, n99621, n99622, n99623, n99624, n99625,
         n99626, n99627, n99628, n99629, n99630, n99631, n99632, n99633,
         n99634, n99635, n99636, n99637, n99638, n99639, n99640, n99641,
         n99642, n99643, n99644, n99645, n99646, n99647, n99648, n99649,
         n99650, n99651, n99652, n99653, n99654, n99655, n99656, n99657,
         n99658, n99659, n99660, n99661, n99662, n99663, n99664, n99665,
         n99666, n99667, n99668, n99669, n99670, n99671, n99672, n99673,
         n99674, n99675, n99676, n99677, n99678, n99679, n99680, n99681,
         n99682, n99683, n99684, n99685, n99686, n99687, n99688, n99689,
         n99690, n99691, n99692, n99693, n99694, n99695, n99696, n99697,
         n99698, n99699, n99700, n99701, n99702, n99703, n99704, n99705,
         n99706, n99707, n99708, n99709, n99710, n99711, n99712, n99713,
         n99714, n99715, n99716, n99717, n99718, n99719, n99720, n99721,
         n99722, n99723, n99724, n99725, n99726, n99727, n99728, n99729,
         n99730, n99731, n99732, n99733, n99734, n99735, n99736, n99737,
         n99738, n99739, n99740, n99741, n99742, n99743, n99744, n99745,
         n99746, n99747, n99748, n99749, n99750, n99751, n99752, n99753,
         n99754, n99755, n99756, n99757, n99758, n99759, n99760, n99761,
         n99762, n99763, n99764, n99765, n99766, n99767, n99768, n99769,
         n99770, n99771, n99772, n99773, n99774, n99775, n99776, n99777,
         n99778, n99779, n99780, n99781, n99782, n99783, n99784, n99785,
         n99786, n99787, n99788, n99789, n99790, n99791, n99792, n99793,
         n99794, n99795, n99796, n99797, n99798, n99799, n99800, n99801,
         n99802, n99803, n99804, n99805, n99806, n99807, n99808, n99809,
         n99810, n99811, n99812, n99813, n99814, n99815, n99816, n99817,
         n99818, n99819, n99820, n99821, n99822, n99823, n99824, n99825,
         n99826, n99827, n99828, n99829, n99830, n99831, n99832, n99833,
         n99834, n99835, n99836, n99837, n99838, n99839, n99840, n99841,
         n99842, n99843, n99844, n99845, n99846, n99847, n99848, n99849,
         n99850, n99851, n99852, n99853, n99854, n99855, n99856, n99857,
         n99858, n99859, n99860, n99861, n99862, n99863, n99864, n99865,
         n99866, n99867, n99868, n99869, n99870, n99871, n99872, n99873,
         n99874, n99875, n99876, n99877, n99878, n99879, n99880, n99881,
         n99882, n99883, n99884, n99885, n99886, n99887, n99888, n99889,
         n99890, n99891, n99892, n99893, n99894, n99895, n99896, n99897,
         n99898, n99899, n99900, n99901, n99902, n99903, n99904, n99905,
         n99906, n99907, n99908, n99909, n99910, n99911, n99912, n99913,
         n99914, n99915, n99916, n99917, n99918, n99919, n99920, n99921,
         n99922, n99923, n99924, n99925, n99926, n99927, n99928, n99929,
         n99930, n99931, n99932, n99933, n99934, n99935, n99936, n99937,
         n99938, n99939, n99940, n99941, n99942, n99943, n99944, n99945,
         n99946, n99947, n99948, n99949, n99950, n99951, n99952, n99953,
         n99954, n99955, n99956, n99957, n99958, n99959, n99960, n99961,
         n99962, n99963, n99964, n99965, n99966, n99967, n99968, n99969,
         n99970, n99971, n99972, n99973, n99974, n99975, n99976, n99977,
         n99978, n99979, n99980, n99981, n99982, n99983, n99984, n99985,
         n99986, n99987, n99988, n99989, n99990, n99991, n99992, n99993,
         n99994, n99995, n99996, n99997, n99998, n99999, n100000, n100001,
         n100002, n100003, n100004, n100005, n100006, n100007, n100008,
         n100009, n100010, n100011, n100012, n100013, n100014, n100015,
         n100016, n100017, n100018, n100019, n100020, n100021, n100022,
         n100023, n100024, n100025, n100026, n100027, n100028, n100029,
         n100030, n100031, n100032, n100033, n100034, n100035, n100036,
         n100037, n100038, n100039, n100040, n100041, n100042, n100043,
         n100044, n100045, n100046, n100047, n100048, n100049, n100050,
         n100051, n100052, n100053, n100054, n100055, n100056, n100057,
         n100058, n100059, n100060, n100061, n100062, n100063, n100064,
         n100065, n100066, n100067, n100068, n100069, n100070, n100071,
         n100072, n100073, n100074, n100075, n100076, n100077, n100078,
         n100079, n100080, n100081, n100082, n100083, n100084, n100085,
         n100086, n100089, n100090, n100091, n100092, n100093, n100094,
         n100095, n100096, n100097, n100098, n100099, n100100, n100101,
         n100102, n100103, n100104, n100105, n100106, n100107, n100108,
         n100109, n100110, n100111, n100112, n100113, n100114, n100115,
         n100116, n100117, n100118, n100119, n100120, n100121, n100122,
         n100123, n100124, n100125, n100126, n100127, n100128, n100129,
         n100130, n100131, n100132, n100133, n100134, n100135, n100136,
         n100137, n100138, n100139, n100140, n100141, n100142, n100144,
         n100145, n100146, n100147, n100148, n100149, n100150, n100151,
         n100153, n100154, n100156, n100157, n100158, n100159, n100160,
         n100161, n100162, n100163, n100164, n100165, n100166, n100167,
         n100168, n100169, n100170, n100171, n100172, n100173, n100174,
         n100175, n100176, n100177, n100178, n100179, n100180, n100181,
         n100182, n100183, n100184, n100185, n100186, n100187, n100188,
         n100189, n100190, n100191, n100192, n100193, n100194, n100195,
         n100196, n100197, n100198, n100199, n100200, n100201, n100202,
         n100203, n100204, n100205, n100206, n100207, n100208, n100209,
         n100210, n100211, n100212, n100213, n100214, n100215, n100216,
         n100217, n100218, n100219, n100220, n100221, n100222, n100223,
         n100224, n100225, n100228, n100229, n100230, n100231, n100232,
         n100233, n100234, n100235, n100236, n100237, n100238, n100239,
         n100240, n100241, n100242, n100243, n100244, n100245, n100246,
         n100247, n100248, n100249, n100250, n100251, n100252, n100253,
         n100254, n100255, n100256, n100257, n100258, n100259, n100260,
         n100261, n100262, n100263, n100264, n100265, n100266, n100268,
         n100269, n100270, n100271, n100272, n100273, n100274, n100275,
         n100276, n100277, n100278, n100280, n100281, n100282, n100283,
         n100284, n100285, n100286, n100287, n100288, n100289, n100290,
         n100291, n100292, n100295, n100296, n100297, n100298, n100300,
         n100301, n100302, n100303, n100304, n100305, n100306, n100307,
         n100308, n100309, n100310, n100311, n100312, n100313, n100314,
         n100315, n100316, n100317, n100318, n100319, n100320, n100321,
         n100322, n100323, n100324, n100325, n100326, n100327, n100328,
         n100329, n100330, n100331, n100332, n100333, n100334, n100335,
         n100336, n100337, n100338, n100339, n100340, n100341, n100342,
         n100343, n100344, n100345, n100346, n100347, n100348, n100349,
         n100350, n100351, n100352, n100353, n100354, n100355, n100356,
         n100357, n100358, n100359, n100361, n100362, n100363, n100365,
         n100366, n100367, n100368, n100369, n100370, n100371, n100372,
         n100373, n100374, n100375, n100376, n100377, n100378, n100379,
         n100380, n100381, n100382, n100383, n100384, n100385, n100386,
         n100387, n100388, n100389, n100390, n100391, n100392, n100393,
         n100394, n100395, n100396, n100397, n100398, n100399, n100400,
         n100401, n100402, n100403, n100404, n100405, n100406, n100407,
         n100408, n100409, n100410, n100411, n100412, n100413, n100414,
         n100415, n100416, n100417, n100418, n100419, n100420, n100422,
         n100423, n100424, n100426, n100427, n100428, n100429, n100430,
         n100460, n100462, n100463, n100496, n100561, n100562, n100563,
         n100564, n100565, n100566, n100567, n100568, n100569, n100570,
         n100571, n100572, n100573, n100574, n100575, n100576, n100577,
         n100578, n100579, n100580, n100581, n100582, n100583, n100584,
         n100585, n100586, n100587, n100588, n100589, n100590, n100591,
         n100592, n100593, n100594, n100595, n100596, n100597, n100598,
         n100599, n100600, n100601, n100602, n100603, n100604, n100605,
         n100606, n100607, n100608, n100609, n100610, n100611, n100612,
         n100613, n100614, n100615, n100616, n100617, n100618, n100619,
         n100620, n100621, n100622, n100623, n100624, n100629, n100630,
         n100631, n100632, n100633, n100634, n100635, n100636, n100637,
         n100638, n100639, n100640, n100641, n100642, n100643, n100644,
         n100645, n100646, n100647, n100648, n100649, n100651, n100653,
         n100655, n100657, n100659, n100661, n100663, n100665, n100667,
         n100669, n100671, n100673, n100675, n100677, n100679, n100681,
         n100683, n100685, n100687, n100689, n100691, n100693, n100695,
         n100697, n100699, n100701, n100703, n100705, n100707, n100709,
         n100711, n100717, n100718, n100719, n100762, n100767, n100770,
         n100771, n100775, n100779, n100784, n100794, n100795, n100796,
         n100799, n100800, n100801, n100892, n100893, n100894, n100992,
         n100993, n100994, n100997, n100998, n100999, n101000, n101001,
         n101002, n101003, n101004, n101005, n101006, n101007, n101008,
         n101009, n101010, n101012, n101013, n101014, n101015, n101016,
         n101017, n101018, n101019, n101020, n101021, n101022, n101023,
         n101024, n101025, n101026, n101027, n101028, n101029, n101030,
         n101031, n101032, n101033, n101034, n101035, n101036, n101037,
         n101038, n101039, n101040, n101041, n101042, n101043, n101044,
         n101045, n101046, n101047, n101048, n101049, n101050, n101051,
         n101052, n101054, n101055, n101056, n101057, n101058, n101059,
         n101060, n101061, n101062, n101063, n101064, n101065, n101066,
         n101067, n101148, n101149, n101150, n101151, n101152, n101153,
         n101154, n101155, n101156, n101157, n101158, n101159, n101160,
         n101161, n101162, n101163, n101164, n101165, n101166, n101167,
         n101168, n101169, n101170, n101171, n101172, n101173, n101174,
         n101175, n101176, n101177, n101178, n101179, n101624, n101661,
         n101665, n101666, n101679, n101683, n101684, n101697, n101701,
         n101702, n101715, n101719, n101720, n101733, n101737, n101738,
         n101751, n101755, n101756, n101769, n101771, n101772, n101785,
         n101789, n101790, n101803, n101805, n101806, n101819, n101823,
         n101824, n101837, n101841, n101842, n101855, n101857, n101858,
         n101871, n101875, n101876, n101889, n101891, n101892, n101905,
         n101907, n101908, n101921, n101923, n101924, n101937, n101939,
         n101940, n101953, n101955, n101956, n101969, n101971, n101972,
         n101985, n101987, n101988, n102001, n102005, n102006, n102019,
         n102023, n102024, n102036, n102040, n102041, n102052, n102056,
         n102057, n102070, n102074, n102075, n102087, n102091, n102092,
         n102101, n102105, n102106, n102115, n102119, n102120, n102131,
         n102133, n102134, n102145, n102149, n102150, n102160, n102164,
         n102165, n102174, n102178, n102179, n102188, n102190, n102197,
         n102199, n102208, n102210, n102217, n102219, n102228, n102230,
         n102237, n102239, n102247, n102249, n102256, n102258, n102267,
         n102269, n102276, n102278, n102286, n102288, n102295, n102297,
         n102306, n102308, n102315, n102317, n102318, n102326, n102328,
         n102335, n102337, n102346, n102348, n102355, n102357, n102366,
         n102373, n102375, n102384, n102386, n102393, n102395, n102404,
         n102406, n102413, n102415, n102424, n102426, n102433, n102435,
         n102444, n102451, n102453, n102462, n102464, n102471, n102473,
         n102482, n102489, n102491, n102500, n102507, n102509, n102518,
         n102520, n102526, n102528, n102537, n102543, n102545, n102554,
         n102560, n102562, n102570, n102576, n102578, n102585, n102591,
         n102593, n102600, n102606, n102608, n102614, n102620, n102622,
         n102630, n102637, n102639, n102646, n102653, n102655, n102663,
         n102665, n102672, n102673, n102679, n102686, n102688, n102694,
         n102700, n102702, n102708, n102710, n102716, n102718, n102725,
         n102727, n102733, n102734, n102739, n102741, n102745, n102747,
         n102752, n102754, n102756, n102759, n102763, n102766, n102767,
         n102772, n102774, n102776, n102779, n102783, n102786, n102787,
         n102792, n102794, n102796, n102799, n102803, n102806, n102807,
         n102812, n102814, n102816, n102819, n102823, n102826, n102827,
         n102832, n102834, n102836, n102839, n102843, n102846, n102847,
         n102852, n102854, n102856, n102859, n102863, n102866, n102867,
         n102872, n102874, n102876, n102879, n102883, n102886, n102887,
         n102892, n102894, n102896, n102899, n102903, n102906, n102907,
         n102912, n102914, n102916, n102919, n102923, n102926, n102927,
         n102932, n102934, n102936, n102939, n102943, n102946, n102947,
         n102952, n102954, n102956, n102959, n102963, n102966, n102967,
         n102971, n102973, n102975, n102980, n102983, n102984, n102989,
         n102991, n102993, n102996, n103000, n103003, n103004, n103009,
         n103011, n103013, n103016, n103020, n103023, n103024, n103029,
         n103031, n103033, n103036, n103040, n103043, n103044, n103049,
         n103051, n103053, n103056, n103060, n103063, n103064, n103069,
         n103071, n103073, n103076, n103080, n103083, n103084, n103089,
         n103091, n103093, n103096, n103100, n103103, n103104, n103109,
         n103111, n103113, n103116, n103120, n103123, n103124, n103129,
         n103131, n103133, n103138, n103141, n103142, n103147, n103149,
         n103151, n103154, n103158, n103161, n103162, n103167, n103169,
         n103171, n103173, n103177, n103180, n103181, n103186, n103188,
         n103190, n103192, n103196, n103199, n103200, n103205, n103207,
         n103209, n103211, n103214, n103217, n103218, n103223, n103225,
         n103227, n103229, n103233, n103236, n103237, n103242, n103244,
         n103246, n103248, n103252, n103255, n103256, n103261, n103263,
         n103265, n103267, n103271, n103274, n103275, n103280, n103282,
         n103284, n103286, n103290, n103293, n103294, n103301, n103303,
         n103307, n103310, n103311, n103316, n103318, n103320, n103326,
         n103327, n103332, n103337, n103338, n103342, n103344, n103350,
         n103351, n103354, n103358, n103367, n103369, n103374, n103378,
         n103387, n103389, n103394, n103398, n103407, n103409, n103414,
         n103418, n103427, n103429, n103434, n103438, n103447, n103449,
         n103454, n103458, n103467, n103469, n103473, n103477, n103486,
         n103488, n103492, n103496, n103505, n103507, n103511, n103515,
         n103524, n103526, n103530, n103533, n103542, n103544, n103548,
         n103552, n103559, n103562, n103566, n103569, n103578, n103579,
         n103583, n103587, n103595, n103597, n103601, n103605, n103614,
         n103616, n103620, n103624, n103632, n103634, n103638, n103642,
         n103650, n103651, n103655, n103659, n103667, n103669, n103673,
         n103677, n103685, n103687, n103691, n103695, n103703, n103704,
         n103708, n103712, n103720, n103721, n103726, n103729, n103736,
         n103737, n103742, n103746, n103753, n103754, n103759, n103763,
         n103770, n103771, n103776, n103780, n103787, n103788, n103793,
         n103796, n103804, n103805, n103812, n103820, n103821, n103829,
         n103835, n103837, n103843, n103850, n103851, n103855, n103860,
         n103867, n103869, n103874, n103878, n103885, n103886, n103890,
         n103893, n103900, n103901, n103911, n103912, n103915, n103916,
         n103917, n103918, n103919, n103920, n103921, n103922, n103923,
         n103924, n103925, n103926, n103927, n103928, n103929, n103930,
         n103931, n103932, n103933, n103934, n103935, n103936, n103937,
         n103938, n103939, n103940, n103942, n103943, n103944, n103945,
         n103946, n103947, n103948, n103949, n103950, n103951, n103952,
         n103953, n103954, n103955, n103956, n103957, n103958, n103959,
         n103960, n103961, n103962, n103963, n103964, n103965, n103966,
         n103967, n103968, n103969, n103970, n103971, n103972, n103973,
         n103974, n103975, n103976, n103977, n103978, n103979, n103980,
         n103981, n103982, n103983, n103984, n103985, n103986, n103987,
         n103988, n103989, n103990, n103991, n103992, n103993, n103994,
         n103995, n103996, n103997, n103998, n103999, n104000, n104001,
         n104002, n104003, n104004, n104005, n104006, n104007, n104008,
         n104009, n104010, n104011, n104012, n104013, n104014, n104015,
         n104016, n104017, n104018, n104019, n104020, n104021, n104022,
         n104023, n104024, n104025, n104026, n104027, n104028, n104029,
         n104030, n104031, n104032, n104033, n104034, n104035, n104036,
         n104037, n104038, n104039, n104040, n104041, n104042, n104043,
         n104044, n104045, n104046, n104047, n104048, n104049, n104050,
         n104051, n104052, n104053, n104054, n104055, n104056, n104057,
         n104058, n104059, n104060, n104061, n104062, n104063, n104064,
         n104065, n104066, n104067, n104068, n104069, n104070, n104071,
         n104072, n104073, n104074, n104075, n104076, n104077, n104078,
         n104079, n104080, n104081, n104082, n104083, n104084, n104085,
         n104086, n104087, n104088, n104089, n104090, n104091, n104092,
         n104093, n104094, n104095, n104096, n104097, n104098, n104099,
         n104100, n104101, n104102, n104103, n104104, n104105, n104106,
         n104107, n104108, n104109, n104110, n104111, n104112, n104113,
         n104114, n104115, n104116, n104117, n104118, n104119, n104120,
         n104121, n104122, n104123, n104124, n104125, n104126, n104127,
         n104128, n104129, n104130, n104131, n104132, n104133, n104134,
         n104135, n104136, n104137, n104138, n104139, n104140, n104141,
         n104142, n104143, n104144, n104145, n104146, n104147, n104148,
         n104149, n104150, n104151, n104152, n104153, n104154, n104155,
         n104156, n104157, n104158, n104159, n104160, n104161, n104162,
         n104163, n104164, n104165, n104166, n104167, n104168, n104169,
         n104170, n104171, n104172, n104173, n104174, n104175, n104176,
         n104177, n104178, n104179, n104180, n104181, n104182, n104183,
         n104184, n104185, n104186, n104187, n104188, n104189, n104190,
         n104191, n104192, n104193, n104194, n104195, n104196, n104197,
         n104198, n104199, n104200, n104201, n104202, n104203, n104204,
         n104205, n104206, n104207, n104208, n104209, n104210, n104211,
         n104212, n104213, n104214, n104215, n104216, n104217, n104218,
         n104219, n104220, n104221, n104222, n104223, n104224, n104225,
         n104226, n104227, n104228, n104229, n104230, n104231, n104232,
         n104233, n104234, n104235, n104236, n104237, n104238, n104239,
         n104240, n104241, n104242, n104243, n104244, n104245, n104246,
         n104247, n104248, n104249, n104250, n104251, n104252, n104253,
         n104254, n104255, n104256, n104257, n104258, n104259, n104260,
         n104261, n104262, n104263, n104264, n104265, n104266, n104267,
         n104268, n104269, n104270, n104271, n104272, n104273, n104274,
         n104275, n104276, n104277, n104278, n104279, n104280, n104281,
         n104282, n104283, n104284, n104285, n104286, n104287, n104288,
         n104289, n104290, n104291, n104292, n104293, n104294, n104295,
         n104296, n104297, n104298, n104299, n104300, n104301, n104302,
         n104303, n104304, n104305, n104306, n104307, n104308, n104309,
         n104310, n104311, n104312, n104313, n104314, n104315, n104316,
         n104317, n104320, n104321, n104322, n104323, n104324, n104325,
         n104326, n104327, n104328, n104329, n104330, n104331, n104332,
         n104333, n104334, n104335, n104336, n104337, n104338, n104339,
         n104340, n104341, n104342, n104343, n104344, n104345, n104346,
         n104347, n104348, n104349, n104350, n104351, n104352, n104353,
         n104354, n104355, n104356, n104357, n104358, n104359, n104360,
         n104361, n104362, n104363, n104364, n104365, n104366, n104367,
         n104368, n104369, n104370, n104371, n104372, n104373, n104374,
         n104375, n104376, net67007, net67008, net68722, net68723, net71745,
         net73629, net82027, net112354, net112358, net112383, net112469,
         net112601, net113159, net113157, net113156, net113155, net113154,
         net113153, net113152, net113102, net113091, net113081, net113538,
         n82424, n82423, n82422, n82091, n104377, n104378, n104379, n104380,
         n104381, n104382, n104383, n104384, n104385, n104386, n104387,
         n104388, n104389, n104390, n104391, n104392, n104393, n104394,
         n104395, n104396, n104397, n104398, n104399, n104400, n104401,
         n104402, n104403, n104404, n104405, n104406, n104407, n104408,
         n104409, n104410, n104411, n104412, n104413, n104414, n104415,
         n104416, n104417, n104418, n104419, n104420, n104421, n104422,
         n104423, n104424, n104425, n104426, n104427, n104428, n104429,
         n104430, n104431, n104432, n104433, n104434, n104435, n104436,
         n104437, n104438, n104439, n104440, n104441, n104442, n104443,
         n104444, n104445, n104446, n104447, n104448, n104449, n104450,
         n104451, n104452, n104453, n104454, n104455, n104456, n104457,
         n104458, n104459, n104460, n104461, n104462, n104463, n104464,
         n104465, n104466, n104467, n104468, n104469, n104470, n104471,
         n104472, n104473, n104474, n104475, n104476, n104477, n104478,
         n104479, n104480, n104481, n104482, n104483, n104484, n104485,
         n104486, n104487, n104488, n104489, n104490, n104491, n104492,
         n104493, n104494, n104495, n104496, n104497, n104498, n104499,
         n104500, n104501, n104502, n104503, n104504, n104505, n104506,
         n104507, n104508, n104509, n104510, n104511, n104512, n104513,
         n104514, n104515, n104516, n104517, n104518, n104519, n104520,
         n104521, n104522, n104523, n104524, n104525, n104526, n104527,
         n104528, n104529, n104530, n104531, n104532, n104533, n104534,
         n104535, n104536, n104537, n104538, n104539, n104540, n104541,
         n104542, n104543, n104544, n104545, n104546, n104547, n104548,
         n104549, n104550, n104551, n104552, n104553, n104554, n104555,
         n104556, n104557, n104558, n104559, n104560, n104561, n104562,
         n104563, n104564, n104565, n104566, n104567, n104568, n104569,
         n104570, n104571, n104572, n104573, n104574, n104575, n104576,
         n104577, n104578, n104579, n104580, n104581, n104582, n104583,
         n104584, n104585, n104586, n104587, n104588, n104589, n104590,
         n104591, n104592, n104593, n104594, n104595, n104596, n104597,
         n104598, n104599, n104600, n104601, n104602, n104603, n104604,
         n104605, n104606, n104607, n104608, n104609, n104610, n104611,
         n104612, n104613, n104614, n104615, n104616, n104617, n104618,
         n104619, n104620, n104621, n104622, n104623, n104624, n104625,
         n104626, n104627, n104628, n104629, n104630, n104631, n104632,
         n104633, n104634, n104635, n104636, n104637, n104638, n104639,
         n104640, n104641, n104642, n104643, n104644, n104645, n104646,
         n104647, n104648, n104649, n104650, n104651, n104652, n104653,
         n104654, n104655, n104656, n104657, n104658, n104659, n104660,
         n104661, n104662, n104663, n104664, n104665, n104666, n104667,
         n104668, n104669, n104670, n104671, n104687, n104688, n104689,
         n104690, n104691, n104692, n104693, n104694, n104695, n104696,
         n104697, n104698, n104699, n104700, n104701, n104702, n104703,
         n104704, n104705, n104706, n104707, n104708, n104709, n104710,
         n104711, n104712, n104713, n104714, n104715, n104716, n104717,
         n104718, n104719, n104720, n104721, n104722, n104723, n104724,
         n104725, n104726, n104727, n104728, n104729, n104730, n104731,
         n104732, n104733, n104734, n104735, n104736, n104737, n104738,
         n104739, n104740, n104741, n104743, n104744, n104745, n104746,
         n104747, n104748, n104749, n104750, n104751, n104752, n104753,
         n104754, n104755, n104756, n104757, n104758, n104759, n104760,
         n104761, n104762, n104763, n104764, n104765, n104766, n104767,
         n104768, n104769, n104770, n104771, n104772, n104773, n104774,
         n104775, n104776, n104777, n104778, n104779, n104780, n104781,
         n104782, n104783, n104784, n104785, n104786, n104787, n104788,
         n104789, n104790, n104791, n104792, n104793, n104794, n104795,
         n104796, n104797, n104798, n104799, n104800, n104801, n104802,
         n104803, n104804, n104805, n104806, n104807, n104808, n104809,
         n104810, n104811, n104812, n104813, n104814, n104815, n104816,
         n104817, n104818, n104819, n104820, n104821, n104822, n104823,
         n104824, n104825, n104826, n104827, n104828, n104829, n104830,
         n104831, n104832, n104833, n104835, n104836, n104837, n104838,
         n104839, n104840, n104841, n104842, n104843, n104844, n104845,
         n104846, n104847, n104848, n104849, n104850, n104851, n104852,
         n104853, n104854, n104855, n104856, n104857, n104858, n104859,
         n104860, n104861, n104862, n104863, n104864, n104865, n104866,
         n104867, n104868, n104869, n104870, n104871, n104872, n104873,
         n104874, n104875, n104876, n104877, n104878, n104879, n104880,
         n104881, n104882, n104883, n104884, n104885, n104886, n104887,
         n104888, n104889, n104890, n104891, n104892, n104893, n104894,
         n104895, n104896, n104897, n104898, n104899, n104900, n104901,
         n104902, n104903, n104904, n104905, n104906, n104907, n104908,
         n104909, n104910, n104911, n104912, n104913, n104914, n104915,
         n104916, n104917, n104918, n104919, n104920, n104921, n104922,
         n104923, n104924, n104925, n104926, n104927, n104928, n104929,
         n104930, n104931, n104932, n104933, n104934, n104935, n104936,
         n104937, n104938, n104939, n104940, n104941, n104942, n104943,
         n104944, n104945, n104946, n104947, n104948, n104949, n104950,
         n104951, n104952, n104953, n104954, n104955, n104956, n104957,
         n104958, n104959, n104960, n104961, n104962, n104963, n104964,
         n104965, n104966, n104967, n104968, n104969, n104970, n104971,
         n104972, n104973, n104974, n104975, n104976, n104977, n104978,
         n104979, n104980, n104981, n104982, n104983, n104984, n104985,
         n104986, n104987, n104988, n104989, n104990, n104991, n104992,
         n104993, n104994, n104995, n104996, n104997, n104998, n104999,
         n105000, n105001, n105002, n105003, n105004, n105005, n105006,
         n105007, n105008, n105009, n105010, n105011, n105012, n105013,
         n105014, n105015, n105016, n105017, n105018, n105019, n105020,
         n105021, n105022, n105023, n105024, n105025, n105026, n105027,
         n105028, n105029, n105030, n105031, n105032, n105033, n105034,
         n105035, n105036, n105037, n105038, n105039, n105040, n105041,
         n105042, n105043, n105044, n105045, n105046, n105047, n105048,
         n105049, n105050, n105051, n105052, n105053, n105054, n105055,
         n105056, n105057, n105058, n105059, n105060, n105061, n105062,
         n105063, n105064, n105065, n105066, n105067, n105068, n105069,
         n105071, n105072, n105073, n105074, n105075, n105076, n105077,
         n105078, n105079, n105080, n105081, n105082, n105083, n105085,
         n105086, n105087, n105088, n105089, n105090, n105091, n105092,
         n105093, n105094, n105095, n105096, n105097, n105098, n105099,
         n105100, n105101, n105102, n105103, n105104, n105105, n105106,
         n105107, n105108, n105109, n105110, n105111, n105112, n105113,
         n105114, n105115, n105116, n105117, n105118, n105119, n105120,
         n105121, n105122, n105123, n105124, n105125, n105126, n105127,
         n105128, n105129, n105130, n105131, n105132, n105133, n105134,
         n105135, n105136, n105137, n105138, n105139, n105140, n105141,
         n105142, n105143, n105144, n105145, n105146, n105147, n105148,
         n105149, n105150, n105151, n105152, n105153, n105154, n105155,
         n105156, n105157, n105158, n105159, n105160, n105161, n105162,
         n105163, n105164, n105165, n105166, n105167, n105168, n105169,
         n105170, n105171, n105172, n105173, n105174, n105175, n105176,
         n105177, n105178, n105179, n105180, n105181, n105182, n105183,
         n105184, n105185, n105186, n105187, n105188, n105189, n105190,
         n105191, n105192, n105193, n105194, n105195, n105196, n105197,
         n105198, n105199, n105200, n105201, n105202, n105203, n105204,
         n105205, n105206, n105207, n105208, n105209, n105210, n105211,
         n105212, n105213, n105214, n105215, n105216, n105217, n105218,
         n105219, n105220, n105221, n105222, n105223, n105224, n105225,
         n105226, n105227, n105228, n105229, n105230, n105231, n105232,
         n105233, n105234, n105235, n105236, n105237, n105238, n105239,
         n105240, n105241, n105242, n105243, n105244, n105245, n105246,
         n105247, n105248, n105249, n105250, n105251, n105252, n105253,
         n105254, n105255, n105256, n105257, n105258, n105259, n105260,
         n105261, n105262, n105263, n105264, n105265, n105266, n105267,
         n105268, n105269, n105270, n105271, n105272, n105273, n105274,
         n105275, n105276, n105277, n105278, n105279, n105280, n105281,
         n105282, n105283, n105284, n105285, n105286, n105287, n105288,
         n105289, n105290, n105291, n105292, n105293, n105294, n105295,
         n105296, n105297, n105298, n105299, n105300, n105301, n105302,
         n105303, n105304, n105305, n105306, n105307, n105308, n105309,
         n105310, n105311, n105312, n105313, n105314, n105315, n105316,
         n105317, n105318, n105319, n105320, n105321, n105322, n105323,
         n105324, n105325, n105326, n105327, n105328, n105329, n105330,
         n105331, n105332, n105333, n105334, n105335, n105336, n105337,
         n105338, n105339, n105340, n105341, n105342, n105343, n105344,
         n105345, n105346, n105347, n105348, n105349, n105350, n105351,
         n105352, n105353, n105354, n105355, n105356, n105357, n105358,
         n105359, n105360, n105361, n105362, n105363, n105364, n105365,
         n105366, n105367, n105368, n105369, n105370, n105371, n105372,
         n105373, n105374, n105375, n105376, n105377, n105378, n105379,
         n105380, n105381, n105382, n105383, n105384, n105385, n105386,
         n105387, n105388, n105389, n105390, n105391, n105392, n105393,
         n105394, n105395, n105396, n105397, n105398, n105399, n105400,
         n105401, n105402, n105403, n105404, n105405, n105406, n105407,
         n105408, n105409, n105410, n105411, n105412, n105413, n105414,
         n105415, n105416, n105417, n105418, n105419, n105420, n105421,
         n105422, n105423, n105424, n105425, n105426, n105427, n105428,
         n105429, n105430, n105431, n105432, n105433, n105434, n105435,
         n105436, n105437, n105438, n105439, n105440, n105441, n105442,
         n105443, n105444, n105445, n105446, n105447, n105448, n105449,
         n105450, n105451, n105452, n105453, n105454, n105455, n105456,
         n105457, n105458, n105459, n105460, n105461, n105462, n105463,
         n105464, n105465, n105466, n105467, n105468, n105469, n105470,
         n105471, n105472, n105473, n105474, n105475, n105476, n105477,
         n105478, n105479, n105480, n105481, n105482, n105483, n105484,
         n105485, n105486, n105487, n105488, n105489, n105490, n105491,
         n105492, n105493, n105494, n105495, n105496, n105497, n105498,
         n105499, n105500, n105501, n105502, n105503, n105504, n105505,
         n105506, n105507, n105508, n105509, n105510, n105511, n105512,
         n105513, n105514, n105515, n105516, n105517, n105518, n105519,
         n105520, n105521, n105522, n105523, n105524, n105525, n105526,
         n105527, n105528, n105529, n105530, n105531, n105532, n105533,
         n105534, n105535, n105536, n105537, n105538, n105539, n105540,
         n105541, n105542, n105543, n105544, n105545, n105546, n105547,
         n105548, n105549, n105550, n105551, n105552, n105553, n105554,
         n105555, n105556, n105557, n105558, n105559, n105560, n105561,
         n105562, n105563, n105564, n105565, n105566, n105567, n105568,
         n105569, n105570, n105571, n105572, n105573, n105574, n105575,
         n105576, n105577, n105578, n105579, n105580, n105581, n105582,
         n105583, n105584, n105585, n105586, n105587, n105588, n105589,
         n105590, n105591, n105592, n105593, n105594, n105595, n105596,
         n105597, n105598, n105599, n105600, n105601, n105602, n105603,
         n105604, n105605, n105606, n105607, n105608, n105609, n105610,
         n105611, n105612, n105613, n105614, n105615, n105616, n105617,
         n105618, n105619, n105620, n105621, n105622, n105623, n105624,
         n105625, n105626, n105627, n105628, n105629, n105630, n105631,
         n105632, n105633, n105634, n105635, n105636, n105637, n105638,
         n105639, n105640, n105641, n105642, n105643, n105644, n105645,
         n105646, n105647, n105648, n105649, n105650, n105651, n105652,
         n105653, n105654, n105655, n105656, n105657, n105658, n105659,
         n105660, n105661, n105662, n105663, n105664, n105665, n105666,
         n105667, n105668, n105669, n105670, n105671, n105672, n105673,
         n105674, n105675, n105676, n105677, n105678, n105679, n105680,
         n105681, n105682, n105683, n105684, n105685, n105686, n105687,
         n105688, n105689, n105690, n105691, n105692, n105693, n105694,
         n105695, n105696, n105697, n105698, n105699, n105700, n105701,
         n105702, n105703, n105704, n105705, n105706, n105707, n105708,
         n105709, n105710, n105711, n105712, n105713, n105714, n105715,
         n105716, n105717, n105718, n105719, n105720, n105721, n105722,
         n105723, n105724, n105725, n105726, n105727, n105728, n105729,
         n105730, n105731, n105732, n105733, n105734, n105735, n105736,
         n105737, n105738, n105739, n105740, n105741, n105742, n105743,
         n105744, n105745, n105746, n105747, n105748, n105749, n105750,
         n105751, n105752, n105753, n105754, n105755, n105756, n105757,
         n105758, n105759, n105760, n105761, n105762, n105763, n105764,
         n105765, n105766, n105767, n105768, n105769, n105770, n105771,
         n105772, n105773, n105774, n105775, n105776, n105777, n105778,
         n105779, n105780, n105781, n105782, n105783, n105784, n105785,
         n105786, n105787, n105788, n105789, n105790, n105791, n105792,
         n105793, n105794, n105795, n105796, n105797, n105798, n105799,
         n105800, n105801, n105802, n105803, n105804, n105805, n105806,
         n105807, n105808, n105809, n105810, n105811, n105812, n105813,
         n105814, n105815, n105816, n105817, n105818, n105819, n105820,
         n105821, n105822, n105823, n105824, n105825, n105826, n105827,
         n105828, n105829, n105830, n105831, n105832, n105833, n105834,
         n105835, n105836, n105837, n105838, n105839, n105840, n105841,
         n105842, n105843, n105844, n105845, n105846, n105847, n105848,
         n105849, n105850, n105851, n105852, n105853, n105854, n105855,
         n105856, n105857, n105858, n105859, n105860, n105861, n105862,
         n105863, n105864, n105865, n105866, n105867, n105868, n105869,
         n105870, n105871, n105872, n105873, n105874, n105875, n105876,
         n105877, n105878, n105879, n105880, n105881, n105882, n105883,
         n105884, n105885, n105886, n105887, n105888, n105889, n105890,
         n105891, n105892, n105893, n105894, n105895, n105896, n105897,
         n105898, n105899, n105900, n105901, n105902, n105903, n105904,
         n105905, n105906, n105907, n105908, n105909, n105910, n105911,
         n105912, n105913, n105914, n105915, n105916, n105917, n105918,
         n105919, n105920, n105921, n105922, n105923, n105924, n105925,
         n105926, n105927, n105928, n105929, n105930, n105931, n105932,
         n105933, n105934, n105935, n105936, n105937, n105938, n105939,
         n105940, n105941, n105942, n105943, n105944, n105945, n105946,
         n105947, n105948, n105949, n105950, n105951, n105952, n105953,
         n105954, n105955, n105956, n105957, n105958, n105959, n105960,
         n105961, n105962, n105963, n105964, n105965, n105966, n105967,
         n105968, n105969, n105970, n105971, n105972, n105973, n105974,
         n105975, n105976, n105977, n105978, n105979, n105980, n105981,
         n105982, n105983, n105984, n105985, n105986, n105987, n105988,
         n105989, n105990, n105991, n105992, n105993, n105994, n105995,
         n105996, n105997, n105998, n105999, n106000, n106001, n106002,
         n106003, n106004, n106005, n106006, n106007, n106008, n106009,
         n106010, n106011, n106012, n106013, n106014, n106015, n106016,
         n106017, n106018, n106019, n106020, n106021, n106022, n106023,
         n106024, n106025, n106026, n106027, n106028, n106029, n106030,
         n106031, n106032, n106033, n106034, n106035, n106036, n106037,
         n106038, n106039, n106040, n106041, n106042, n106043, n106044,
         n106045, n106046, n106047, n106048, n106049, n106050, n106051,
         n106052, n106053, n106054, n106055, n106056, n106057, n106058,
         n106059, n106060, n106061, n106062, n106063, n106064, n106065,
         n106066, n106067, n106068, n106069, n106070, n106071, n106072,
         n106073, n106074, n106075, n106076, n106077, n106078, n106079,
         n106080, n106081, n106082, n106083, n106084, n106085, n106086,
         n106087, n106088, n106089, n106090, n106091, n106092, n106093,
         n106094, n106095, n106096, n106097, n106098, n106099, n106100,
         n106101, n106102, n106103, n106104, n106105, n106106, n106107,
         n106108, n106109, n106110, n106111, n106112, n106113, n106114,
         n106115, n106116, n106117, n106118, n106119, n106120, n106121,
         n106122, n106123, n106124, n106125, n106126, n106127, n106128,
         n106129, n106130, n106131, n106132, n106133, n106134, n106135,
         n106136, n106137, n106138, n106139, n106140, n106141, n106142,
         n106143, n106144, n106145, n106146, n106147, n106148, n106149,
         n106150, n106151, n106152, n106153, n106154, n106155, n106156,
         n106157, n106158, n106159, n106160, n106161, n106162, n106163,
         n106164, n106165, n106166, n106167, n106168, n106169, n106170,
         n106171, n106172, n106173, n106174, n106175, n106176, n106177,
         n106178, n106179, n106180, n106181, n106182, n106183, n106184,
         n106185, n106186, n106187, n106188, n106189, n106190, n106191,
         n106192, n106193, n106194, n106195, n106196, n106197, n106198,
         n106199, n106200, n106201, n106202, n106203, n106204, n106205,
         n106206, n106207, n106208, n106209, n106210, n106211, n106212,
         n106213, n106214, n106215, n106216, n106217, n106218, n106219,
         n106220, n106221, n106222, n106223, n106224, n106225, n106226,
         n106227, n106228, n106229, n106230, n106231, n106232, n106233,
         n106234, n106235, n106236, n106237, n106238, n106239, n106240,
         n106241, n106242, n106243, n106244, n106245, n106246, n106247,
         n106248, n106249, n106250, n106251, n106252, n106253, n106254,
         n106255, n106256, n106257, n106258, n106259, n106260, n106261,
         n106262, n106263, n106264, n106265, n106266, n106267, n106268,
         n106269, n106270, n106271, n106272, n106273, n106274, n106275,
         n106276, n106277, n106278, n106279, n106280, n106281, n106282,
         n106283, n106284, n106285, n106286, n106287, n106288, n106289,
         n106290, n106291, n106292, n106293, n106294, n106295, n106296,
         n106297, n106298, n106299, n106300, n106301, n106302, n106303,
         n106304, n106305, n106306, n106307, n106308, n106309, n106310,
         n106311, n106312, n106313, n106314, n106315, n106316, n106317,
         n106318, n106319, n106320, n106321, n106322, n106323, n106324,
         n106325, n106326, n106327, n106328, n106329, n106330, n106331,
         n106332, n106333, n106334, n106335, n106336, n106337, n106338,
         n106339, n106340, n106341, n106342, n106343, n106344, n106345,
         n106346, n106347, n106348, n106349, n106350, n106351, n106352,
         n106353, n106354, n106355, n106356, n106357, n106358, n106359,
         n106360, n106361, n106362, n106363, n106364, n106365, n106366,
         n106367, n106368, n106369, n106370, n106371, n106372, n106373,
         n106374, n106375, n106376, n106377, n106378, n106379, n106380,
         n106381, n106382, n106383, n106384, n106385, n106386, n106387,
         n106388, n106389, n106390, n106391, n106392, n106393, n106394,
         n106395, n106396, n106397, n106398, n106399, n106400, n106401,
         n106402, n106403, n106404, n106405, n106406, n106407, n106408,
         n106409, n106410, n106411, n106412, n106413, n106414, n106415,
         n106416, n106417, n106418, n106419, n106420, n106421, n106422,
         n106423, n106424, n106425, n106426, n106427, n106428, n106429,
         n106430, n106431, n106432, n106433, n106434, n106435, n106436,
         n106437, n106438, n106439, n106440, n106441, n106442, n106443,
         n106444, n106445, n106446, n106447, n106448, n106449, n106450,
         n106451, n106452, n106453, n106454, n106455, n106456, n106457,
         n106458, n106459, n106460, n106461, n106462, n106463, n106464,
         n106465, n106466, n106467, n106468, n106469, n106470, n106471,
         n106472, n106473, n106474, n106475, n106476, n106477, n106478,
         n106479, n106480, n106481, n106482, n106483, n106484, n106485,
         n106486, n106487, n106488, n106489, n106490, n106491, n106492,
         n106493, n106494, n106495, n106496, n106497, n106498, n106499,
         n106500, n106501, n106502, n106503, n106504, n106505, n106506,
         n106507, n106508, n106509, n106510, n106511, n106512, n106513,
         n106514, n106515, n106516, n106517, n106518, n106519, n106520,
         n106521, n106522, n106523, n106524, n106525, n106526, n106527,
         n106528, n106529, n106530, n106531, n106532, n106533, n106534,
         n106535, n106536, n106537, n106538, n106539, n106540, n106541,
         n106542, n106543, n106544, n106545, n106546, n106547, n106548,
         n106549, n106550, n106551, n106552, n106553, n106554, n106555,
         n106556, n106557, n106558, n106559, n106560, n106561, n106562,
         n106563, n106564, n106565, n106566, n106567, n106568, n106569,
         n106570, n106571, n106572, n106573, n106574, n106575, n106576,
         n106577, n106578, n106579, n106580, n106581, n106582, n106583,
         n106584, n106585, n106586, n106587, n106588, n106589, n106590,
         n106591, n106592, n106593, n106594, n106595, n106596, n106597,
         n106598, n106599, n106600, n106601, n106602, n106603, n106604,
         n106605, n106606, n106607, n106608, n106609, n106610, n106611,
         n106612, n106613, n106614, n106615, n106616, n106617, n106618,
         n106619, n106620, n106621, n106622, n106623, n106624, n106625,
         n106626, n106627, n106628, n106629, n106630, n106631, n106632,
         n106633, n106634, n106635, n106636, n106637, n106638, n106639,
         n106640, n106641, n106642, n106643, n106644, n106645, n106646,
         n106647, n106648, n106649, n106650, n106651, n106652, n106653,
         n106654, n106655, n106656, n106657, n106658, n106659, n106660,
         n106661, n106662, n106663, n106664, n106665, n106666, n106667,
         n106668, n106669, n106670, n106671, n106672, n106673, n106674,
         n106675, n106676, n106677, n106678, n106679, n106680, n106681,
         n106682, n106683, n106684, n106685, n106686, n106687, n106688,
         n106689, n106690, n106691, n106692, n106693, n106694, n106695,
         n106696, n106697, n106698, n106699, n106700, n106701, n106702,
         n106703, n106704, n106705, n106706, n106707, n106708, n106709,
         n106710, n106711, n106712, n106713, n106714, n106715, n106716,
         n106717, n106718, n106719, n106720, n106721, n106722, n106723,
         n106724, n106725, n106726, n106727, n106728, n106729, n106730,
         n106731, n106732, n106733, n106734, n106735, n106736, n106737,
         n106738, n106739, n106740, n106741, n106742, n106743, n106744,
         n106745, n106746, n106747, n106748, n106749, n106750, n106751,
         n106752, n106753, n106754, n106755, n106756, n106757, n106758,
         n106759, n106760, n106761, n106762, n106763, n106764, n106765,
         n106766, n106767, n106768, n106769, n106770, n106771, n106772,
         n106773, n106774, n106775, n106776, n106777, n106778, n106779,
         n106780, n106781, n106782, n106783, n106784, n106785, n106786,
         n106787, n106788, n106789, n106790, n106791, n106792, n106793,
         n106794, n106795, n106796, n106797, n106798, n106799, n106800,
         n106801, n106802, n106803, n106804, n106805, n106806, n106807,
         n106808, n106809, n106810, n106811, n106812, n106813, n106814,
         n106815, n106816, n106817, n106818, n106819, n106820, n106821,
         n106822, n106823, n106824, n106825, n106826, n106827, n106828,
         n106829, n106830, n106831, n106832, n106833, n106834, n106835,
         n106836, n106837, n106838, n106839, n106840, n106841, n106842,
         n106843, n106844, n106845, n106846, n106847, n106848, n106849,
         n106850, n106851, n106852, n106853, n106854, n106855, n106856,
         n106857, n106858, n106859, n106860, n106861, n106862, n106863,
         n106864, n106865, n106866, n106867, n106868, n106869, n106870,
         n106871, n106872, n106873, n106874, n106875, n106876, n106877,
         n106878, n106879, n106880, n106881, n106882, n106883, n106884,
         n106885, n106886, n106887, n106888, n106889, n106890, n106891,
         n106892, n106893, n106894, n106895, n106896, n106897, n106898,
         n106899, n106900, n106901, n106902, n106903, n106904, n106905,
         n106906, n106907, n106908, n106909, n106910, n106911, n106912,
         n106913, n106914, n106915, n106916, n106917, n106918, n106919,
         n106920, n106921, n106922, n106923, n106924, n106925, n106926,
         n106927, n106928, n106929, n106930, n106931, n106932, n106933,
         n106934, n106935, n106936, n106937, n106938, n106939, n106940,
         n106941, n106942, n106943, n106944, n106945, n106946, n106947,
         n106948, n106949, n106950, n106951, n106952, n106953, n106954,
         n106955, n106956, n106957, n106958, n106959, n106960, n106961,
         n106962, n106963, n106964, n106965, n106966, n106967, n106968,
         n106969, n106970, n106971, n106972, n106973, n106974, n106975,
         n106976, n106977, n106978, n106979, n106980, n106981, n106982,
         n106983, n106984, n106985, n106986, n106987, n106988, n106989,
         n106990, n106991, n106992, n106993, n106994, n106995, n106996,
         n106997, n106998, n106999, n107000, n107001, n107002, n107003,
         n107004, n107005, n107006, n107007, n107008, n107009, n107010,
         n107011, n107012, n107013, n107014, n107015, n107016, n107017,
         n107018, n107019, n107020, n107021, n107022, n107023, n107024,
         n107025, n107026, n107027, n107028, n107029, n107030, n107031,
         n107032, n107033, n107034, n107035, n107036, n107037, n107038,
         n107039, n107040, n107041, n107042, n107043, n107044, n107045,
         n107046, n107047, n107048, n107049, n107050, n107051, n107052,
         n107053, n107054, n107055, n107056, n107057, n107058, n107059,
         n107060, n107061, n107062, n107063, n107064, n107065, n107066,
         n107067, n107068, n107069, n107070, n107071, n107072, n107073,
         n107074, n107075, n107076, n107077, n107078, n107079, n107080,
         n107081, n107082, n107083, n107084, n107085, n107086, n107087,
         n107088, n107089, n107090, n107091, n107092, n107093, n107094,
         n107095, n107096, n107097, n107098, n107099, n107100, n107101,
         n107102, n107103, n107104, n107105, n107106, n107107, n107108,
         n107109, n107110, n107111, n107112, n107113, n107114, n107115,
         n107116, n107117, n107118, n107119, n107120, n107121, n107122,
         n107123, n107124, n107125, n107126, n107127, n107128, n107129,
         n107130, n107131, n107132, n107133, n107134, n107135, n107136,
         n107137, n107138, n107139, n107140, n107141, n107142, n107143,
         n107144, n107145, n107146, n107147, n107148, n107149, n107150,
         n107151, n107152, n107153, n107154, n107155, n107156, n107157,
         n107158, n107159, n107160, n107161, n107162, n107163, n107164,
         n107165, n107166, n107167, n107168, n107169, n107170, n107171,
         n107172, n107173, n107174, n107175, n107176, n107177, n107178,
         n107179, n107180, n107181, n107182, n107183, n107184, n107185,
         n107186, n107187, n107188, n107189, n107190, n107191, n107192,
         n107193, n107194, n107195, n107196, n107197, n107198, n107199,
         n107200, n107201, n107202, n107203, n107204, n107205, n107206,
         n107207, n107208, n107209, n107210, n107211, n107212, n107213,
         n107214, n107215, n107216, n107217, n107218, n107219, n107220,
         n107221, n107222, n107223, n107224, n107225, n107226, n107227,
         n107228, n107229, n107230, n107231, n107232, n107233, n107234,
         n107235, n107236, n107237, n107238, n107239, n107240, n107241,
         n107242, n107243, n107244, n107245, n107246, n107247, n107248,
         n107249, n107250, n107251, n107252, n107253, n107254, n107255,
         n107256, n107257, n107258, n107259, n107260, n107261, n107262,
         n107263, n107264, n107265, n107266, n107267, n107268, n107269,
         n107270, n107271, n107272, n107273, n107274, n107275, n107276,
         n107277, n107278, n107279, n107280, n107281, n107282, n107283,
         n107284, n107285, n107286, n107287, n107288, n107289, n107290,
         n107291, n107292, n107293, n107294, n107295, n107296, n107297,
         n107298, n107299, n107300, n107301, n107302, n107303, n107304,
         n107305, n107306, n107307, n107308, n107309, n107310, n107311,
         n107312, n107313, n107314, n107315, n107316, n107317, n107318,
         n107319, n107320, n107321, n107322, n107323, n107324, n107325,
         n107326, n107327, n107328, n107329, n107330, n107331, n107332,
         n107333, n107334, n107335, n107336, n107337, n107338, n107339,
         n107340, n107341, n107342, n107343, n107344, n107345, n107346,
         n107347, n107348, n107349, n107350, n107351, n107352, n107353,
         n107354, n107355, n107356, n107357, n107358, n107359, n107360,
         n107361, n107362, n107363, n107364, n107365, n107366, n107367,
         n107368, n107369, n107370, n107371, n107372, n107373, n107374,
         n107375, n107376, n107377, n107378, n107379, n107380, n107381,
         n107382, n107383, n107384, n107385, n107386, n107387, n107388,
         n107389, n107390, n107391, n107392, n107393, n107394, n107395,
         n107396, n107397, n107398, n107399, n107400, n107401, n107402,
         n107403, n107404, n107405, n107406, n107407, n107408, n107409,
         n107410, n107411, n107412, n107413, n107414, n107415, n107416,
         n107417, n107418, n107419, n107420, n107421, n107422, n107423,
         n107424, n107425, n107426, n107427, n107428, n107429, n107430,
         n107431, n107432, n107433, n107434, n107435, n107436, n107437,
         n107438, n107439, n107440, n107441, n107442, n107443, n107444,
         n107445, n107446, n107447, n107448, n107449, n107450, n107451,
         n107452, n107453, n107454, n107455, n107456, n107457, n107458,
         n107459, n107460, n107461, n107462, n107463, n107464, n107465,
         n107466, n107467, n107468, n107469, n107470, n107471, n107472,
         n107473, n107474, n107475, n107476, n107477, n107478, n107479,
         n107480, n107481, n107482, n107483, n107484, n107485, n107486,
         n107487, n107488, n107489, n107490, n107491, n107492, n107493,
         n107494, n107495, n107496, n107497, n107498, n107499, n107500,
         n107501, n107502, n107503, n107504, n107505, n107506, n107507,
         n107508, n107509, n107510, n107511, n107512, n107513, n107514,
         n107515, n107516, n107517, n107518, n107519, n107520, n107521,
         n107522, n107523, n107524, n107525, n107526, n107527, n107528,
         n107529, n107530, n107531, n107532, n107533, n107534, n107535,
         n107536, n107537, n107538, n107539, n107540, n107541, n107542,
         n107543, n107544, n107545, n107546, n107547, n107548, n107549,
         n107550, n107551, n107552, n107553, n107554, n107555, n107556,
         n107557, n107558, n107559, n107560, n107561, n107562, n107563,
         n107564, n107565, n107566, n107567, n107568, n107569, n107570,
         n107571, n107572, n107573, n107574, n107575, n107576, n107577,
         n107578, n107579, n107580, n107581, n107582, n107583, n107584,
         n107585, n107586, n107587, n107588, n107589, n107590, n107591,
         n107592, n107593, n107594, n107595, n107596, n107597, n107598,
         n107599, n107600, n107601, n107602, n107603, n107604, n107605,
         n107606, n107607, n107608, n107609, n107610, n107611, n107612,
         n107613, n107614, n107615, n107616, n107617, n107618, n107619,
         n107620, n107621, n107622, n107623, n107624, n107625, n107626,
         n107627, n107628, n107629, n107630, n107631, n107632, n107633,
         n107634, n107635, n107636, n107637, n107638, n107639, n107640,
         n107641, n107642, n107643, n107644, n107645, n107646, n107647,
         n107648, n107649, n107650, n107651, n107652, n107653, n107654,
         n107655, n107656, n107657, n107658, n107659, n107660, n107661,
         n107662, n107663, n107664, n107665, n107666, n107667, n107668,
         n107669, n107670, n107671, n107672, n107673, n107674, n107675,
         n107676, n107677, n107678, n107679, n107680, n107681, n107682,
         n107683, n107684, n107685, n107686, n107687, n107688, n107689,
         n107690, n107691, n107692, n107693, n107694, n107695, n107696,
         n107697, n107698, n107699, n107700, n107701, n107702, n107703,
         n107704, n107705, n107706, n107707, n107708, n107709, n107710,
         n107711, n107712, n107713, n107714, n107715, n107716, n107717,
         n107718, n107719, n107720, n107721, n107722, n107723, n107724,
         n107725, n107726, n107727, n107728, n107729, n107730, n107731,
         n107732, n107733, n107734, n107735, n107736, n107737, n107738,
         n107739, n107740, n107741, n107742, n107743, n107744, n107745,
         n107746, n107747, n107748, n107749, n107750, n107751, n107752,
         n107753, n107754, n107755, n107756, n107757, n107758, n107759,
         n107760, n107761, n107762, n107763, n107764, n107765, n107766,
         n107767, n107768, n107769, n107770, n107771, n107772, n107773,
         n107774, n107775, n107776, n107777, n107778, n107779, n107780,
         n107781, n107782, n107783, n107784, n107785, n107786, n107787,
         n107788, n107789, n107790, n107791, n107792, n107793, n107794,
         n107795, n107796, n107797, n107798, n107799, n107800, n107801,
         n107802, n107803, n107804, n107805, n107806, n107807, n107808,
         n107809, n107810, n107811, n107812, n107813, n107814, n107815,
         n107816, n107817, n107818, n107819, n107820, n107821, n107822,
         n107823, n107824, n107825, n107826, n107827, n107828, n107829,
         n107830, n107831, n107832, n107833, n107834, n107835, n107836,
         n107837, n107838, n107839, n107840, n107841, n107842, n107843,
         n107844, n107845, n107846, n107847, n107848, n107849, n107850,
         n107851, n107852, n107853, n107854, n107855, n107856, n107857,
         n107858, n107859, n107860, n107861, n107862, n107863, n107864,
         n107865, n107866, n107867, n107868, n107869, n107870, n107871,
         n107872, n107873, n107874, n107875, n107876, n107877, n107878,
         n107879, n107880, n107881, n107882, n107883, n107884, n107885,
         n107886, n107887, n107888, n107889, n107890, n107891, n107892,
         n107893, n107894, n107895, n107896, n107897, n107898, n107899,
         n107900, n107901, n107902, n107903, n107904, n107905, n107906,
         n107907, n107908, n107909, n107910, n107911, n107912, n107913,
         n107914, n107915, n107916, n107917, n107918, n107919, n107920,
         n107921, n107922, n107923, n107924, n107925, n107926, n107927,
         n107928, n107929, n107930, n107931, n107932, n107933, n107934,
         n107935, n107936, n107937, n107938, n107939, n107940, n107941,
         n107942, n107943, n107944, n107945, n107946, n107947, n107948,
         n107949, n107950, n107951, n107952, n107953, n107954, n107955,
         n107956, n107957, n107958, n107959, n107960, n107961, n107962,
         n107963, n107964, n107965, n107966, n107967, n107968, n107969,
         n107970, n107971, n107972, n107973, n107974, n107975, n107976,
         n107977, n107978, n107979, n107980, n107981, n107982, n107983,
         n107984, n107985, n107986, n107987, n107988, n107989, n107990,
         n107991, n107992, n107993, n107994, n107995, n107996, n107997,
         n107998, n107999, n108000, n108001, n108002, n108003, n108004,
         n108005, n108006, n108007, n108008, n108009, n108010, n108011,
         n108012, n108013, n108014, n108015, n108016, n108017, n108018,
         n108019, n108020, n108021, n108022, n108023, n108024, n108025,
         n108026, n108027, n108028, n108029, n108030, n108031, n108032,
         n108033, n108034, n108035, n108036, n108037, n108038, n108039,
         n108040, n108041, n108042, n108043, n108044, n108045, n108046,
         n108047, n108048, n108049, n108050, n108051, n108052, n108053,
         n108054, n108055, n108056, n108057, n108058, n108059, n108060,
         n108061, n108062, n108063, n108064, n108065, n108066, n108067,
         n108068, n108069, n108070, n108071, n108072, n108073, n108074,
         n108075, n108076, n108077, n108078, n108079, n108080, n108081,
         n108082, n108083, n108084, n108085, n108086, n108087, n108088,
         n108089, n108090, n108091, n108092, n108093, n108094, n108095,
         n108096, n108097, n108098, n108099, n108100, n108101, n108102,
         n108103, n108104, n108105, n108106, n108107, n108108, n108109,
         n108110, n108111, n108112, n108113, n108114, n108115, n108116,
         n108117, n108118, n108119, n108120, n108121, n108122, n108123,
         n108124, n108125, n108126, n108127, n108128, n108129, n108130,
         n108131, n108132, n108133, n108134, n108135, n108136, n108137,
         n108138, n108139, n108140, n108141, n108142, n108143, n108144,
         n108145, n108146, n108147, n108148, n108149, n108150, n108151,
         n108152, n108153, n108154, n108155, n108156, n108157, n108158,
         n108159, n108160, n108161, n108162, n108163, n108164, n108165,
         n108166, n108167, n108168, n108169, n108170, n108171, n108172,
         n108173, n108174, n108175, n108176, n108177, n108178, n108179,
         n108180, n108181, n108182, n108183, n108184, n108185, n108186,
         n108187, n108188, n108189, n108190, n108191, n108192, n108193,
         n108194, n108195, n108196, n108197, n108198, n108199, n108200,
         n108201, n108202, n108203, n108204, n108205, n108206, n108207,
         n108208, n108209, n108210, n108211, n108212, n108213, n108214,
         n108215, n108216, n108217, n108218, n108219, n108220, n108221,
         n108222, n108223, n108224, n108225, n108226, n108227, n108228,
         n108229, n108230, n108231, n108232, n108233, n108234, n108235,
         n108236, n108237, n108238, n108239, n108240, n108241, n108242,
         n108243, n108244, n108245, n108246, n108247, n108248, n108249,
         n108250, n108251, n108252, n108253, n108254, n108255, n108256,
         n108257, n108258, n108259, n108260, n108261, n108262, n108263,
         n108264, n108265, n108266, n108267, n108268, n108269, n108270,
         n108271, n108272, n108273, n108274, n108275, n108276, n108277,
         n108278, n108279, n108280, n108281, n108282, n108283, n108284,
         n108285, n108286, n108287, n108288, n108289, n108290, n108291,
         n108292, n108293, n108294, n108295, n108296, n108297, n108298,
         n108299, n108300, n108301, n108302, n108303, n108304, n108305,
         n108306, n108307, n108308, n108309, n108310, n108311, n108312,
         n108313, n108314, n108315, n108316, n108317, n108318, n108319,
         n108320, n108321, n108322, n108323, n108324, n108325, n108326,
         n108327, n108328, n108329, n108330, n108331, n108332, n108333,
         n108334, n108335, n108336, n108337, n108338, n108339, n108340,
         n108341, n108342, n108343, n108344, n108345, n108346, n108347,
         n108348, n108349, n108350, n108351, n108352, n108353, n108354,
         n108355, n108356, n108357, n108358, n108359, n108360, n108361,
         n108362, n108363, n108364, n108365, n108366, n108367, n108368,
         n108369, n108370, n108371, n108372, n108373, n108374, n108375,
         n108376, n108377, n108378, n108379, n108380, n108381, n108382,
         n108383, n108384, n108385, n108386, n108387, n108388, n108389,
         n108390, n108391, n108392, n108393, n108394, n108395, n108396,
         n108397, n108398, n108399, n108400, n108401, n108402, n108403,
         n108404, n108405, n108406, n108407, n108408, n108409, n108410,
         n108411, n108412, n108413, n108414, n108415, n108416, n108417,
         n108418, n108419, n108420, n108421, n108422, n108423, n108424,
         n108425, n108426, n108427, n108428, n108429, n108430, n108431,
         n108432, n108433, n108434, n108435, n108436, n108437, n108438,
         n108439, n108440, n108441, n108442, n108443, n108444, n108445,
         n108446, n108447, n108448, n108449, n108450, n108451, n108452,
         n108453, n108454, n108455, n108456, n108457, n108458, n108459,
         n108460, n108461, n108462, n108463, n108464, n108465, n108466,
         n108467, n108468, n108469, n108470, n108471, n108472, n108473,
         n108474, n108475, n108476, n108477, n108478, n108479, n108480,
         n108481, n108482, n108483, n108484, n108485, n108486, n108487,
         n108488, n108489, n108490, n108491, n108492, n108493, n108494,
         n108495, n108496, n108497, n108498, n108499, n108500, n108501,
         n108502, n108503, n108504, n108505, n108506, n108507, n108508,
         n108509, n108510, n108511, n108512, n108513, n108514, n108515,
         n108516, n108517, n108518, n108519, n108520, n108521, n108522,
         n108523, n108524, n108525, n108526, n108527, n108528, n108529,
         n108530, n108531, n108532, n108533, n108534, n108535, n108536,
         n108537, n108538, n108539, n108540, n108541, n108542, n108543,
         n108544, n108545, n108546, n108547, n108548, n108549, n108550,
         n108551, n108552, n108553, n108554, n108555, n108556, n108557,
         n108558, n108559, n108560, n108561, n108562, n108563, n108564,
         n108565, n108566, n108567, n108568, n108569, n108570, n108571,
         n108572, n108573, n108574, n108575, n108576, n108577, n108578,
         n108579, n108580, n108581, n108582, n108583, n108584, n108585,
         n108586, n108587, n108588, n108589, n108590, n108591, n108592,
         n108593, n108594, n108595, n108596, n108597, n108598, n108599,
         n108600, n108601, n108602, n108603, n108604, n108605, n108606,
         n108607, n108608, n108609, n108610, n108611, n108612, n108613,
         n108614, n108615, n108616, n108617, n108618, n108619, n108620,
         n108621, n108622, n108623, n108624, n108625, n108626, n108627,
         n108628, n108629, n108630, n108631, n108632, n108633, n108634,
         n108635, n108636, n108637, n108638, n108639, n108640, n108641,
         n108642, n108643, n108644, n108645, n108646, n108647, n108648,
         n108649, n108650, n108651, n108652, n108653, n108654, n108655,
         n108656, n108657, n108658, n108659, n108660, n108661, n108662,
         n108663, n108664, n108665, n108666, n108667, n108668, n108669,
         n108670, n108671, n108672, n108673, n108674, n108675, n108676,
         n108677, n108678, n108679, n108680, n108681, n108682, n108683,
         n108684, n108685, n108686, n108687, n108688, n108689, n108690,
         n108691, n108692, n108693, n108694, n108695, n108696, n108697,
         n108698, n108699, n108700, n108701, n108702, n108703, n108704,
         n108705, n108706, n108707, n108708, n108709, n108710, n108711,
         n108712, n108713, n108714, n108715, n108716, n108717, n108718,
         n108719, n108720, n108721, n108722, n108723, n108724, n108725,
         n108726, n108727, n108728, n108729, n108730, n108731, n108732,
         n108733, n108734, n108735, n108736, n108737, n108738, n108739,
         n108740, n108741, n108742, n108743, n108744, n108745, n108746,
         n108747, n108748, n108749, n108750, n108751, n108752, n108753,
         n108754, n108755, n108756, n108757, n108758, n108759, n108760,
         n108761, n108762, n108763, n108764, n108765, n108766, n108767,
         n108768, n108769, n108770, n108771, n108772, n108773, n108774,
         n108775, n108776, n108777, n108778, n108779, n108780, n108781,
         n108782, n108783, n108784, n108785, n108786, n108787, n108788,
         n108789, n108790, n108791, n108792, n108793, n108794, n108795,
         n108796, n108797, n108798, n108799, n108800, n108801, n108802,
         n108803, n108804, n108805, n108806, n108807, n108808, n108809,
         n108810, n108811, n108812, n108813, n108814, n108815, n108816,
         n108817, n108818, n108819, n108820, n108821, n108822, n108823,
         n108824, n108825, n108826, n108827, n108828, n108829, n108830,
         n108831, n108832, n108833, n108834, n108835, n108836, n108837,
         n108838, n108839, n108840, n108841, n108842, n108843, n108844,
         n108845, n108846, n108847, n108848, n108849, n108850, n108851,
         n108852, n108853, n108854, n108855, n108856, n108857, n108858,
         n108859, n108860, n108861, n108862, n108863, n108864, n108865,
         n108866, n108867, n108868, n108869, n108870, n108871, n108872,
         n108873, n108874, n108875, n108876, n108877, n108878, n108879,
         n108880, n108881, n108882, n108883, n108884, n108885, n108886,
         n108887, n108888, n108889, n108890, n108891, n108892, n108893,
         n108894, n108895, n108896, n108897, n108898, n108899, n108900,
         n108901, n108902, n108903, n108904, n108905, n108906, n108907,
         n108908, n108909, n108910, n108911, n108912, n108913, n108914,
         n108915, n108916, n108917, n108918, n108919, n108920, n108921,
         n108922, n108923, n108924, n108925, n108926, n108927, n108928,
         n108929, n108930, n108931, n108932, n108933, n108934, n108935,
         n108936, n108937, n108938, n108939, n108940, n108941, n108942,
         n108943, n108944, n108945, n108946, n108947, n108948, n108949,
         n108950, n108951, n108952, n108953, n108954, n108955, n108956,
         n108957, n108958, n108959, n108960, n108961, n108962, n108963,
         n108964, n108965, n108966, n108967, n108968, n108969, n108970,
         n108971, n108972, n108973, n108974, n108975, n108976, n108977,
         n108978, n108979, n108980, n108981, n108982, n108983, n108984,
         n108985, n108986, n108987, n108988, n108989, n108990, n108991,
         n108992, n108993, n108994, n108995, n108996, n108997, n108998,
         n108999, n109000, n109001, n109002, n109003, n109004, n109005,
         n109006, n109007, n109008, n109009, n109010, n109011, n109012,
         n109013, n109014, n109015, n109016, n109017, n109018, n109019,
         n109020, n109021, n109022, n109023, n109024, n109025, n109026,
         n109027, n109028, n109029, n109030, n109031, n109032, n109033,
         n109034, n109035, n109036, n109037, n109038, n109039, n109040,
         n109041, n109042, n109043, n109044, n109045, n109046, n109047,
         n109048, n109049, n109050, n109051, n109052, n109053, n109054,
         n109055, n109056, n109057, n109058, n109059, n109060, n109061,
         n109062, n109063, n109064, n109065, n109066, n109067, n109068,
         n109069, n109070, n109071, n109072, n109073, n109074, n109075,
         n109076, n109077, n109078, n109079, n109080, n109081, n109082,
         n109083, n109084, n109085, n109086, n109087, n109088, n109089,
         n109090, n109091, n109092, n109093, n109094, n109095, n109096,
         n109097, n109098, n109099, n109100, n109101, n109102, n109103,
         n109104, n109105, n109106, n109107, n109108, n109109, n109110,
         n109111, n109112, n109113, n109114, n109115, n109116, n109117,
         n109118, n109119, n109120, n109121, n109122, n109123, n109124,
         n109125, n109126, n109127, n109128, n109129, n109130, n109131,
         n109132, n109133, n109134, n109135, n109136, n109137, n109138,
         n109139, n109140, n109141, n109142, n109143, n109144, n109145,
         n109146, n109147, n109148, n109149, n109150, n109151, n109152,
         n109153, n109154, n109155, n109156, n109157, n109158, n109159,
         n109160, n109161, n109162, n109163, n109164, n109165, n109166,
         n109167, n109168, n109169, n109170, n109171, n109172, n109173,
         n109174, n109175, n109176, n109177, n109178, n109179, n109180,
         n109181, n109182, n109183, n109184, n109185, n109186, n109187,
         n109188, n109189, n109190, n109191, n109192, n109193, n109194,
         n109195, n109196, n109197, n109198, n109199, n109200, n109201,
         n109202, n109203, n109204, n109205, n109206, n109207, n109208,
         n109209, n109210, n109211, n109212, n109213, n109214, n109215,
         n109216, n109217, n109218, n109219, n109220, n109221, n109222,
         n109223, n109224, n109225, n109226, n109227, n109228, n109229,
         n109230, n109231, n109232, n109233, n109234, n109235, n109236,
         n109237, n109238, n109239, n109240, n109241, n109242, n109243,
         n109244, n109245, n109246, n109247, n109248, n109249, n109250,
         n109251, n109252, n109253, n109254, n109255, n109256, n109257,
         n109258, n109259, n109260, n109261, n109262, n109263, n109264,
         n109265, n109266, n109267, n109268, n109269, n109270, n109271,
         n109272, n109273, n109274, n109275, n109276, n109277, n109278,
         n109279, n109280, n109281, n109282, n109283, n109284, n109285,
         n109286, n109287, n109288, n109289, n109290, n109291, n109292,
         n109293, n109294, n109295, n109296, n109297, n109298, n109299,
         n109300, n109301, n109302, n109303, n109304, n109305, n109306,
         n109307, n109308, n109309, n109310, n109311, n109312, n109313,
         n109314, n109315, n109316, n109317, n109318, n109319, n109320,
         n109321, n109322, n109323, n109324, n109325, n109326, n109327,
         n109328, n109329, n109330, n109331, n109332, n109333, n109334,
         n109335, n109336, n109337, n109338, n109339, n109340, n109341,
         n109342, n109343, n109344, n109345, n109346, n109347, n109348,
         n109349, n109350, n109351, n109352, n109353, n109354, n109355,
         n109356, n109357, n109358, n109359, n109360, n109361, n109362,
         n109363, n109364, n109365, n109366, n109367, n109368, n109369,
         n109370, n109371, n109372, n109373, n109374, n109375, n109376,
         n109377, n109378, n109379, n109380, n109381, n109382, n109383,
         n109384, n109385, n109386, n109387, n109388, n109389, n109390,
         n109391, n109392, n109393, n109394, n109395, n109396, n109397,
         n109398, n109399, n109400, n109401, n109402, n109403, n109404,
         n109405, n109406, n109407, n109408, n109409, n109410, n109411,
         n109412, n109413, n109414, n109415, n109416, n109417, n109418,
         n109419, n109420, n109421, n109422, n109423, n109424, n109425,
         n109426, n109427, n109428, n109429, n109430, n109431, n109432,
         n109433, n109434, n109435, n109436, n109437, n109438, n109439,
         n109440, n109441, n109442, n109443, n109444, n109445, n109446,
         n109447, n109448, n109449, n109450, n109451, n109452, n109453,
         n109454, n109455, n109456, n109457, n109458, n109459, n109460,
         n109461, n109462, n109463, n109464, n109465, n109466, n109467,
         n109468, n109469, n109470, n109471, n109472, n109473, n109474,
         n109475, n109476, n109477, n109478, n109479, n109480, n109481,
         n109482, n109483, n109484, n109485, n109486, n109487, n109488,
         n109489, n109490, n109491, n109492, n109493, n109494, n109495,
         n109496, n109497, n109498, n109499, n109500, n109501, n109502,
         n109503, n109504, n109505, n109506, n109507, n109508, n109509,
         n109510, n109511, n109512, n109513, n109514, n109515, n109516,
         n109517, n109518, n109519, n109520, n109521, n109522, n109523,
         n109524, n109525, n109526, n109527, n109528, n109529, n109530,
         n109531, n109532, n109533, n109534, n109535, n109536, n109537,
         n109538, n109539, n109540, n109541, n109542, n109543, n109544,
         n109545, n109546, n109547, n109548, n109549, n109550, n109551,
         n109552, n109553, n109554, n109555, n109556, n109557, n109558,
         n109559, n109560, n109561, n109562, n109563, n109564, n109565,
         n109566, n109567, n109568, n109569, n109570, n109571, n109572,
         n109573, n109574, n109575, n109576, n109577, n109578, n109579,
         n109580, n109581, n109582, n109583, n109584, n109585, n109586,
         n109587, n109588, n109589, n109590, n109591, n109592, n109593,
         n109594, n109595, n109596, n109597, n109598, n109599, n109600,
         n109601, n109602, n109603, n109604, n109605, n109606, n109607,
         n109608, n109609, n109610, n109611, n109612, n109613, n109614,
         n109615, n109616, n109617, n109618, n109619, n109620, n109621,
         n109622, n109623, n109624, n109625, n109626, n109627, n109628,
         n109629, n109630, n109631, n109632, n109633, n109634, n109635,
         n109636, n109637, n109638, n109639, n109640, n109641, n109642,
         n109643, n109644, n109645, n109646, n109647, n109648, n109649,
         n109650, n109651, n109652, n109653, n109654, n109655, n109656,
         n109657, n109658, n109659, n109660, n109661, n109662, n109663,
         n109664, n109665, n109666, n109667, n109668, n109669, n109670,
         n109671, n109672, n109673, n109674, n109675, n109676, n109677,
         n109678, n109679, n109680, n109681, n109682, n109683, n109684,
         n109685, n109686, n109687, n109688, n109689, n109690, n109691,
         n109692, n109693, n109694, n109695, n109696, n109697, n109698,
         n109699, n109700, n109701, n109702, n109703, n109704, n109705,
         n109706, n109707, n109708, n109709, n109710, n109711, n109712,
         n109713, n109714, n109715, n109716, n109717, n109718, n109719,
         n109720, n109721, n109722, n109723, n109724, n109725, n109726,
         n109727, n109728, n109729, n109730, n109731, n109732, n109733,
         n109734, n109735, n109736, n109737, n109738, n109739, n109740,
         n109741, n109742, n109743, n109744, n109745, n109746, n109747,
         n109748, n109749, n109750, n109751, n109752, n109753, n109754,
         n109755, n109756, n109757, n109758, n109759, n109760, n109761,
         n109762, n109763, n109764, n109765, n109766, n109767, n109768,
         n109769, n109770, n109771, n109772, n109773, n109774, n109775,
         n109776, n109777, n109778, n109779, n109780, n109781, n109782,
         n109783, n109784, n109785, n109786, n109787, n109788, n109789,
         n109790, n109791, n109792, n109793, n109794, n109795, n109796,
         n109797, n109798, n109799, n109800, n109801, n109802, n109803,
         n109804, n109805, n109806, n109807, n109808, n109809, n109810,
         n109811, n109812, n109813, n109814, n109815, n109816, n109817,
         n109818, n109819, n109820, n109821, n109822, n109823, n109824,
         n109825, n109826, n109827, n109828, n109829, n109830, n109831,
         n109832, n109833, n109834, n109835, n109836, n109837, n109838,
         n109839, n109840, n109841, n109842, n109843, n109844, n109845,
         n109846, n109847, n109848, n109849, n109850, n109851, n109852,
         n109853, n109854, n109855, n109856, n109857, n109858, n109859,
         n109860, n109861, n109862, n109863, n109864, n109865, n109866,
         n109867, n109868, n109869, n109870, n109871, n109872, n109873,
         n109874, n109875, n109876, n109877, n109878, n109879, n109880,
         n109881, n109882, n109883, n109884, n109885, n109886, n109887,
         n109888, n109889, n109890, n109891, n109892, n109893, n109894,
         n109895, n109896, n109897, n109898, n109899, n109900, n109901,
         n109902, n109903, n109904, n109905, n109906, n109907, n109908,
         n109909, n109910, n109911, n109912, n109913, n109914, n109915,
         n109916, n109917, n109918, n109919, n109920, n109921, n109922,
         n109923, n109924, n109925, n109926, n109927, n109928, n109929,
         n109930, n109931, n109932, n109933, n109934, n109935, n109936,
         n109937, n109938, n109939, n109940, n109941, n109942, n109943,
         n109944, n109945, n109946, n109947, n109948, n109949, n109950,
         n109951, n109952, n109953, n109954, n109955, n109956, n109957,
         n109958, n109959, n109960, n109961, n109962, n109963, n109964,
         n109965, n109966, n109967, n109968, n109969, n109970, n109971,
         n109972, n109973, n109974, n109975, n109976, n109977, n109978,
         n109979, n109980, n109981, n109982, n109983, n109984, n109985,
         n109986, n109987, n109988, n109989, n109990, n109991, n109992,
         n109993, n109994, n109995, n109996, n109997, n109998, n109999,
         n110000, n110001, n110002, n110003, n110004, n110005, n110006,
         n110007, n110008, n110009, n110010, n110011, n110012, n110013,
         n110014, n110015, n110016, n110017, n110018, n110019, n110020,
         n110021, n110022, n110023, n110024, n110025, n110026, n110027,
         n110028, n110029, n110030, n110031, n110032, n110033, n110034,
         n110035, n110036, n110037, n110038, n110039, n110040, n110041,
         n110042, n110043, n110044, n110045, n110046, n110047, n110048,
         n110049, n110050, n110051, n110052, n110053, n110054, n110055,
         n110056, n110057, n110058, n110059, n110060, n110061, n110062,
         n110063, n110064, n110065, n110066, n110067, n110068, n110069,
         n110070, n110071, n110072, n110073, n110074, n110075, n110076,
         n110077, n110078, n110079, n110080, n110081, n110082, n110083,
         n110084, n110085, n110086, n110087, n110088, n110089, n110090,
         n110091, n110092, n110093, n110094, n110095, n110096, n110097,
         n110098, n110099, n110100, n110101, n110102, n110103, n110104,
         n110105, n110106, n110107, n110108, n110109, n110110, n110111,
         n110112, n110113, n110114, n110115, n110116, n110117, n110118,
         n110119, n110120, n110121, n110122, n110123, n110124, n110125,
         n110126, n110127, n110128, n110129, n110130, n110131, n110132,
         n110133, n110134, n110135, n110136, n110137, n110138, n110139,
         n110140, n110141, n110142, n110143, n110144, n110145, n110146,
         n110147, n110148, n110149, n110150, n110151, n110152, n110153,
         n110154, n110155, n110156, n110157, n110158, n110159, n110160,
         n110161, n110162, n110163, n110164, n110165, n110166, n110167,
         n110168, n110169, n110170, n110171, n110172, n110173, n110174,
         n110175, n110176, n110177, n110178, n110179, n110180, n110181,
         n110182, n110183, n110184, n110185, n110186, n110187, n110188,
         n110189, n110190, n110191, n110192, n110193, n110194, n110195,
         n110196, n110197, n110198, n110199, n110200, n110201, n110202,
         n110203, n110204, n110205, n110206, n110207, n110208, n110209,
         n110210, n110211, n110212, n110213, n110214, n110215, n110216,
         n110217, n110218, n110219, n110220, n110221, n110222, n110223,
         n110224, n110225, n110226, n110227, n110228, n110229, n110230,
         n110231, n110232, n110233, n110234, n110235, n110236, n110237,
         n110238, n110239, n110240, n110241, n110242, n110243, n110244,
         n110245, n110246, n110247, n110248, n110249, n110250, n110251,
         n110252, n110253, n110254, n110255, n110256, n110257, n110258,
         n110259, n110260, n110261, n110262, n110263, n110264, n110265,
         n110266, n110267, n110268, n110269, n110270, n110271, n110272,
         n110273, n110274, n110275, n110276, n110277, n110278, n110279,
         n110280, n110281, n110282, n110283, n110284, n110285, n110286,
         n110287, n110288, n110289, n110290, n110291, n110292, n110293,
         n110294, n110295, n110296, n110297, n110298, n110299, n110300,
         n110301, n110302, n110303, n110304, n110305, n110306, n110307,
         n110308, n110309, n110310, n110311, n110312, n110313, n110314,
         n110315, n110316, n110317, n110318, n110319, n110320, n110321,
         n110322, n110323, n110324, n110325, n110326, n110327, n110328,
         n110329, n110330, n110331, n110332, n110333, n110334, n110335,
         n110336, n110337, n110338, n110339, n110340, n110341, n110342,
         n110343, n110344, n110345, n110346, n110347, n110348, n110349,
         n110350, n110351, n110352, n110353, n110354, n110355, n110356,
         n110357, n110358, n110359, n110360, n110361, n110362, n110363,
         n110364, n110365, n110366, n110367, n110368, n110369, n110370,
         n110371, n110372, n110373, n110374, n110375, n110376, n110377,
         n110378, n110379, n110380, n110381, n110382, n110383, n110384,
         n110385, n110386, n110387, n110388, n110389, n110390, n110391,
         n110392, n110393, n110394, n110395, n110396, n110397, n110398,
         n110399, n110400, n110401, n110402, n110403, n110404, n110405,
         n110406, n110407, n110408, n110409, n110410, n110411, n110412,
         n110413, n110414, n110415, n110416, n110417, n110418, n110419,
         n110420, n110421, n110422, n110423, n110424, n110425, n110426,
         n110427, n110428, n110429, n110430, n110431, n110432, n110433,
         n110434, n110435, n110436, n110437, n110438, n110439, n110440,
         n110441, n110442, n110443, n110444, n110445, n110446, n110447,
         n110448, n110449, n110450, n110451, n110452, n110453, n110454,
         n110455, n110456, n110457, n110458, n110459, n110460, n110461,
         n110462, n110463, n110464, n110465, n110466, n110467, n110468,
         n110469, n110470, n110471, n110472, n110473, n110474, n110475,
         n110476, n110477, n110478, n110479, n110480, n110481, n110482,
         n110483, n110484, n110485, n110486, n110487, n110488, n110489,
         n110490, n110491, n110492, n110493, n110494, n110495, n110496,
         n110497, n110498, n110499, n110500, n110501, n110502, n110503,
         n110504, n110505, n110506, n110507, n110508, n110509, n110510,
         n110511, n110512, n110513, n110514, n110515, n110516, n110517,
         n110518, n110519, n110520, n110521, n110522, n110523, n110524,
         n110525, n110526, n110527, n110528, n110529, n110530, n110531,
         n110532, n110533, n110534, n110535, n110536, n110537, n110538,
         n110539, n110540, n110541, n110542, n110543, n110544, n110545,
         n110546, n110547, n110548, n110549, n110550, n110551, n110552,
         n110553, n110554, n110555, n110556, n110557, n110558, n110559,
         n110560, n110561, n110562, n110563, n110564, n110565, n110566,
         n110567, n110568, n110569, n110570, n110571, n110572, n110573,
         n110574, n110575, n110576, n110577, n110578, n110579, n110580,
         n110581, n110582, n110583, n110584, n110585, n110586, n110587,
         n110588, n110589, n110590, n110591, n110592, n110593, n110594,
         n110595, n110596, n110597, n110598, n110599, n110600, n110601,
         n110602, n110603, n110604, n110605, n110606, n110607, n110608,
         n110609, n110610, n110611, n110612, n110613, n110614, n110615,
         n110616, n110617, n110618, n110619, n110620, n110621, n110622,
         n110623, n110624, n110625, n110626, n110627, n110628, n110629,
         n110630, n110631, n110632, n110633, n110634, n110635, n110636,
         n110637, n110638, n110639, n110640, n110641, n110642, n110643,
         n110644, n110645, n110646, n110647, n110648, n110649, n110650,
         n110651, n110652, n110653, n110654, n110655, n110656, n110657,
         n110658, n110659, n110660, n110661, n110662, n110663, n110664,
         n110665, n110666, n110667, n110668, n110669, n110670, n110671,
         n110672, n110673, n110674, n110675, n110676, n110677, n110678,
         n110679, n110680, n110681, n110682, n110683, n110684, n110685,
         n110686, n110687, n110688, n110689, n110690, n110691, n110692,
         n110693, n110694, n110695, n110696, n110697, n110698, n110699,
         n110700, n110701, n110702, n110703, n110704, n110705, n110706,
         n110707, n110708, n110709, n110710, n110711, n110712, n110713,
         n110714, n110715, n110716, n110717, n110718, n110719, n110720,
         n110721, n110722, n110723, n110724, n110725, n110726, n110727,
         n110728, n110729, n110730, n110731, n110732, n110733, n110734,
         n110735, n110736, n110737, n110738, n110739, n110740, n110741,
         n110742, n110743, n110744, n110745, n110746, n110747, n110748,
         n110749, n110750, n110751, n110752, n110753, n110754, n110755,
         n110756, n110757, n110758, n110759, n110760, n110761, n110762,
         n110763, n110764, n110765, n110766, n110767, n110768, n110769,
         n110770, n110771, n110772, n110773, n110774, n110775, n110776,
         n110777, n110778, n110779, n110780, n110781, n110782, n110783,
         n110784, n110785, n110786, n110787, n110788, n110789, n110790,
         n110791, n110792, n110793, n110794, n110795, n110796, n110797,
         n110798, n110799, n110800, n110801, n110802, n110803, n110804,
         n110805, n110806, n110807, n110808, n110809, n110810, n110811,
         n110812, n110813, n110814, n110815, n110816, n110817, n110818,
         n110819, n110820, n110821, n110822, n110823, n110824, n110825,
         n110826, n110827, n110828, n110829, n110830, n110831, n110832,
         n110833, n110834, n110835, n110836, n110837, n110838, n110839,
         n110840, n110841, n110842, n110843, n110844, n110845, n110846,
         n110847, n110848, n110849, n110850, n110851, n110852, n110853,
         n110854, n110855, n110856, n110857, n110858, n110859, n110860,
         n110861, n110862, n110863, n110864, n110865, n110866, n110867,
         n110868, n110869, n110870, n110871, n110872, n110873, n110874,
         n110875, n110876, n110877, n110878, n110879, n110880, n110881,
         n110882, n110883, n110884, n110885, n110886, n110887, n110888,
         n110889, n110890, n110891, n110892, n110893, n110894, n110895,
         n110896, n110897, n110898, n110899, n110900, n110901, n110902,
         n110903, n110904, n110905, n110906, n110907, n110908, n110909,
         n110910, n110911, n110912, n110913, n110914, n110915, n110916,
         n110917, n110918, n110919, n110920, n110921, n110922, n110923,
         n110924, n110925, n110926, n110927, n110928, n110929, n110930,
         n110931, n110932, n110933, n110934, n110935, n110936, n110937,
         n110938, n110939, n110940, n110941, n110942, n110943, n110944,
         n110945, n110946, n110947, n110948, n110949, n110950, n110951,
         n110952, n110953, n110954, n110955, n110956, n110957, n110958,
         n110959, n110960, n110961, n110962, n110963, n110964, n110965,
         n110966, n110967, n110968, n110969, n110970, n110971, n110972,
         n110973, n110974, n110975, n110976, n110977, n110978, n110979,
         n110980, n110981, n110982, n110983, n110984, n110985, n110986,
         n110987, n110988, n110989, n110990, n110991, n110992, n110993,
         n110994, n110995, n110996, n110997, n110998, n110999, n111000,
         n111001, n111002, n111003, n111004, n111005, n111006, n111007,
         n111008, n111009, n111010, n111011, n111012, n111013, n111014,
         n111015, n111016, n111017, n111018, n111019, n111020, n111021,
         n111022, n111023, n111024, n111025, n111026, n111027, n111028,
         n111029, n111030, n111031, n111032, n111033, n111034, n111035,
         n111036, n111037, n111038, n111039, n111040, n111041, n111042,
         n111043, n111044, n111045, n111046, n111047, n111048, n111049,
         n111050, n111051, n111052, n111053, n111054, n111055, n111056,
         n111057, n111058, n111059, n111060, n111061, n111062, n111063,
         n111064, n111065, n111066, n111067, n111068, n111069, n111070,
         n111071, n111072, n111073, n111074, n111075, n111076, n111077,
         n111078, n111079, n111080, n111081, n111082, n111083, n111084,
         n111085, n111086, n111087, n111088, n111089, n111090, n111091,
         n111092, n111093, n111094, n111095, n111096, n111097, n111098,
         n111099, n111100, n111101, n111102, n111103, n111104, n111105,
         n111106, n111107, n111108, n111109, n111110, n111111, n111112,
         n111113, n111114, n111115, n111116, n111117, n111118, n111119,
         n111120, n111121, n111122, n111123, n111124, n111125, n111126,
         n111127, n111128, n111129, n111130, n111131, n111132, n111133,
         n111134, n111135, n111136, n111137, n111138, n111139, n111140,
         n111141, n111142, n111143, n111144, n111145, n111146, n111147,
         n111148, n111149, n111150, n111151, n111152, n111153, n111154,
         n111155, n111156, n111157, n111158, n111159, n111160, n111161;
  wire   [31:0] \DLX_Datapath/next_ALUOut_EXMEM ;
  wire   [31:0] \DLX_Datapath/MUX_HDU_ALUInB ;
  wire   [31:0] \DLX_Datapath/MUX_HDU_ALUInA ;
  wire   [31:0] \DLX_Datapath/next_B_IDEX ;
  wire   [1:0] \DLX_Datapath/RegisterFile/next_to_transfer ;
  wire   [2:0] \DLX_Datapath/RegisterFile/old_CWP1 ;
  wire   [1:0] \DLX_Datapath/ArithLogUnit/sel_shf ;
  wire   [4:0] \DLX_Datapath/ArithLogUnit/B_shf ;
  wire   [31:0] \DLX_Datapath/ArithLogUnit/A_shf ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/sel_log ;
  wire   [31:0] \DLX_Datapath/ArithLogUnit/B_log ;
  wire   [31:0] \DLX_Datapath/ArithLogUnit/A_log ;
  wire   [31:0] \DLX_Datapath/ArithLogUnit/Sum_cmp ;
  wire   [15:0] \DLX_Datapath/ArithLogUnit/B_mul ;
  wire   [31:0] \DLX_Datapath/ArithLogUnit/B_add ;
  wire   [31:0] \DLX_Datapath/ArithLogUnit/A_add ;
  wire   [3:0] \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 ;
  wire   [3:0] \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_1 ;
  wire   [3:0] \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_0 ;
  wire   [3:0] \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_1 ;
  wire   [3:0] \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_0 ;
  wire   [3:0] \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_1 ;
  wire   [3:0] \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_0 ;
  wire   [3:0] \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 ;
  wire   [3:0] \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 ;
  wire   [3:0] \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 ;
  wire   [3:0] \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 ;
  wire   [3:0] \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 ;
  wire   [3:0] \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 ;
  wire   [3:0] \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_1 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_0 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_1 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_0 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_1 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_0 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_1 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_0 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_1 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_0 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_1 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_0 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_1 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_0 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_1 ;
  wire   [3:0] \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_0 ;
  wire   [4:0] \DLX_ControlUnit/ALUop2 ;
  wire   [4:0] \DLX_ControlUnit/cw4 ;
  wire   [13:0] \DLX_ControlUnit/cw3 ;
  wire   [17:0] \DLX_ControlUnit/cw2 ;
  tri   [127:0] stackBus_Out;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign PC_out[7] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0  [3];
  assign PC_out[6] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0  [2];
  assign PC_out[5] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0  [1];
  assign PC_out[4] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0  [0];
  assign PC_out[11] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0  [3];
  assign PC_out[10] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0  [2];
  assign PC_out[9] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0  [1];
  assign PC_out[8] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0  [0];
  assign PC_out[15] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0  [3];
  assign PC_out[14] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0  [2];
  assign PC_out[13] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0  [1];
  assign PC_out[12] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0  [0];
  assign PC_out[19] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0  [3];
  assign PC_out[18] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0  [2];
  assign PC_out[17] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0  [1];
  assign PC_out[16] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0  [0];
  assign PC_out[23] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0  [3];
  assign PC_out[22] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0  [2];
  assign PC_out[21] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0  [1];
  assign PC_out[20] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0  [0];
  assign PC_out[27] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0  [3];
  assign PC_out[26] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0  [2];
  assign PC_out[25] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0  [1];
  assign PC_out[24] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0  [0];
  assign PC_out[31] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0  [3];
  assign PC_out[30] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0  [2];
  assign PC_out[29] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0  [1];
  assign PC_out[28] = \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0  [0];

  DFFR_X2 \DLX_Datapath/RegisterFile/SWP_reg[2]  ( .D(n60369), .CK(Clk), .RN(
        n106373), .Q(n106753), .QN(n59515) );
  DFFR_X2 \DLX_Datapath/RegisterFile/SWP_reg[1]  ( .D(n60370), .CK(Clk), .RN(
        n106436), .Q(n106764), .QN(n59514) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[0]  ( .D(n106549), .CK(Clk), .RN(Rst), 
        .Q(n106765), .QN(n100462) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[0]  ( .D(n106631), .CK(Clk), .RN(Rst), 
        .Q(n69289) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[0]  ( .D(n59081), .CK(Clk), .RN(Rst), 
        .Q(n106766), .QN(n100416) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26827 ), .CK(Clk), .RN(Rst), .Q(n106767), 
        .QN(n102767) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[0]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(
        \DLX_Datapath/RegisterFile/N46866 ), .Q(\DLX_Datapath/next_B_IDEX [0])
         );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[0]  ( .D(n106663), .CK(Clk), .RN(Rst), .Q(
        n69292) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[0]  ( .D(
        \DLX_Datapath/ArithLogUnit/N193 ), .GN(n106360), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [0]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[0]  ( .D(n104325), .CK(Clk), .RN(Rst), 
        .Q(DataAddr[0]), .QN(n58728) );
  DFFR_X2 \DLX_Datapath/PC_reg[0]  ( .D(n60325), .CK(Clk), .RN(Rst), .Q(
        PC_out[0]), .QN(net2465273) );
  DFFR_X2 \DLX_Datapath/PC_IFID_reg[0]  ( .D(n60229), .CK(Clk), .RN(Rst), .Q(
        n106809), .QN(n59420) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[25][1]  ( .D(n60211), 
        .CK(Clk), .RN(Rst), .Q(n106812) );
  DFFR_X2 \DLX_Datapath/PC_reg[1]  ( .D(n60324), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_0/S_0[1] ), .QN(net2465147)
         );
  DFFR_X2 \DLX_Datapath/PC_reg[11]  ( .D(n60314), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [3]), .QN(n104499) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[19]  ( .D(n106530), .CK(Clk), .RN(Rst), 
        .Q(n106822) );
  DFFR_X2 \DLX_Datapath/PC_reg[19]  ( .D(n60306), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [3]), .QN(n57424) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[23]  ( .D(n106526), .CK(Clk), .RN(Rst), 
        .Q(n106824) );
  DFFR_X2 \DLX_Datapath/PC_reg[23]  ( .D(n60302), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [3]), .QN(n62191) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[31]  ( .D(n106518), .CK(Clk), .RN(Rst), 
        .Q(n106825) );
  DFFR_X2 \DLX_Datapath/PC_reg[31]  ( .D(n60294), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0 [3]), .QN(n57431) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[30]  ( .D(n106519), .CK(Clk), .RN(Rst), 
        .Q(n106826) );
  DFFR_X2 \DLX_Datapath/PC_reg[30]  ( .D(n60295), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0 [2]), .QN(n57430) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[28]  ( .D(n106521), .CK(Clk), .RN(Rst), 
        .Q(n106827) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[29]  ( .D(n106520), .CK(Clk), .RN(Rst), 
        .Q(n106828) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[29]  ( .D(n106641), .CK(Clk), .RN(Rst), 
        .Q(n69303) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[29]  ( .D(n59078), .CK(Clk), .RN(Rst), 
        .Q(n106830), .QN(n61904) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26856 ), .CK(Clk), .RN(Rst), .Q(n106838), 
        .QN(n103327) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[29]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n106836), .Q(
        \DLX_Datapath/next_B_IDEX [29]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[29]  ( .D(n106687), .CK(Clk), .RN(Rst), .Q(
        n69307), .QN(n104669) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[29]  ( .D(n106839), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [29]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[29]  ( .D(n104327), .CK(Clk), .RN(Rst), .Q(DataAddr[29]), .QN(n58724) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[11]  ( .D(n103931), .CK(Clk), .RN(Rst), 
        .Q(n106842) );
  DFFS_X2 \DLX_Datapath/IR_IFID_reg[30]  ( .D(n60366), .CK(Clk), .SN(n106508), 
        .Q(n69313), .QN(n106847) );
  DFFS_X2 \DLX_Datapath/IR_IDEX_reg[30]  ( .D(\DLX_Datapath/N357 ), .CK(Clk), 
        .SN(Rst), .Q(n69315) );
  DFFS_X2 \DLX_Datapath/IR_MEMWB_reg[30]  ( .D(n111022), .CK(Clk), .SN(n106508), .Q(n69319), .QN(n104443) );
  DFFS_X2 \DLX_Datapath/IR_IFID_reg[28]  ( .D(n60367), .CK(Clk), .SN(Rst), .Q(
        n69321), .QN(n106936) );
  DFFS_X2 \DLX_Datapath/IR_IDEX_reg[28]  ( .D(\DLX_Datapath/N355 ), .CK(Clk), 
        .SN(n106508), .Q(n69322), .QN(n106937) );
  DFFS_X2 \DLX_Datapath/IR_EXMEM_reg[28]  ( .D(n69322), .CK(Clk), .SN(Rst), 
        .Q(n69323), .QN(n106940) );
  DFFS_X2 \DLX_Datapath/IR_MEMWB_reg[28]  ( .D(n69323), .CK(Clk), .SN(n106508), 
        .Q(n69324), .QN(n104442) );
  DFFS_X2 \DLX_Datapath/IR_IFID_reg[26]  ( .D(n60368), .CK(Clk), .SN(Rst), .Q(
        n69325), .QN(n106942) );
  DFFS_X2 \DLX_Datapath/IR_IDEX_reg[26]  ( .D(\DLX_Datapath/N353 ), .CK(Clk), 
        .SN(n106508), .Q(n69326), .QN(n104427) );
  DFFS_X2 \DLX_Datapath/IR_EXMEM_reg[26]  ( .D(n69326), .CK(Clk), .SN(Rst), 
        .Q(n106943), .QN(n57378) );
  DFFS_X2 \DLX_Datapath/IR_MEMWB_reg[26]  ( .D(n106943), .CK(Clk), .SN(Rst), 
        .Q(n106944), .QN(n100762) );
  DFFR_X2 \DLX_ControlUnit/ALUop2_reg[4]  ( .D(n106554), .CK(Clk), .RN(Rst), 
        .Q(\DLX_ControlUnit/ALUop2 [4]) );
  DFFR_X2 \DLX_ControlUnit/ALUop2_reg[3]  ( .D(n60327), .CK(Clk), .RN(Rst), 
        .Q(\DLX_ControlUnit/ALUop2 [3]) );
  DFFR_X2 \DLX_Datapath/RegisterFile/SWP_reg[0]  ( .D(n60371), .CK(Clk), .RN(
        Rst), .Q(n107027), .QN(\dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ) );
  DFFR_X2 \DLX_Datapath/RegisterFile/CWP_reg[0]  ( .D(n60374), .CK(Clk), .RN(
        Rst), .Q(n105044), .QN(n59516) );
  DFF_X2 \DLX_Datapath/CWP_EXMEM_reg[0]  ( .D(n59073), .CK(Clk), .Q(n69346), 
        .QN(n107104) );
  DFF_X2 \DLX_Datapath/CWP_MEMWB_reg[0]  ( .D(n59072), .CK(Clk), .Q(n107105), 
        .QN(n58722) );
  DFFR_X2 \DLX_Datapath/RegisterFile/CWP_reg[1]  ( .D(n60373), .CK(Clk), .RN(
        Rst), .Q(\DLX_Datapath/CWP_IDEX[1] ), .QN(n59517) );
  DFF_X2 \DLX_Datapath/CWP_EXMEM_reg[1]  ( .D(n59071), .CK(Clk), .Q(n69347), 
        .QN(n104950) );
  DFF_X2 \DLX_Datapath/CWP_MEMWB_reg[1]  ( .D(n59070), .CK(Clk), .Q(n107107), 
        .QN(n58720) );
  DFFR_X2 \DLX_Datapath/RegisterFile/CWP_reg[2]  ( .D(n60372), .CK(Clk), .RN(
        Rst), .Q(\DLX_Datapath/CWP_IDEX[2] ), .QN(n59518) );
  DFF_X2 \DLX_Datapath/CWP_MEMWB_reg[2]  ( .D(n59068), .CK(Clk), .QN(n107109)
         );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[0]  ( .D(n106571), .CK(Clk), .RN(Rst), .Q(
        n69349), .QN(n104564) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[1]  ( .D(n106594), .CK(Clk), .RN(Rst), .Q(
        n69350), .QN(n104563) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[3]  ( .D(n106592), .CK(Clk), .RN(Rst), .Q(
        n69352), .QN(n104562) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[4]  ( .D(n106570), .CK(Clk), .RN(Rst), .Q(
        n69353), .QN(n104561) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[5]  ( .D(n106569), .CK(Clk), .RN(Rst), .Q(
        n69354), .QN(n104560) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[7]  ( .D(n106578), .CK(Clk), .RN(Rst), .Q(
        n69356), .QN(n104559) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[9]  ( .D(n106567), .CK(Clk), .RN(Rst), .Q(
        n69358), .QN(n104558) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[10]  ( .D(n106577), .CK(Clk), .RN(Rst), 
        .Q(n69359), .QN(n104557) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[11]  ( .D(n106591), .CK(Clk), .RN(Rst), 
        .Q(\DLX_Datapath/IR_IFID[11] ), .QN(n57380) );
  SDFFR_X2 \DLX_Datapath/IR_IDEX_reg[11]  ( .D(1'b0), .SI(net113091), .SE(
        \DLX_Datapath/IR_IFID[11] ), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/HazardDetUnit/N109 ), .QN(n100424) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[11]  ( .D(
        \DLX_Datapath/HazardDetUnit/N137 ), .CK(Clk), .RN(Rst), .QN(n54614) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[12]  ( .D(n106576), .CK(Clk), .RN(Rst), 
        .Q(\DLX_Datapath/IR_IFID[12] ), .QN(n57381) );
  SDFFR_X2 \DLX_Datapath/IR_IDEX_reg[12]  ( .D(1'b0), .SI(net113102), .SE(
        \DLX_Datapath/IR_IFID[12] ), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/HazardDetUnit/N110 ), .QN(n100426) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[12]  ( .D(
        \DLX_Datapath/HazardDetUnit/N138 ), .CK(Clk), .RN(Rst), .QN(n54616) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[13]  ( .D(n106566), .CK(Clk), .RN(Rst), 
        .Q(\DLX_Datapath/IR_IFID[13] ), .QN(n57382) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[13]  ( .D(
        \DLX_Datapath/HazardDetUnit/N139 ), .CK(Clk), .RN(Rst), .QN(n54618) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[14]  ( .D(n106590), .CK(Clk), .RN(Rst), 
        .Q(n69362), .QN(n104501) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[14]  ( .D(
        \DLX_Datapath/HazardDetUnit/N112 ), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/HazardDetUnit/N140 ), .QN(n62662) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[14]  ( .D(
        \DLX_Datapath/HazardDetUnit/N140 ), .CK(Clk), .RN(Rst), .Q(n107129), 
        .QN(n100894) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[15]  ( .D(\DLX_Datapath/IR_IDEX[15] ), 
        .CK(Clk), .RN(Rst), .Q(\DLX_Datapath/IR_EXMEM[15] ), .QN(n62661) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[15]  ( .D(\DLX_Datapath/IR_EXMEM[15] ), 
        .CK(Clk), .RN(Rst), .Q(n104497), .QN(n54623) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[16]  ( .D(n106588), .CK(Clk), .RN(Rst), 
        .Q(n107132), .QN(n59435) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[16]  ( .D(\DLX_Datapath/N343 ), .CK(Clk), 
        .RN(Rst), .Q(\DLX_Datapath/HazardDetUnit/N95 ), .QN(n62496) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[16]  ( .D(
        \DLX_Datapath/HazardDetUnit/N123 ), .CK(Clk), .RN(Rst), .Q(n107133), 
        .QN(n100632) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[17]  ( .D(n106587), .CK(Clk), .RN(Rst), 
        .Q(n107134), .QN(n59441) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[17]  ( .D(
        \DLX_Datapath/HazardDetUnit/N124 ), .CK(Clk), .RN(Rst), .Q(n107135), 
        .QN(n100631) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[18]  ( .D(n106565), .CK(Clk), .RN(Rst), 
        .Q(n107137), .QN(n59442) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[18]  ( .D(
        \DLX_Datapath/HazardDetUnit/N125 ), .CK(Clk), .RN(Rst), .Q(n107138), 
        .QN(n100630) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[19]  ( .D(n106586), .CK(Clk), .RN(Rst), 
        .Q(n107139), .QN(n59443) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[19]  ( .D(\DLX_Datapath/N346 ), .CK(Clk), 
        .RN(Rst), .Q(\DLX_Datapath/HazardDetUnit/N98 ), .QN(n64247) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[19]  ( .D(
        \DLX_Datapath/HazardDetUnit/N98 ), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/HazardDetUnit/N126 ), .QN(n64267) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[19]  ( .D(
        \DLX_Datapath/HazardDetUnit/N126 ), .CK(Clk), .RN(Rst), .Q(n105037), 
        .QN(n54620) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[20]  ( .D(n106564), .CK(Clk), .RN(Rst), 
        .Q(n107142), .QN(n59444) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[20]  ( .D(\DLX_Datapath/N347 ), .CK(Clk), 
        .RN(n106434), .Q(\DLX_Datapath/IR_IDEX[20] ), .QN(n64246) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[20]  ( .D(\DLX_Datapath/IR_IDEX[20] ), 
        .CK(Clk), .RN(n106434), .Q(\DLX_Datapath/IR_EXMEM[20] ), .QN(n64266)
         );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[20]  ( .D(\DLX_Datapath/IR_EXMEM[20] ), 
        .CK(Clk), .RN(n106434), .Q(n107143), .QN(n100892) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[21]  ( .D(n106563), .CK(Clk), .RN(n106434), 
        .Q(n107144), .QN(n59445) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[22]  ( .D(n106562), .CK(Clk), .RN(n106434), 
        .Q(n107145), .QN(n59451) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[23]  ( .D(n106561), .CK(Clk), .RN(n106434), 
        .Q(n105061), .QN(n59452) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[24]  ( .D(n106585), .CK(Clk), .RN(n106434), 
        .Q(n104707), .QN(n59453) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[25]  ( .D(n106575), .CK(Clk), .RN(n106434), 
        .Q(n104495), .QN(n59454) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[27]  ( .D(n106584), .CK(Clk), .RN(n106434), 
        .Q(n69377), .QN(n104496) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[27]  ( .D(\DLX_Datapath/N354 ), .CK(Clk), 
        .RN(n106434), .Q(\DLX_Datapath/IR_IDEX[27] ), .QN(n59415) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[27]  ( .D(\DLX_Datapath/IR_IDEX[27] ), 
        .CK(Clk), .RN(n106434), .Q(\DLX_Datapath/IR_EXMEM[27] ), .QN(n59323)
         );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[29]  ( .D(n106583), .CK(Clk), .RN(n106483), 
        .Q(n69379), .QN(n104498) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[29]  ( .D(\DLX_Datapath/N356 ), .CK(Clk), 
        .RN(n106430), .Q(\DLX_Datapath/IR_IDEX[29] ), .QN(n59417) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[29]  ( .D(\DLX_Datapath/IR_IDEX[29] ), 
        .CK(Clk), .RN(Rst), .Q(\DLX_Datapath/IR_EXMEM[29] ), .QN(n59325) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[25][0]  ( .D(n60212), 
        .CK(Clk), .RN(n106479), .Q(n107150) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[31]  ( .D(\DLX_Datapath/N358 ), .CK(Clk), 
        .RN(Rst), .Q(\DLX_Datapath/IR_IDEX[31] ), .QN(n59419) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[31]  ( .D(n106662), .CK(Clk), .RN(n106482), .Q(n69413) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[30]  ( .D(n106661), .CK(Clk), .RN(n106505), .Q(n69414) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[28]  ( .D(n106652), .CK(Clk), .RN(n106507), .Q(n69415) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[23]  ( .D(n106639), .CK(Clk), .RN(n106423), .Q(n69416) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[19]  ( .D(n106658), .CK(Clk), .RN(n106489), .Q(n69417) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[31]  ( .D(n59061), .CK(Clk), .RN(Rst), 
        .Q(n107152), .QN(n100794) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[30]  ( .D(n59060), .CK(Clk), .RN(Rst), 
        .Q(n107153), .QN(n100800) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[28]  ( .D(n59059), .CK(Clk), .RN(Rst), 
        .Q(n107154), .QN(n58713) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[23]  ( .D(n59058), .CK(Clk), .RN(Rst), 
        .Q(n107156), .QN(n59346) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[19]  ( .D(n59057), .CK(Clk), .RN(Rst), 
        .Q(n107161), .QN(n59342) );
  DFFR_X2 \DLX_ControlUnit/cw5_reg[3]  ( .D(\DLX_ControlUnit/cw4 [3]), .CK(Clk), .RN(Rst), .QN(n105059) );
  DFFR_X2 \DLX_ControlUnit/cw5_reg[2]  ( .D(\DLX_ControlUnit/cw4 [2]), .CK(Clk), .RN(Rst), .Q(n105048), .QN(n105060) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[4]  ( .D(n103930), .CK(Clk), .RN(Rst), .QN(
        n100770) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][29]  ( .D(n106834), 
        .CK(Clk), .RN(Rst), .Q(n107168), .QN(n102150) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][0]  ( .D(n106990), 
        .CK(Clk), .RN(Rst), .Q(n107169), .QN(n101666) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26760 ), .CK(Clk), .RN(Rst), .Q(n69429), 
        .QN(n104554) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26731 ), .CK(Clk), .RN(Rst), .Q(n69430), 
        .QN(n104528) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26728 ), .CK(Clk), .RN(Rst), .Q(n107170), 
        .QN(n103326) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26699 ), .CK(Clk), .RN(Rst), .Q(n107171), 
        .QN(n102766) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26696 ), .CK(Clk), .RN(Rst), .Q(n107172), 
        .QN(n102718) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26667 ), .CK(Clk), .RN(Rst), .Q(n107173), 
        .QN(n102199) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][29]  ( .D(n106833), 
        .CK(Clk), .RN(Rst), .Q(n107174) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][0]  ( .D(n106959), 
        .CK(Clk), .RN(Rst), .Q(n107175) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26632 ), .CK(Clk), .RN(Rst), .Q(n107176)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26603 ), .CK(Clk), .RN(Rst), .Q(n107177)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26600 ), .CK(Clk), .RN(Rst), .Q(n107178)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26571 ), .CK(Clk), .RN(Rst), .Q(n107179)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26539 ), .CK(Clk), .RN(Rst), .Q(n107181)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26536 ), .CK(Clk), .RN(Rst), .Q(n107182)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26507 ), .CK(Clk), .RN(Rst), .Q(n107183)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26504 ), .CK(Clk), .RN(Rst), .Q(n107184), 
        .QN(n103886) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26475 ), .CK(Clk), .RN(Rst), .Q(n107185), 
        .QN(n103369) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26472 ), .CK(Clk), .RN(Rst), .Q(n107186)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26443 ), .CK(Clk), .RN(Rst), .Q(n107187)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26440 ), .CK(Clk), .RN(Rst), .Q(n107188)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26408 ), .CK(Clk), .RN(Rst), .Q(n107190)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26379 ), .CK(Clk), .RN(Rst), .Q(n107191)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26376 ), .CK(Clk), .RN(Rst), .Q(n107192)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26347 ), .CK(Clk), .RN(Rst), .Q(n107193)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26344 ), .CK(Clk), .RN(Rst), .Q(n107194)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26315 ), .CK(Clk), .RN(Rst), .Q(n107195)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26312 ), .CK(Clk), .RN(Rst), .Q(n107196)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26283 ), .CK(Clk), .RN(Rst), .Q(n107197)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26280 ), .CK(Clk), .RN(Rst), .Q(n69459) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26251 ), .CK(Clk), .RN(Rst), .Q(n69460) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26248 ), .CK(Clk), .RN(Rst), .Q(n107198)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26219 ), .CK(Clk), .RN(Rst), .Q(n107199)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26216 ), .CK(Clk), .RN(Rst), .Q(n69463) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26187 ), .CK(Clk), .RN(n106433), .Q(n69464) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][29]  ( .D(n104244), 
        .CK(Clk), .RN(n106433), .Q(n69465) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26155 ), .CK(Clk), .RN(n106433), .Q(n69466) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26152 ), .CK(Clk), .RN(n106433), .Q(
        n107200), .QN(n102149) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26123 ), .CK(Clk), .RN(n106433), .Q(
        n107201), .QN(n101665) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26091 ), .CK(Clk), .RN(n106433), .Q(n69470) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26088 ), .CK(Clk), .RN(n106433), .Q(
        n107202) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26059 ), .CK(Clk), .RN(n106433), .Q(
        n107203) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26056 ), .CK(Clk), .RN(n106433), .Q(
        n107204) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][0]  ( .D(n104232), 
        .CK(Clk), .RN(n106433), .Q(n107205) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26024 ), .CK(Clk), .RN(n106433), .Q(
        n107206) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25995 ), .CK(Clk), .RN(n106434), .Q(
        n107207) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25992 ), .CK(Clk), .RN(n106436), .Q(
        n107208), .QN(n103885) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25963 ), .CK(Clk), .RN(n106436), .Q(
        n107209), .QN(n103367) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25960 ), .CK(Clk), .RN(n106436), .Q(
        n107210) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25931 ), .CK(Clk), .RN(n106436), .Q(
        n107211) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][29]  ( .D(n104265), 
        .CK(Clk), .RN(n106436), .Q(n107212) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][0]  ( .D(n104259), 
        .CK(Clk), .RN(n106436), .Q(n107213) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25896 ), .CK(Clk), .RN(n106436), .Q(n69483) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25867 ), .CK(Clk), .RN(n106436), .Q(n69484) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25864 ), .CK(Clk), .RN(n106436), .Q(n69486) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25832 ), .CK(Clk), .RN(n106436), .Q(
        n107214) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25800 ), .CK(Clk), .RN(n106441), .Q(
        n107215) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25768 ), .CK(Clk), .RN(n106482), .Q(
        n107216) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25704 ), .CK(Clk), .RN(Rst), .Q(n107217)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25640 ), .CK(Clk), .RN(n106485), .Q(
        n107218) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25608 ), .CK(Clk), .RN(n106484), .Q(
        n107219) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25576 ), .CK(Clk), .RN(n106483), .Q(
        n107220) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25544 ), .CK(Clk), .RN(n106442), .Q(
        n107221) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25512 ), .CK(Clk), .RN(Rst), .Q(n107222), 
        .QN(n100563) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25480 ), .CK(Clk), .RN(Rst), .Q(n69498) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25448 ), .CK(Clk), .RN(Rst), .Q(n107223)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25416 ), .CK(Clk), .RN(n106439), .Q(
        n107224) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25384 ), .CK(Clk), .RN(Rst), .Q(n107225)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][29]  ( .D(n104309), 
        .CK(Clk), .RN(n106456), .Q(n107226) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25288 ), .CK(Clk), .RN(n106399), .Q(
        n107228), .QN(n102716) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25256 ), .CK(Clk), .RN(n106371), .Q(
        n107229), .QN(n102145) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25224 ), .CK(Clk), .RN(Rst), .Q(n107230)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25192 ), .CK(Clk), .RN(Rst), .Q(n69507) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25160 ), .CK(Clk), .RN(Rst), .Q(n107231)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][29]  ( .D(n104283), 
        .CK(Clk), .RN(Rst), .Q(n107232) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25064 ), .CK(Clk), .RN(n106383), .Q(n69511), .QN(n104613) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][29]  ( .D(n104206), 
        .CK(Clk), .RN(n106430), .Q(n107233) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25000 ), .CK(Clk), .RN(Rst), .Q(n107234), 
        .QN(n100595) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24968 ), .CK(Clk), .RN(Rst), .Q(n69514) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24936 ), .CK(Clk), .RN(Rst), .Q(n69515) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24904 ), .CK(Clk), .RN(Rst), .Q(n107235), 
        .QN(n101151) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24872 ), .CK(Clk), .RN(Rst), .Q(n107236)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24840 ), .CK(Clk), .RN(Rst), .Q(n107237)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24808 ), .CK(Clk), .RN(Rst), .Q(n69519) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24776 ), .CK(Clk), .RN(Rst), .Q(n107238)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24712 ), .CK(Clk), .RN(Rst), .Q(n107239)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24680 ), .CK(Clk), .RN(Rst), .Q(n107240), 
        .QN(n103320) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24648 ), .CK(Clk), .RN(n106464), .Q(n69524) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24616 ), .CK(Clk), .RN(n106463), .Q(
        n107241) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24552 ), .CK(Clk), .RN(n106462), .Q(
        n107242) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24520 ), .CK(Clk), .RN(Rst), .Q(n107243), 
        .QN(n102710) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24488 ), .CK(Clk), .RN(n106487), .Q(n69529), .QN(n104634) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24456 ), .CK(Clk), .RN(Rst), .Q(n107244)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24424 ), .CK(Clk), .RN(Rst), .Q(n107245)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24392 ), .CK(Clk), .RN(Rst), .Q(n107246)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24360 ), .CK(Clk), .RN(n106436), .Q(
        n107247) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24328 ), .CK(Clk), .RN(n106474), .Q(
        n107248) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24296 ), .CK(Clk), .RN(n106396), .Q(
        n107249), .QN(n103318) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24264 ), .CK(Clk), .RN(Rst), .Q(n107250)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24232 ), .CK(Clk), .RN(n106493), .Q(
        n107251) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24168 ), .CK(Clk), .RN(Rst), .Q(n107252)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24136 ), .CK(Clk), .RN(Rst), .Q(n107253)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24072 ), .CK(Clk), .RN(n106398), .Q(
        n107254) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24040 ), .CK(Clk), .RN(Rst), .Q(n69543) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24008 ), .CK(Clk), .RN(Rst), .Q(n107255), 
        .QN(n102708) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23976 ), .CK(Clk), .RN(Rst), .Q(n69545) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23944 ), .CK(Clk), .RN(Rst), .Q(n107256), 
        .QN(n103878) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23912 ), .CK(Clk), .RN(n106494), .Q(
        n107257), .QN(n103316) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23880 ), .CK(Clk), .RN(n106456), .Q(
        n107258) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23816 ), .CK(Clk), .RN(n106441), .Q(
        n107259) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23784 ), .CK(Clk), .RN(Rst), .Q(n107260), 
        .QN(n101023) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][29]  ( .D(n104041), 
        .CK(Clk), .RN(n106487), .Q(n107261) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23720 ), .CK(Clk), .RN(n106487), .Q(n69553) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23688 ), .CK(Clk), .RN(n106490), .Q(
        n107262), .QN(n100994) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23656 ), .CK(Clk), .RN(Rst), .Q(n69555) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23624 ), .CK(Clk), .RN(Rst), .Q(n107263)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23592 ), .CK(Clk), .RN(Rst), .Q(n107264)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23560 ), .CK(Clk), .RN(n106395), .Q(
        n107265), .QN(n103874) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23528 ), .CK(Clk), .RN(n106435), .Q(
        n107266) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23496 ), .CK(Clk), .RN(n106435), .Q(n69560) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23464 ), .CK(Clk), .RN(n106435), .Q(n69561) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23432 ), .CK(Clk), .RN(n106435), .Q(
        n107267) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23400 ), .CK(Clk), .RN(n106435), .Q(
        n107268) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23368 ), .CK(Clk), .RN(n106435), .Q(n69564) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23336 ), .CK(Clk), .RN(n106435), .Q(
        n107269) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23304 ), .CK(Clk), .RN(n106435), .Q(
        n107270) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23240 ), .CK(Clk), .RN(n106435), .Q(
        n107272) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23208 ), .CK(Clk), .RN(n106435), .Q(
        n107273) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23176 ), .CK(Clk), .RN(n106435), .Q(
        n107274) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23112 ), .CK(Clk), .RN(Rst), .Q(n107275)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23080 ), .CK(Clk), .RN(Rst), .Q(n107276)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23048 ), .CK(Clk), .RN(Rst), .Q(n107277)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23016 ), .CK(Clk), .RN(Rst), .Q(n107278)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22984 ), .CK(Clk), .RN(Rst), .Q(n107279)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22952 ), .CK(Clk), .RN(n106507), .Q(n69577) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22920 ), .CK(Clk), .RN(Rst), .Q(n69578) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22888 ), .CK(Clk), .RN(n106464), .Q(
        n107280) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22856 ), .CK(Clk), .RN(Rst), .Q(n107281)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22824 ), .CK(Clk), .RN(Rst), .Q(n69581) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22792 ), .CK(Clk), .RN(Rst), .Q(n107282)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22760 ), .CK(Clk), .RN(Rst), .Q(n69583) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22728 ), .CK(Clk), .RN(Rst), .Q(n107283)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22696 ), .CK(Clk), .RN(Rst), .Q(n107284)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22664 ), .CK(Clk), .RN(Rst), .Q(n107285)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22632 ), .CK(Clk), .RN(Rst), .Q(n107286)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22600 ), .CK(Clk), .RN(Rst), .Q(n69588) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25835 ), .CK(Clk), .RN(Rst), .Q(n69591) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25803 ), .CK(Clk), .RN(Rst), .Q(n107288)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25771 ), .CK(Clk), .RN(Rst), .Q(n107289)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25739 ), .CK(Clk), .RN(Rst), .Q(n107290)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25675 ), .CK(Clk), .RN(Rst), .Q(n107291)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25611 ), .CK(Clk), .RN(Rst), .Q(n107292)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25579 ), .CK(Clk), .RN(Rst), .Q(n107293)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25547 ), .CK(Clk), .RN(Rst), .Q(n107294)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25515 ), .CK(Clk), .RN(Rst), .Q(n107295)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25483 ), .CK(Clk), .RN(Rst), .Q(n107296), 
        .QN(n100592) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25451 ), .CK(Clk), .RN(Rst), .Q(n69603) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25419 ), .CK(Clk), .RN(Rst), .Q(n107297)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25387 ), .CK(Clk), .RN(Rst), .Q(n107298)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25355 ), .CK(Clk), .RN(Rst), .Q(n107299)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25323 ), .CK(Clk), .RN(Rst), .Q(n107300)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25291 ), .CK(Clk), .RN(Rst), .Q(n107301), 
        .QN(n102763) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25259 ), .CK(Clk), .RN(Rst), .Q(n107302), 
        .QN(n102197) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25227 ), .CK(Clk), .RN(Rst), .Q(n107303), 
        .QN(n101661) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25195 ), .CK(Clk), .RN(Rst), .Q(n107304)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25163 ), .CK(Clk), .RN(Rst), .Q(n69612) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25131 ), .CK(Clk), .RN(Rst), .Q(n107305)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25067 ), .CK(Clk), .RN(Rst), .Q(n107306)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25035 ), .CK(Clk), .RN(Rst), .Q(n69616), 
        .QN(n104584) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25003 ), .CK(Clk), .RN(Rst), .Q(n107307)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24971 ), .CK(Clk), .RN(Rst), .Q(n107308), 
        .QN(n100624) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24939 ), .CK(Clk), .RN(Rst), .Q(n107309)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24907 ), .CK(Clk), .RN(Rst), .Q(n69620) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24875 ), .CK(Clk), .RN(Rst), .Q(n107310), 
        .QN(n101179) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24843 ), .CK(Clk), .RN(Rst), .Q(n107311)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24811 ), .CK(Clk), .RN(Rst), .Q(n107312)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24779 ), .CK(Clk), .RN(Rst), .Q(n69624) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24747 ), .CK(Clk), .RN(Rst), .Q(n107313)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24683 ), .CK(Clk), .RN(Rst), .Q(n107314)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24651 ), .CK(Clk), .RN(Rst), .Q(n107315), 
        .QN(n102759) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24619 ), .CK(Clk), .RN(Rst), .Q(n69629) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24587 ), .CK(Clk), .RN(Rst), .Q(n107316)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24523 ), .CK(Clk), .RN(Rst), .Q(n107317)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24491 ), .CK(Clk), .RN(Rst), .Q(n107318), 
        .QN(n102190) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24459 ), .CK(Clk), .RN(Rst), .Q(n69634), 
        .QN(n104637) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24427 ), .CK(Clk), .RN(Rst), .Q(n107319)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24395 ), .CK(Clk), .RN(Rst), .Q(n107320)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24363 ), .CK(Clk), .RN(Rst), .Q(n107321)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24331 ), .CK(Clk), .RN(Rst), .Q(n107322)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24299 ), .CK(Clk), .RN(Rst), .Q(n107323)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24267 ), .CK(Clk), .RN(Rst), .Q(n107324), 
        .QN(n102756) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24235 ), .CK(Clk), .RN(Rst), .Q(n107325)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24203 ), .CK(Clk), .RN(Rst), .Q(n107326)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24139 ), .CK(Clk), .RN(Rst), .Q(n107327)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24107 ), .CK(Clk), .RN(Rst), .Q(n107328)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24043 ), .CK(Clk), .RN(Rst), .Q(n107329)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24011 ), .CK(Clk), .RN(Rst), .Q(n69648) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23979 ), .CK(Clk), .RN(Rst), .Q(n107330), 
        .QN(n102188) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23947 ), .CK(Clk), .RN(Rst), .Q(n107331)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23915 ), .CK(Clk), .RN(Rst), .Q(n107332), 
        .QN(n103358) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23883 ), .CK(Clk), .RN(Rst), .Q(n107333), 
        .QN(n102754) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23851 ), .CK(Clk), .RN(Rst), .Q(n107334)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23787 ), .CK(Clk), .RN(Rst), .Q(n107335)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23755 ), .CK(Clk), .RN(Rst), .Q(n107336), 
        .QN(n101052) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23723 ), .CK(Clk), .RN(Rst), .Q(n107337)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23691 ), .CK(Clk), .RN(Rst), .Q(n69658) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23659 ), .CK(Clk), .RN(Rst), .Q(n107338), 
        .QN(n101020) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23627 ), .CK(Clk), .RN(Rst), .Q(n69660) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23595 ), .CK(Clk), .RN(Rst), .Q(n107339)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23563 ), .CK(Clk), .RN(Rst), .Q(n107340)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23531 ), .CK(Clk), .RN(Rst), .Q(n107341), 
        .QN(n103354) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23499 ), .CK(Clk), .RN(Rst), .Q(n107342)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23467 ), .CK(Clk), .RN(Rst), .Q(n69665) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23435 ), .CK(Clk), .RN(Rst), .Q(n69666) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23403 ), .CK(Clk), .RN(Rst), .Q(n107343)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23371 ), .CK(Clk), .RN(Rst), .Q(n107344)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23339 ), .CK(Clk), .RN(Rst), .Q(n107345)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23307 ), .CK(Clk), .RN(Rst), .Q(n107346)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23275 ), .CK(Clk), .RN(Rst), .Q(n107347)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23243 ), .CK(Clk), .RN(Rst), .Q(n107348), 
        .QN(n102752) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23211 ), .CK(Clk), .RN(Rst), .Q(n107349)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23179 ), .CK(Clk), .RN(Rst), .Q(n107350)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23147 ), .CK(Clk), .RN(Rst), .Q(n107351)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23115 ), .CK(Clk), .RN(Rst), .Q(n107352)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23083 ), .CK(Clk), .RN(Rst), .Q(n107353)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23051 ), .CK(Clk), .RN(Rst), .Q(n107354)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][0]  ( .D(n103990), 
        .CK(Clk), .RN(Rst), .Q(n107355) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22987 ), .CK(Clk), .RN(Rst), .Q(n107356)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][0]  ( .D(n104012), 
        .CK(Clk), .RN(Rst), .Q(n107357) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22923 ), .CK(Clk), .RN(Rst), .Q(n69682) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][0]  ( .D(n103993), 
        .CK(Clk), .RN(Rst), .Q(n69683) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22859 ), .CK(Clk), .RN(Rst), .Q(n107358)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22827 ), .CK(Clk), .RN(Rst), .Q(n107359)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22795 ), .CK(Clk), .RN(Rst), .Q(n107360)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22763 ), .CK(Clk), .RN(Rst), .Q(n107361)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22731 ), .CK(Clk), .RN(Rst), .Q(n69688) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22667 ), .CK(Clk), .RN(Rst), .Q(n107362)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22635 ), .CK(Clk), .RN(Rst), .Q(n107363)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22603 ), .CK(Clk), .RN(Rst), .Q(n107364)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22571 ), .CK(Clk), .RN(Rst), .Q(n107365)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22539 ), .CK(Clk), .RN(Rst), .Q(n69694), 
        .QN(n104512) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[11]  ( .D(n59093), .CK(Clk), .RN(n106430), 
        .Q(\DLX_ControlUnit/cw2 [11]), .QN(n57390) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[29]  ( .D(n59013), .CK(Clk), .RN(n106430), 
        .Q(n107414) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[0]  ( .D(n59012), .CK(Clk), .RN(n106430), 
        .Q(n107415) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[16]  ( .D(n62245), .CK(Clk), .RN(n106430), 
        .QN(n62247) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[17]  ( .D(n59084), .CK(Clk), .RN(n106430), 
        .Q(\DLX_ControlUnit/cw2 [17]), .QN(n57393) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[20]  ( .D(n106558), .CK(Clk), .RN(n106430), 
        .Q(n107417) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[21]  ( .D(n106572), .CK(Clk), .RN(Rst), .Q(
        n104506), .QN(n100463) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[0]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(
        \DLX_Datapath/RegisterFile/N46424 ), .Q(\DLX_Datapath/next_A_IDEX[0] )
         );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[0]  ( .D(n106599), .CK(Clk), .RN(Rst), .Q(
        n107419) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[29]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n106835), .Q(
        \DLX_Datapath/next_A_IDEX[29] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[29]  ( .D(n106629), .CK(Clk), .RN(Rst), .Q(
        n107420) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[10]  ( .D(n60346), .CK(Clk), .RN(Rst), 
        .QN(n100638) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[9]  ( .D(n60347), .CK(Clk), .RN(Rst), 
        .QN(n100639) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[8]  ( .D(n60348), .CK(Clk), .RN(Rst), 
        .QN(n100640) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[7]  ( .D(n60349), .CK(Clk), .RN(Rst), 
        .QN(n100641) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[6]  ( .D(n60350), .CK(Clk), .RN(Rst), 
        .QN(n100642) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[5]  ( .D(n60351), .CK(Clk), .RN(Rst), 
        .QN(n100643) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[4]  ( .D(n60352), .CK(Clk), .RN(Rst), 
        .QN(n100644) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[3]  ( .D(n60353), .CK(Clk), .RN(Rst), 
        .QN(n100645) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[2]  ( .D(n60354), .CK(Clk), .RN(Rst), 
        .QN(n100646) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[1]  ( .D(n60355), .CK(Clk), .RN(Rst), 
        .QN(n100647) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[0]  ( .D(n60356), .CK(Clk), .RN(Rst), 
        .QN(n100648) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[15]  ( .D(n59220), .CK(Clk), .RN(Rst), 
        .QN(n100633) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[14]  ( .D(n59219), .CK(Clk), .RN(Rst), 
        .QN(n100634) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[13]  ( .D(n59218), .CK(Clk), .RN(Rst), 
        .QN(n100635) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[12]  ( .D(n59217), .CK(Clk), .RN(Rst), 
        .QN(n100636) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[11]  ( .D(n59216), .CK(Clk), .RN(Rst), 
        .QN(n100637) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[26]  ( .D(n60335), .CK(Clk), .RN(Rst), 
        .Q(n69784), .QN(n104570) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[25]  ( .D(n60336), .CK(Clk), .RN(n106490), 
        .Q(n69785), .QN(n104571) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[24]  ( .D(n60337), .CK(Clk), .RN(Rst), 
        .Q(n69786), .QN(n104572) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[23]  ( .D(n60338), .CK(Clk), .RN(Rst), 
        .Q(n69787), .QN(n104573) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[22]  ( .D(n60339), .CK(Clk), .RN(Rst), 
        .Q(n69788), .QN(n104574) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[21]  ( .D(n60340), .CK(Clk), .RN(Rst), 
        .Q(n69789), .QN(n104575) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[20]  ( .D(n60341), .CK(Clk), .RN(Rst), 
        .Q(n69790), .QN(n104576) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[19]  ( .D(n60342), .CK(Clk), .RN(Rst), 
        .Q(n69791), .QN(n104577) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[18]  ( .D(n60343), .CK(Clk), .RN(Rst), 
        .Q(n69792), .QN(n104578) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[17]  ( .D(n60344), .CK(Clk), .RN(Rst), 
        .Q(n69793), .QN(n104579) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[16]  ( .D(n60345), .CK(Clk), .RN(Rst), 
        .Q(n69794), .QN(n104580) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[31]  ( .D(n60330), .CK(Clk), .RN(n106393), 
        .Q(n69795), .QN(n104565) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[30]  ( .D(n60331), .CK(Clk), .RN(Rst), 
        .Q(n69796), .QN(n104566) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[29]  ( .D(n60332), .CK(Clk), .RN(n106429), 
        .Q(n69797), .QN(n104567) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[28]  ( .D(n60333), .CK(Clk), .RN(n106429), 
        .Q(n69798), .QN(n104568) );
  DFFR_X2 \DLX_Datapath/Imm_IDEX_reg[27]  ( .D(n60334), .CK(Clk), .RN(n106429), 
        .Q(n69799), .QN(n104569) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[0]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [0]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[0]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [0]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [0]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/sel_shf_reg[1]  ( .D(n60443), .GN(n106949), 
        .Q(\DLX_Datapath/ArithLogUnit/sel_shf [1]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/sel_shf_reg[0]  ( .D(n60442), .GN(n105198), 
        .Q(\DLX_Datapath/ArithLogUnit/sel_shf [0]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_shf_reg[0]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [0]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/B_shf [0]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[29]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [29]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [29]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[0]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [0]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [0]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[0]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [0]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [0]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[29]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [29]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [29]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[0]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [0]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [0]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[29]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [29]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [29]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/sel_log_reg[1]  ( .G(n106369), .D(
        \DLX_Datapath/ArithLogUnit/N179 ), .Q(
        \DLX_Datapath/ArithLogUnit/sel_log [1]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/sel_log_reg[2]  ( .G(n106370), .D(
        \DLX_Datapath/ArithLogUnit/N179 ), .Q(
        \DLX_Datapath/ArithLogUnit/sel_log [2]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/sel_log_reg[3]  ( .G(n106369), .D(
        \DLX_Datapath/ArithLogUnit/N180 ), .Q(
        \DLX_Datapath/ArithLogUnit/sel_log [3]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/Cin_add_reg  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N177 ), .Q(\DLX_Datapath/ArithLogUnit/Cin_add ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[0]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N145 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [0]) );
  DFFR_X2 \DLX_Datapath/PC_reg[2]  ( .D(n60323), .CK(Clk), .RN(n106429), .Q(
        n74605), .QN(net2465245) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[11]  ( .D(n106538), .CK(Clk), .RN(n106429), .Q(n107621) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[11]  ( .D(n106635), .CK(Clk), .RN(n106429), .Q(n69991) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[11]  ( .D(n59009), .CK(Clk), .RN(n106429), .Q(n107622), .QN(n59334) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25847 ), .CK(Clk), .RN(n106449), .Q(n69994) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25815 ), .CK(Clk), .RN(n106431), .Q(
        n107632) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25783 ), .CK(Clk), .RN(Rst), .Q(n107633)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25751 ), .CK(Clk), .RN(n106479), .Q(
        n107634) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25687 ), .CK(Clk), .RN(Rst), .Q(n107635)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25623 ), .CK(Clk), .RN(Rst), .Q(n107636)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25591 ), .CK(Clk), .RN(n106489), .Q(
        n107637) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25559 ), .CK(Clk), .RN(n106488), .Q(
        n107638) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25527 ), .CK(Clk), .RN(n106490), .Q(
        n107639) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25495 ), .CK(Clk), .RN(n106410), .Q(
        n107640), .QN(n100580) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25463 ), .CK(Clk), .RN(Rst), .Q(n70006) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25431 ), .CK(Clk), .RN(n106432), .Q(
        n107641) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25399 ), .CK(Clk), .RN(n106432), .Q(
        n107642) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25367 ), .CK(Clk), .RN(n106432), .Q(
        n107643) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25335 ), .CK(Clk), .RN(n106432), .Q(
        n107644) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25303 ), .CK(Clk), .RN(n106432), .Q(
        n107645), .QN(n103000) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25271 ), .CK(Clk), .RN(n106432), .Q(
        n107646), .QN(n102433) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25239 ), .CK(Clk), .RN(n106432), .Q(
        n107647), .QN(n101871) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25207 ), .CK(Clk), .RN(n106432), .Q(
        n107648) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25175 ), .CK(Clk), .RN(n106432), .Q(n70015) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25143 ), .CK(Clk), .RN(n106432), .Q(
        n107649) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25079 ), .CK(Clk), .RN(Rst), .Q(n107650)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25047 ), .CK(Clk), .RN(Rst), .Q(n70019), 
        .QN(n104596) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25015 ), .CK(Clk), .RN(n106465), .Q(
        n107651) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24983 ), .CK(Clk), .RN(Rst), .Q(n107652), 
        .QN(n100612) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24951 ), .CK(Clk), .RN(Rst), .Q(n107653)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24919 ), .CK(Clk), .RN(Rst), .Q(n70023) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24887 ), .CK(Clk), .RN(Rst), .Q(n107654), 
        .QN(n101167) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24855 ), .CK(Clk), .RN(n106425), .Q(
        n107655) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24823 ), .CK(Clk), .RN(n106392), .Q(
        n107656) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24791 ), .CK(Clk), .RN(Rst), .Q(n70027) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24759 ), .CK(Clk), .RN(Rst), .Q(n107657)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24695 ), .CK(Clk), .RN(Rst), .Q(n107658)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24663 ), .CK(Clk), .RN(Rst), .Q(n107659), 
        .QN(n102996) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24631 ), .CK(Clk), .RN(Rst), .Q(n70032) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24599 ), .CK(Clk), .RN(Rst), .Q(n107660)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24535 ), .CK(Clk), .RN(Rst), .Q(n107661)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24503 ), .CK(Clk), .RN(Rst), .Q(n107662), 
        .QN(n102426) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24471 ), .CK(Clk), .RN(Rst), .Q(n70037), 
        .QN(n104617) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24439 ), .CK(Clk), .RN(Rst), .Q(n107663)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24407 ), .CK(Clk), .RN(Rst), .Q(n107664)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24375 ), .CK(Clk), .RN(Rst), .Q(n107665)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24343 ), .CK(Clk), .RN(Rst), .Q(n107666)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24311 ), .CK(Clk), .RN(Rst), .Q(n107667)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24279 ), .CK(Clk), .RN(Rst), .Q(n107668), 
        .QN(n102993) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24247 ), .CK(Clk), .RN(n106508), .Q(
        n107669) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24215 ), .CK(Clk), .RN(n106430), .Q(
        n107670) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24151 ), .CK(Clk), .RN(n106470), .Q(
        n107671) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][12]  ( .D(n104117), 
        .CK(Clk), .RN(n106505), .Q(n107672) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][12]  ( .D(n104080), 
        .CK(Clk), .RN(Rst), .Q(n107673) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24023 ), .CK(Clk), .RN(Rst), .Q(n70051) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23991 ), .CK(Clk), .RN(Rst), .Q(n107674), 
        .QN(n102424) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23959 ), .CK(Clk), .RN(Rst), .Q(n107675)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][12]  ( .D(n104091), 
        .CK(Clk), .RN(n106431), .Q(n107676), .QN(n103587) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23895 ), .CK(Clk), .RN(n106431), .Q(
        n107677), .QN(n102991) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][12]  ( .D(n104129), 
        .CK(Clk), .RN(n106431), .Q(n107678) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23799 ), .CK(Clk), .RN(n106431), .Q(
        n107679) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23767 ), .CK(Clk), .RN(n106431), .Q(
        n107680), .QN(n101040) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23735 ), .CK(Clk), .RN(n106431), .Q(
        n107681) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23703 ), .CK(Clk), .RN(n106431), .Q(n70061) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23671 ), .CK(Clk), .RN(n106431), .Q(
        n107682), .QN(n101009) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23639 ), .CK(Clk), .RN(n106431), .Q(n70063) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23607 ), .CK(Clk), .RN(n106431), .Q(
        n107683) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23575 ), .CK(Clk), .RN(n106431), .Q(
        n107684) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23543 ), .CK(Clk), .RN(Rst), .Q(n107685), 
        .QN(n103583) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23511 ), .CK(Clk), .RN(Rst), .Q(n107686)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23479 ), .CK(Clk), .RN(Rst), .Q(n70068) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23447 ), .CK(Clk), .RN(Rst), .Q(n70069) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23415 ), .CK(Clk), .RN(Rst), .Q(n107687)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23383 ), .CK(Clk), .RN(Rst), .Q(n107688)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23351 ), .CK(Clk), .RN(Rst), .Q(n107689)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23319 ), .CK(Clk), .RN(Rst), .Q(n107690)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23287 ), .CK(Clk), .RN(Rst), .Q(n107691)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23255 ), .CK(Clk), .RN(Rst), .Q(n107692), 
        .QN(n102989) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23223 ), .CK(Clk), .RN(Rst), .Q(n107693)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23191 ), .CK(Clk), .RN(Rst), .Q(n107694)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23159 ), .CK(Clk), .RN(Rst), .Q(n107695)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23127 ), .CK(Clk), .RN(Rst), .Q(n107696)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23095 ), .CK(Clk), .RN(Rst), .Q(n107697)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23063 ), .CK(Clk), .RN(Rst), .Q(n107698)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23031 ), .CK(Clk), .RN(Rst), .Q(n107699)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22999 ), .CK(Clk), .RN(Rst), .Q(n107700)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22967 ), .CK(Clk), .RN(Rst), .Q(n107701)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22935 ), .CK(Clk), .RN(Rst), .Q(n70085) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22903 ), .CK(Clk), .RN(Rst), .Q(n70086) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22871 ), .CK(Clk), .RN(Rst), .Q(n107702)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22839 ), .CK(Clk), .RN(Rst), .Q(n107703)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22807 ), .CK(Clk), .RN(Rst), .Q(n107704)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22775 ), .CK(Clk), .RN(Rst), .Q(n107705)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22743 ), .CK(Clk), .RN(Rst), .Q(n70091) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22711 ), .CK(Clk), .RN(Rst), .Q(n107706)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22679 ), .CK(Clk), .RN(Rst), .Q(n107707)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22647 ), .CK(Clk), .RN(Rst), .Q(n107708)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22615 ), .CK(Clk), .RN(Rst), .Q(n107709)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22583 ), .CK(Clk), .RN(Rst), .Q(n107710)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][12]  ( .D(
        \DLX_Datapath/RegisterFile/N22551 ), .CK(Clk), .RN(Rst), .Q(n70097), 
        .QN(n104523) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25879 ), .CK(Clk), .RN(Rst), .Q(n70098) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][12]  ( .D(n104270), 
        .CK(Clk), .RN(Rst), .Q(n107711) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25943 ), .CK(Clk), .RN(Rst), .Q(n107712)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25975 ), .CK(Clk), .RN(n106417), .Q(
        n107713), .QN(n103595) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26007 ), .CK(Clk), .RN(Rst), .Q(n107714)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][12]  ( .D(n104228), 
        .CK(Clk), .RN(n106493), .Q(n107715) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26071 ), .CK(Clk), .RN(Rst), .Q(n107716)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26103 ), .CK(Clk), .RN(n106372), .Q(n70105) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26135 ), .CK(Clk), .RN(n106506), .Q(
        n107717), .QN(n101875) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26167 ), .CK(Clk), .RN(Rst), .Q(n70107) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26199 ), .CK(Clk), .RN(Rst), .Q(n70108) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26231 ), .CK(Clk), .RN(Rst), .Q(n107718)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26263 ), .CK(Clk), .RN(Rst), .Q(n70110) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][12]  ( .D(n104238), 
        .CK(Clk), .RN(n106504), .Q(n107719) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26327 ), .CK(Clk), .RN(n106372), .Q(
        n107720) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26359 ), .CK(Clk), .RN(Rst), .Q(n107721)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26391 ), .CK(Clk), .RN(Rst), .Q(n107722)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26455 ), .CK(Clk), .RN(Rst), .Q(n107724)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26487 ), .CK(Clk), .RN(Rst), .Q(n107725), 
        .QN(n103597) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26519 ), .CK(Clk), .RN(Rst), .Q(n107726)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26551 ), .CK(Clk), .RN(Rst), .Q(n107727)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26583 ), .CK(Clk), .RN(Rst), .Q(n107728)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26615 ), .CK(Clk), .RN(Rst), .Q(n107729)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][12]  ( .D(n106971), 
        .CK(Clk), .RN(n106505), .Q(n107730) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26679 ), .CK(Clk), .RN(n106507), .Q(
        n107731), .QN(n102435) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26711 ), .CK(Clk), .RN(n106508), .Q(
        n107732), .QN(n103003) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26743 ), .CK(Clk), .RN(Rst), .Q(n70125), 
        .QN(n104537) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][12]  ( .D(n107002), 
        .CK(Clk), .RN(Rst), .Q(n107733), .QN(n101876) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26839 ), .CK(Clk), .RN(Rst), .Q(n107735), 
        .QN(n103004) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[12]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107074), .Q(
        \DLX_Datapath/next_A_IDEX[12] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[12]  ( .D(n106620), .CK(Clk), .RN(Rst), .Q(
        n107736) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[12]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107040), .Q(
        \DLX_Datapath/next_B_IDEX [12]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[12]  ( .D(n106670), .CK(Clk), .RN(Rst), .Q(
        n70130) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[12]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [12]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [12]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[12]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [12]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [12]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[12]  ( .D(n103919), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [12]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[12]  ( .D(n104329), .CK(Clk), .RN(Rst), .Q(DataAddr[12]), .QN(n58698) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[12]  ( .D(n59005), .CK(Clk), .RN(Rst), .Q(
        n107741) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[12]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [12]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[12]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [12]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [12]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[12]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [12]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [12]) );
  DFFR_X2 \DLX_Datapath/PC_reg[12]  ( .D(n60313), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [0]), .QN(n104494) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[18]  ( .D(n103944), .CK(Clk), .RN(Rst), 
        .Q(n107744) );
  DFFR_X2 \DLX_Datapath/PC_reg[18]  ( .D(n60307), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [2]), .QN(n57425) );
  DFFR_X2 \DLX_Datapath/PC_reg[27]  ( .D(n60298), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [3]), .QN(n59478) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[27]  ( .D(n106522), .CK(Clk), .RN(Rst), 
        .Q(n107747) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[27]  ( .D(n106651), .CK(Clk), .RN(Rst), 
        .Q(n70142) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[27]  ( .D(n59004), .CK(Clk), .RN(Rst), 
        .Q(n107748), .QN(n59350) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25863 ), .CK(Clk), .RN(Rst), .Q(n70147) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25831 ), .CK(Clk), .RN(Rst), .Q(n107752)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25799 ), .CK(Clk), .RN(Rst), .Q(n107753)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25767 ), .CK(Clk), .RN(Rst), .Q(n107754)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25703 ), .CK(Clk), .RN(Rst), .Q(n107755)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25639 ), .CK(Clk), .RN(Rst), .Q(n107756)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25607 ), .CK(Clk), .RN(Rst), .Q(n107757), 
        .QN(n103867) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25575 ), .CK(Clk), .RN(Rst), .Q(n107758)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25543 ), .CK(Clk), .RN(Rst), .Q(n107759)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25511 ), .CK(Clk), .RN(Rst), .Q(n107760), 
        .QN(n100564) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25479 ), .CK(Clk), .RN(Rst), .Q(n70159) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25447 ), .CK(Clk), .RN(Rst), .Q(n107761)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25415 ), .CK(Clk), .RN(Rst), .Q(n107762)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25383 ), .CK(Clk), .RN(Rst), .Q(n107763)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][28]  ( .D(n104308), 
        .CK(Clk), .RN(Rst), .Q(n107764) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25319 ), .CK(Clk), .RN(n106432), .Q(
        n107765), .QN(n103307) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25287 ), .CK(Clk), .RN(Rst), .Q(n107766), 
        .QN(n102700) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25255 ), .CK(Clk), .RN(Rst), .Q(n107767), 
        .QN(n102131) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25223 ), .CK(Clk), .RN(Rst), .Q(n107768)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25191 ), .CK(Clk), .RN(Rst), .Q(n70168) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25159 ), .CK(Clk), .RN(Rst), .Q(n107769)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][28]  ( .D(n104282), 
        .CK(Clk), .RN(Rst), .Q(n107770) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25063 ), .CK(Clk), .RN(Rst), .Q(n70172), 
        .QN(n104612) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][28]  ( .D(n104210), 
        .CK(Clk), .RN(Rst), .Q(n107771) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24999 ), .CK(Clk), .RN(Rst), .Q(n107772), 
        .QN(n100596) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][28]  ( .D(n104293), 
        .CK(Clk), .RN(Rst), .Q(n107773) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24935 ), .CK(Clk), .RN(Rst), .Q(n70176) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24903 ), .CK(Clk), .RN(n106502), .Q(
        n107774), .QN(n101152) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24871 ), .CK(Clk), .RN(n106418), .Q(
        n107775) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][28]  ( .D(n104154), 
        .CK(Clk), .RN(n106443), .Q(n107776) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24807 ), .CK(Clk), .RN(n106425), .Q(n70180) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][28]  ( .D(n104188), 
        .CK(Clk), .RN(n106397), .Q(n107777) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][28]  ( .D(n104161), 
        .CK(Clk), .RN(n106486), .Q(n107778) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24679 ), .CK(Clk), .RN(n106490), .Q(
        n107779), .QN(n103303) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24647 ), .CK(Clk), .RN(n106488), .Q(n70185) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24615 ), .CK(Clk), .RN(n106441), .Q(
        n107780) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24551 ), .CK(Clk), .RN(n106484), .Q(
        n107781) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24519 ), .CK(Clk), .RN(Rst), .Q(n107782), 
        .QN(n102694) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24487 ), .CK(Clk), .RN(Rst), .Q(n70190), 
        .QN(n104633) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24455 ), .CK(Clk), .RN(Rst), .Q(n107783)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24423 ), .CK(Clk), .RN(n106395), .Q(
        n107784) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24391 ), .CK(Clk), .RN(Rst), .Q(n107785)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24359 ), .CK(Clk), .RN(Rst), .Q(n107786)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24327 ), .CK(Clk), .RN(Rst), .Q(n107787)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24295 ), .CK(Clk), .RN(n106449), .Q(
        n107788), .QN(n103301) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24263 ), .CK(Clk), .RN(n106422), .Q(
        n107789) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24231 ), .CK(Clk), .RN(n106421), .Q(
        n107790) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24167 ), .CK(Clk), .RN(n106420), .Q(
        n107791) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24135 ), .CK(Clk), .RN(n106473), .Q(
        n107792) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24071 ), .CK(Clk), .RN(n106426), .Q(
        n107793), .QN(n103860) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24039 ), .CK(Clk), .RN(Rst), .Q(n70204) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24007 ), .CK(Clk), .RN(Rst), .Q(n107794), 
        .QN(n101054) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23975 ), .CK(Clk), .RN(n106372), .Q(n70206) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23943 ), .CK(Clk), .RN(n106458), .Q(
        n107795) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23911 ), .CK(Clk), .RN(n106457), .Q(n70208), .QN(n104652) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23879 ), .CK(Clk), .RN(n106475), .Q(n70209) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][28]  ( .D(n104025), 
        .CK(Clk), .RN(Rst), .Q(n107796) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23783 ), .CK(Clk), .RN(n106373), .Q(
        n107797), .QN(n101024) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][28]  ( .D(n104040), 
        .CK(Clk), .RN(Rst), .Q(n107798) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23719 ), .CK(Clk), .RN(Rst), .Q(n70214) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23687 ), .CK(Clk), .RN(Rst), .Q(n107799)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23655 ), .CK(Clk), .RN(Rst), .Q(n70216) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23623 ), .CK(Clk), .RN(Rst), .Q(n107800)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23591 ), .CK(Clk), .RN(Rst), .Q(n107801)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][28]  ( .D(n104034), 
        .CK(Clk), .RN(Rst), .Q(n107802), .QN(n103855) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23527 ), .CK(Clk), .RN(Rst), .Q(n107803)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][28]  ( .D(n104053), 
        .CK(Clk), .RN(Rst), .Q(n70221) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23463 ), .CK(Clk), .RN(Rst), .Q(n70222) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23431 ), .CK(Clk), .RN(Rst), .Q(n107804)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23399 ), .CK(Clk), .RN(Rst), .Q(n107805)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23367 ), .CK(Clk), .RN(n106381), .Q(n70225) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23335 ), .CK(Clk), .RN(n106406), .Q(
        n107806) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23303 ), .CK(Clk), .RN(Rst), .Q(n107807)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23239 ), .CK(Clk), .RN(n106378), .Q(
        n107809) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23207 ), .CK(Clk), .RN(n106382), .Q(
        n107810) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][28]  ( .D(n104002), 
        .CK(Clk), .RN(n106371), .Q(n107811) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23143 ), .CK(Clk), .RN(n106445), .Q(
        n107812) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23111 ), .CK(Clk), .RN(n106417), .Q(
        n107813) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23079 ), .CK(Clk), .RN(Rst), .Q(n107814)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23047 ), .CK(Clk), .RN(Rst), .Q(n107815)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23015 ), .CK(Clk), .RN(Rst), .Q(n107816)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22983 ), .CK(Clk), .RN(Rst), .Q(n107817)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22951 ), .CK(Clk), .RN(n106481), .Q(n70238) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22919 ), .CK(Clk), .RN(n106431), .Q(n70239) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22887 ), .CK(Clk), .RN(Rst), .Q(n107818)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22855 ), .CK(Clk), .RN(n106503), .Q(
        n107819) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22823 ), .CK(Clk), .RN(n106419), .Q(n70242) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22791 ), .CK(Clk), .RN(n106480), .Q(
        n107820) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22759 ), .CK(Clk), .RN(n106501), .Q(n70244) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22727 ), .CK(Clk), .RN(n106491), .Q(
        n107821) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22695 ), .CK(Clk), .RN(Rst), .Q(n107822)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22663 ), .CK(Clk), .RN(Rst), .Q(n107823)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22631 ), .CK(Clk), .RN(n106412), .Q(
        n107824) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22599 ), .CK(Clk), .RN(n106413), .Q(n70249) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25895 ), .CK(Clk), .RN(n106383), .Q(n70251) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][28]  ( .D(n104264), 
        .CK(Clk), .RN(n106403), .Q(n107826) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25959 ), .CK(Clk), .RN(n106384), .Q(
        n107827) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25991 ), .CK(Clk), .RN(n106404), .Q(
        n107828) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26023 ), .CK(Clk), .RN(n106408), .Q(
        n107829) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26055 ), .CK(Clk), .RN(n106387), .Q(
        n107830) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26087 ), .CK(Clk), .RN(n106388), .Q(
        n107831) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26151 ), .CK(Clk), .RN(n106389), .Q(
        n107833), .QN(n102133) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][28]  ( .D(n104242), 
        .CK(Clk), .RN(n106380), .Q(n70260) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26215 ), .CK(Clk), .RN(Rst), .Q(n70261) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26247 ), .CK(Clk), .RN(Rst), .Q(n107834)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26279 ), .CK(Clk), .RN(Rst), .Q(n70263) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26311 ), .CK(Clk), .RN(n106371), .Q(
        n107835) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26343 ), .CK(Clk), .RN(Rst), .Q(n107836)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26375 ), .CK(Clk), .RN(Rst), .Q(n107837)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26407 ), .CK(Clk), .RN(Rst), .Q(n107838)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26439 ), .CK(Clk), .RN(Rst), .Q(n107839)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26471 ), .CK(Clk), .RN(Rst), .Q(n107840)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26503 ), .CK(Clk), .RN(n106378), .Q(
        n107841), .QN(n103869) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26535 ), .CK(Clk), .RN(n106379), .Q(
        n107842) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26599 ), .CK(Clk), .RN(n106448), .Q(
        n107844) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26631 ), .CK(Clk), .RN(n106448), .Q(
        n107845) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][28]  ( .D(n106987), 
        .CK(Clk), .RN(n106448), .Q(n107846) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26695 ), .CK(Clk), .RN(n106448), .Q(
        n107847), .QN(n102702) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26727 ), .CK(Clk), .RN(n106448), .Q(
        n107848), .QN(n103310) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26759 ), .CK(Clk), .RN(n106448), .Q(n70278), .QN(n104553) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][28]  ( .D(n107018), 
        .CK(Clk), .RN(n106448), .Q(n107849), .QN(n102134) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26855 ), .CK(Clk), .RN(n106448), .Q(
        n107851), .QN(n103311) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[28]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107090), .Q(
        \DLX_Datapath/next_A_IDEX[28] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[28]  ( .D(n106613), .CK(Clk), .RN(n106448), 
        .Q(n107852) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[28]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107056), .Q(
        \DLX_Datapath/next_B_IDEX [28]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[28]  ( .D(n106686), .CK(Clk), .RN(n106448), 
        .Q(n70283), .QN(n104668) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[28]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [28]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [28]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[28]  ( .D(n103915), .GN(n60158), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [28]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[28]  ( .D(n104330), .CK(Clk), .RN(
        n106447), .Q(DataAddr[28]), .QN(n58691) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[28]  ( .D(n58998), .CK(Clk), .RN(n106447), 
        .Q(n107853) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[28]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [28]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [28]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[28]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [28]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [28]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[28]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N141 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [28]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[31]  ( .D(n106925), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [31]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[31]  ( .D(n104331), .CK(Clk), .RN(
        n106447), .Q(DataAddr[31]), .QN(n58688) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25866 ), .CK(Clk), .RN(n106447), .Q(n70291) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25834 ), .CK(Clk), .RN(n106447), .Q(
        n107855) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25802 ), .CK(Clk), .RN(n106447), .Q(
        n107856) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25770 ), .CK(Clk), .RN(n106447), .Q(
        n107857) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25706 ), .CK(Clk), .RN(n106447), .Q(
        n107858) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25642 ), .CK(Clk), .RN(n106447), .Q(
        n107859) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25610 ), .CK(Clk), .RN(n106446), .Q(
        n107860) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25578 ), .CK(Clk), .RN(n106446), .Q(
        n107861) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25546 ), .CK(Clk), .RN(n106446), .Q(
        n107862) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25514 ), .CK(Clk), .RN(n106446), .Q(
        n107863), .QN(n100561) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25482 ), .CK(Clk), .RN(n106446), .Q(n70303) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25450 ), .CK(Clk), .RN(n106446), .Q(n70304) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25418 ), .CK(Clk), .RN(n106446), .Q(
        n107864) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25386 ), .CK(Clk), .RN(n106446), .Q(
        n107865) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][31]  ( .D(n104306), 
        .CK(Clk), .RN(n106446), .Q(n107866) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25290 ), .CK(Clk), .RN(n106446), .Q(
        n107868), .QN(n102745) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25258 ), .CK(Clk), .RN(n106446), .Q(
        n107869), .QN(n102174) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25226 ), .CK(Clk), .RN(n106445), .Q(
        n107870) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25194 ), .CK(Clk), .RN(n106445), .Q(n70312) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25162 ), .CK(Clk), .RN(n106445), .Q(
        n107871) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][31]  ( .D(n104288), 
        .CK(Clk), .RN(n106445), .Q(n107872) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25066 ), .CK(Clk), .RN(n106445), .Q(n70316), .QN(n104583) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][31]  ( .D(n104213), 
        .CK(Clk), .RN(n106445), .Q(n70317) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25002 ), .CK(Clk), .RN(n106445), .Q(
        n107873), .QN(n100593) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][31]  ( .D(n104294), 
        .CK(Clk), .RN(n106445), .Q(n107874) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24938 ), .CK(Clk), .RN(n106445), .Q(n70320) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24906 ), .CK(Clk), .RN(n106445), .Q(n70321), .QN(n104655) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24874 ), .CK(Clk), .RN(n106445), .Q(
        n107875) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24842 ), .CK(Clk), .RN(n106456), .Q(
        n107876) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24810 ), .CK(Clk), .RN(n106372), .Q(n70324) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24778 ), .CK(Clk), .RN(n106480), .Q(
        n107877) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][31]  ( .D(n104170), 
        .CK(Clk), .RN(n106457), .Q(n107878) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24682 ), .CK(Clk), .RN(n106491), .Q(
        n107879), .QN(n101148) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24650 ), .CK(Clk), .RN(n106481), .Q(n70329) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24618 ), .CK(Clk), .RN(n106456), .Q(n70330) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24554 ), .CK(Clk), .RN(n106455), .Q(
        n107880) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24522 ), .CK(Clk), .RN(n106458), .Q(
        n107881), .QN(n102741) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24490 ), .CK(Clk), .RN(n106419), .Q(n70334), .QN(n104636) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][31]  ( .D(n104146), 
        .CK(Clk), .RN(Rst), .Q(n107882) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24426 ), .CK(Clk), .RN(Rst), .Q(n107883)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][31]  ( .D(n104190), 
        .CK(Clk), .RN(n106431), .Q(n107884) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24362 ), .CK(Clk), .RN(n106444), .Q(
        n107885) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24330 ), .CK(Clk), .RN(Rst), .Q(n107886)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24298 ), .CK(Clk), .RN(n106477), .Q(
        n107887), .QN(n103344) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24266 ), .CK(Clk), .RN(Rst), .Q(n107888)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24170 ), .CK(Clk), .RN(Rst), .Q(n107889)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24138 ), .CK(Clk), .RN(Rst), .Q(n107890)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][31]  ( .D(n104079), 
        .CK(Clk), .RN(Rst), .Q(n107891) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24042 ), .CK(Clk), .RN(n106492), .Q(n70348) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24010 ), .CK(Clk), .RN(Rst), .Q(n107892), 
        .QN(n102739) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23978 ), .CK(Clk), .RN(Rst), .Q(n70350) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][31]  ( .D(n104090), 
        .CK(Clk), .RN(Rst), .Q(n107893), .QN(n100775) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23914 ), .CK(Clk), .RN(Rst), .Q(n107894), 
        .QN(n103342) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][31]  ( .D(n104126), 
        .CK(Clk), .RN(Rst), .Q(n107895) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23818 ), .CK(Clk), .RN(Rst), .Q(n70355) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23786 ), .CK(Clk), .RN(Rst), .Q(n107896), 
        .QN(n101021) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23754 ), .CK(Clk), .RN(n106377), .Q(
        n107897) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23722 ), .CK(Clk), .RN(Rst), .Q(n70358) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23690 ), .CK(Clk), .RN(n106427), .Q(
        n107898), .QN(n100992) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23658 ), .CK(Clk), .RN(Rst), .Q(n70360) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23626 ), .CK(Clk), .RN(n106394), .Q(
        n107899) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23594 ), .CK(Clk), .RN(n106478), .Q(
        n107900) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][31]  ( .D(n104028), 
        .CK(Clk), .RN(Rst), .Q(n70363) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23530 ), .CK(Clk), .RN(n106477), .Q(n70364) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23498 ), .CK(Clk), .RN(Rst), .Q(n70365) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23466 ), .CK(Clk), .RN(n106376), .Q(n70366) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23434 ), .CK(Clk), .RN(n106452), .Q(n70367) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23402 ), .CK(Clk), .RN(n106400), .Q(
        n107901) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23370 ), .CK(Clk), .RN(n106451), .Q(n70369) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23338 ), .CK(Clk), .RN(n106450), .Q(
        n107902) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23306 ), .CK(Clk), .RN(n106504), .Q(
        n107903) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23242 ), .CK(Clk), .RN(Rst), .Q(n107905)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23210 ), .CK(Clk), .RN(Rst), .Q(n107906)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23178 ), .CK(Clk), .RN(Rst), .Q(n107907)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23114 ), .CK(Clk), .RN(n106432), .Q(
        n107908) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23082 ), .CK(Clk), .RN(Rst), .Q(n107909)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23050 ), .CK(Clk), .RN(n106433), .Q(
        n107910) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23018 ), .CK(Clk), .RN(n106459), .Q(
        n107911) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22986 ), .CK(Clk), .RN(n106434), .Q(
        n107912) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22954 ), .CK(Clk), .RN(Rst), .Q(n70382) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22922 ), .CK(Clk), .RN(n106416), .Q(n70383) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22890 ), .CK(Clk), .RN(n106384), .Q(
        n107913) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22858 ), .CK(Clk), .RN(Rst), .Q(n107914)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22826 ), .CK(Clk), .RN(n106441), .Q(n70386) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22794 ), .CK(Clk), .RN(n106445), .Q(
        n107915) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22762 ), .CK(Clk), .RN(Rst), .Q(n70388) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22730 ), .CK(Clk), .RN(n106379), .Q(
        n107916) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22698 ), .CK(Clk), .RN(n106380), .Q(
        n107917) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22666 ), .CK(Clk), .RN(n106406), .Q(
        n107918) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22634 ), .CK(Clk), .RN(n106378), .Q(
        n107919) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22602 ), .CK(Clk), .RN(n106385), .Q(
        n107920) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][31]  ( .D(n104261), 
        .CK(Clk), .RN(Rst), .Q(n107922) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25962 ), .CK(Clk), .RN(n106387), .Q(
        n107923) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25994 ), .CK(Clk), .RN(n106388), .Q(
        n107924), .QN(n103911) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26026 ), .CK(Clk), .RN(n106389), .Q(
        n107925) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26058 ), .CK(Clk), .RN(n106403), .Q(
        n107926) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26090 ), .CK(Clk), .RN(n106412), .Q(
        n107927) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26154 ), .CK(Clk), .RN(n106407), .Q(
        n107928), .QN(n102178) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][31]  ( .D(n104243), 
        .CK(Clk), .RN(Rst), .Q(n70404) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26218 ), .CK(Clk), .RN(n106414), .Q(n70405) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26250 ), .CK(Clk), .RN(n106461), .Q(
        n107929) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26282 ), .CK(Clk), .RN(n106487), .Q(n70407) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26314 ), .CK(Clk), .RN(n106399), .Q(
        n107930) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26346 ), .CK(Clk), .RN(Rst), .Q(n107931)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26378 ), .CK(Clk), .RN(Rst), .Q(n107932)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26410 ), .CK(Clk), .RN(Rst), .Q(n107933)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26442 ), .CK(Clk), .RN(n106447), .Q(
        n107934) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26474 ), .CK(Clk), .RN(n106375), .Q(
        n107935) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26506 ), .CK(Clk), .RN(n106374), .Q(
        n107936), .QN(n103912) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26538 ), .CK(Clk), .RN(n106384), .Q(
        n107937) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26602 ), .CK(Clk), .RN(n106404), .Q(
        n107939) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26634 ), .CK(Clk), .RN(n106399), .Q(
        n107940) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][31]  ( .D(n106989), 
        .CK(Clk), .RN(n106459), .Q(n107941) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26698 ), .CK(Clk), .RN(n106484), .Q(
        n107942), .QN(n102747) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26730 ), .CK(Clk), .RN(n106443), .Q(
        n107943), .QN(n103350) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26762 ), .CK(Clk), .RN(n106486), .Q(n70422), .QN(n104556) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][31]  ( .D(n107020), 
        .CK(Clk), .RN(n106429), .Q(n107944), .QN(n102179) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26858 ), .CK(Clk), .RN(Rst), .Q(n107946), 
        .QN(n103351) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[31]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107092), .Q(
        \DLX_Datapath/next_A_IDEX[31] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[31]  ( .D(n106614), .CK(Clk), .RN(Rst), .Q(
        n107947) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[31]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107058), .Q(
        \DLX_Datapath/next_B_IDEX [31]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[31]  ( .D(n106688), .CK(Clk), .RN(n106394), 
        .Q(n70427), .QN(n104671) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[31]  ( .D(n58995), .CK(Clk), .RN(n106476), 
        .Q(n107948) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[31]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [31]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [31]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[31]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [31]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [31]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[31]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [31]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [31]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[31]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N176 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [31]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[30]  ( .D(n106923), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [30]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[30]  ( .D(n104332), .CK(Clk), .RN(
        n106444), .Q(DataAddr[30]), .QN(n58685) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25865 ), .CK(Clk), .RN(n106412), .Q(n70433) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25833 ), .CK(Clk), .RN(Rst), .Q(n107952)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][30]  ( .D(n104216), 
        .CK(Clk), .RN(n106446), .Q(n107953) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25769 ), .CK(Clk), .RN(n106407), .Q(
        n107954) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25705 ), .CK(Clk), .RN(n106414), .Q(
        n107955) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25641 ), .CK(Clk), .RN(n106387), .Q(
        n107956) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25609 ), .CK(Clk), .RN(n106389), .Q(
        n107957) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25577 ), .CK(Clk), .RN(n106403), .Q(
        n107958) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25545 ), .CK(Clk), .RN(n106388), .Q(
        n107959) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25513 ), .CK(Clk), .RN(n106419), .Q(
        n107960), .QN(n100562) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25481 ), .CK(Clk), .RN(n106456), .Q(n70445) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25449 ), .CK(Clk), .RN(n106480), .Q(n70446) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25417 ), .CK(Clk), .RN(n106491), .Q(
        n107961) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25385 ), .CK(Clk), .RN(n106481), .Q(
        n107962) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25353 ), .CK(Clk), .RN(Rst), .Q(n107963)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25289 ), .CK(Clk), .RN(n106501), .Q(
        n107965), .QN(n102733) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25257 ), .CK(Clk), .RN(n106455), .Q(
        n107966), .QN(n102160) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25225 ), .CK(Clk), .RN(Rst), .Q(n107967)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25193 ), .CK(Clk), .RN(n106503), .Q(n70454) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25161 ), .CK(Clk), .RN(Rst), .Q(n107968)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25097 ), .CK(Clk), .RN(Rst), .Q(n107969)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25065 ), .CK(Clk), .RN(n106374), .Q(n70458), .QN(n104614) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25033 ), .CK(Clk), .RN(Rst), .Q(n107970)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25001 ), .CK(Clk), .RN(Rst), .Q(n107971), 
        .QN(n100594) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24969 ), .CK(Clk), .RN(Rst), .Q(n70461) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24937 ), .CK(Clk), .RN(n106375), .Q(n70462) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24905 ), .CK(Clk), .RN(n106487), .Q(n70463), .QN(n104654) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24873 ), .CK(Clk), .RN(n106447), .Q(
        n107972) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24841 ), .CK(Clk), .RN(n106461), .Q(
        n107973) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24809 ), .CK(Clk), .RN(n106416), .Q(n70466) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24777 ), .CK(Clk), .RN(n106399), .Q(
        n107974) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24713 ), .CK(Clk), .RN(Rst), .Q(n107975)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24681 ), .CK(Clk), .RN(n106464), .Q(n70470), .QN(n104648) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24649 ), .CK(Clk), .RN(Rst), .Q(n70471) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24617 ), .CK(Clk), .RN(n106396), .Q(n70472) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24521 ), .CK(Clk), .RN(n106435), .Q(
        n107976), .QN(n102727) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24489 ), .CK(Clk), .RN(n106462), .Q(n70476), .QN(n104635) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24457 ), .CK(Clk), .RN(n106440), .Q(
        n107977) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24425 ), .CK(Clk), .RN(n106463), .Q(
        n107978) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24393 ), .CK(Clk), .RN(n106442), .Q(
        n107979) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24361 ), .CK(Clk), .RN(n106446), .Q(
        n107980) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24329 ), .CK(Clk), .RN(Rst), .Q(n107981)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24297 ), .CK(Clk), .RN(n106396), .Q(
        n107982), .QN(n103332) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24265 ), .CK(Clk), .RN(n106435), .Q(
        n107983) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24169 ), .CK(Clk), .RN(n106442), .Q(
        n107984) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24137 ), .CK(Clk), .RN(Rst), .Q(n107985)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24073 ), .CK(Clk), .RN(n106440), .Q(
        n107986) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24041 ), .CK(Clk), .RN(n106462), .Q(n70490) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24009 ), .CK(Clk), .RN(n106464), .Q(
        n107987), .QN(n102725) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23977 ), .CK(Clk), .RN(n106463), .Q(n70492) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23945 ), .CK(Clk), .RN(n106467), .Q(
        n107988), .QN(n103893) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23913 ), .CK(Clk), .RN(Rst), .Q(n70494), 
        .QN(n104653) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23881 ), .CK(Clk), .RN(Rst), .Q(n107989)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23817 ), .CK(Clk), .RN(Rst), .Q(n70497) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23785 ), .CK(Clk), .RN(Rst), .Q(n107990), 
        .QN(n101022) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23753 ), .CK(Clk), .RN(Rst), .Q(n107991)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23721 ), .CK(Clk), .RN(Rst), .Q(n70500) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23689 ), .CK(Clk), .RN(Rst), .Q(n107992), 
        .QN(n100993) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23657 ), .CK(Clk), .RN(n106469), .Q(n70502) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23625 ), .CK(Clk), .RN(Rst), .Q(n107993)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23593 ), .CK(Clk), .RN(Rst), .Q(n107994)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23561 ), .CK(Clk), .RN(n106443), .Q(
        n107995), .QN(n103890) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23529 ), .CK(Clk), .RN(n106443), .Q(n70506) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23497 ), .CK(Clk), .RN(n106443), .Q(n70507) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23465 ), .CK(Clk), .RN(n106443), .Q(n70508) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23433 ), .CK(Clk), .RN(n106443), .Q(
        n107996) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23401 ), .CK(Clk), .RN(n106443), .Q(
        n107997) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23369 ), .CK(Clk), .RN(n106443), .Q(n70511) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23337 ), .CK(Clk), .RN(n106443), .Q(
        n107998) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23305 ), .CK(Clk), .RN(n106443), .Q(
        n107999) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23241 ), .CK(Clk), .RN(n106443), .Q(
        n108001) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23209 ), .CK(Clk), .RN(n106443), .Q(
        n108002) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23177 ), .CK(Clk), .RN(n106442), .Q(
        n108003) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23113 ), .CK(Clk), .RN(n106442), .Q(
        n108004) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23081 ), .CK(Clk), .RN(n106442), .Q(
        n108005) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23049 ), .CK(Clk), .RN(n106442), .Q(
        n108006) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23017 ), .CK(Clk), .RN(n106442), .Q(
        n108007) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22985 ), .CK(Clk), .RN(n106442), .Q(
        n108008) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22953 ), .CK(Clk), .RN(n106442), .Q(n70524) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22921 ), .CK(Clk), .RN(n106442), .Q(n70525) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22889 ), .CK(Clk), .RN(n106442), .Q(
        n108009) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22857 ), .CK(Clk), .RN(n106442), .Q(
        n108010) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22825 ), .CK(Clk), .RN(n106442), .Q(
        n108011) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22793 ), .CK(Clk), .RN(n106441), .Q(
        n108012) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22761 ), .CK(Clk), .RN(n106441), .Q(n70530) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22729 ), .CK(Clk), .RN(n106441), .Q(
        n108013) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22697 ), .CK(Clk), .RN(n106441), .Q(
        n108014) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22665 ), .CK(Clk), .RN(n106441), .Q(
        n108015) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22633 ), .CK(Clk), .RN(n106441), .Q(
        n108016) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22601 ), .CK(Clk), .RN(n106441), .Q(n70535) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25897 ), .CK(Clk), .RN(n106441), .Q(n70537) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][30]  ( .D(n104263), 
        .CK(Clk), .RN(n106441), .Q(n108018) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25961 ), .CK(Clk), .RN(n106441), .Q(
        n108019) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25993 ), .CK(Clk), .RN(n106441), .Q(
        n108020), .QN(n103900) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26025 ), .CK(Clk), .RN(n106440), .Q(
        n108021) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26057 ), .CK(Clk), .RN(n106440), .Q(
        n108022) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26089 ), .CK(Clk), .RN(n106440), .Q(
        n108023) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26153 ), .CK(Clk), .RN(n106440), .Q(
        n108024), .QN(n102164) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][30]  ( .D(n104251), 
        .CK(Clk), .RN(n106440), .Q(n70546) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26217 ), .CK(Clk), .RN(n106440), .Q(n70547) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26249 ), .CK(Clk), .RN(n106440), .Q(
        n108025) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26281 ), .CK(Clk), .RN(n106440), .Q(n70549) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26313 ), .CK(Clk), .RN(n106440), .Q(
        n108026) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26345 ), .CK(Clk), .RN(n106440), .Q(
        n108027) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26377 ), .CK(Clk), .RN(n106440), .Q(
        n108028) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26409 ), .CK(Clk), .RN(Rst), .Q(n108029)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26441 ), .CK(Clk), .RN(Rst), .Q(n108030)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26473 ), .CK(Clk), .RN(Rst), .Q(n108031)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26505 ), .CK(Clk), .RN(Rst), .Q(n108032), 
        .QN(n103901) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26537 ), .CK(Clk), .RN(Rst), .Q(n108033)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26601 ), .CK(Clk), .RN(Rst), .Q(n108035)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26633 ), .CK(Clk), .RN(Rst), .Q(n108036)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][30]  ( .D(n106988), 
        .CK(Clk), .RN(Rst), .Q(n108037) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26697 ), .CK(Clk), .RN(Rst), .Q(n108038), 
        .QN(n102734) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26729 ), .CK(Clk), .RN(Rst), .Q(n108039), 
        .QN(n103337) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26761 ), .CK(Clk), .RN(Rst), .Q(n70564), 
        .QN(n104555) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][30]  ( .D(n107019), 
        .CK(Clk), .RN(Rst), .Q(n108040), .QN(n102165) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26857 ), .CK(Clk), .RN(Rst), .Q(n108042), 
        .QN(n103338) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[30]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107091), .Q(
        \DLX_Datapath/next_A_IDEX[30] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[30]  ( .D(n106630), .CK(Clk), .RN(Rst), .Q(
        n108043) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[30]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107057), .Q(
        \DLX_Datapath/next_B_IDEX [30]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[30]  ( .D(n106674), .CK(Clk), .RN(Rst), .Q(
        n70569), .QN(n104670) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[30]  ( .D(n58992), .CK(Clk), .RN(Rst), .Q(
        n108044) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[30]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [30]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [30]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[30]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [30]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [30]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[27]  ( .D(n106921), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [27]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[27]  ( .D(n104333), .CK(Clk), .RN(Rst), .Q(DataAddr[27]), .QN(n58682) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[27]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [27]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [27]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[27]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N172 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [27]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[26]  ( .D(n106919), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [26]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[26]  ( .D(n104334), .CK(Clk), .RN(Rst), .Q(DataAddr[26]), .QN(n58680) );
  DFFR_X2 \DLX_Datapath/PC_reg[26]  ( .D(n60299), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [2]), .QN(n57427) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[24]  ( .D(n106525), .CK(Clk), .RN(Rst), 
        .Q(net2410613) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[24]  ( .D(n106659), .CK(Clk), .RN(Rst), 
        .Q(n70575) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[24]  ( .D(n58987), .CK(Clk), .RN(n106439), .Q(n108048), .QN(n59347) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[25]  ( .D(n106524), .CK(Clk), .RN(n106439), .Q(n108049) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[25]  ( .D(n106660), .CK(Clk), .RN(n106439), .Q(n70576) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[25]  ( .D(n58986), .CK(Clk), .RN(n106439), .Q(n108050), .QN(n59348) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[26]  ( .D(n106523), .CK(Clk), .RN(n106439), .Q(n108051) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[26]  ( .D(n106640), .CK(Clk), .RN(n106439), .Q(n70577) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[26]  ( .D(n58985), .CK(Clk), .RN(n106439), .Q(n108052), .QN(n59349) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25861 ), .CK(Clk), .RN(n106439), .Q(n70580) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25829 ), .CK(Clk), .RN(n106439), .Q(
        n108054) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25797 ), .CK(Clk), .RN(n106439), .Q(
        n108055) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25765 ), .CK(Clk), .RN(n106438), .Q(
        n108056) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25701 ), .CK(Clk), .RN(n106438), .Q(
        n108057) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25637 ), .CK(Clk), .RN(n106438), .Q(
        n108058) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25605 ), .CK(Clk), .RN(n106438), .Q(
        n108059), .QN(n103835) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25573 ), .CK(Clk), .RN(n106438), .Q(
        n108060) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25541 ), .CK(Clk), .RN(n106438), .Q(
        n108061) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25509 ), .CK(Clk), .RN(n106438), .Q(
        n108062), .QN(n100566) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25477 ), .CK(Clk), .RN(n106438), .Q(n70592) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25445 ), .CK(Clk), .RN(n106438), .Q(
        n108063) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25413 ), .CK(Clk), .RN(n106438), .Q(
        n108064) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25381 ), .CK(Clk), .RN(n106437), .Q(
        n108065) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25349 ), .CK(Clk), .RN(n106437), .Q(
        n108066) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25317 ), .CK(Clk), .RN(n106437), .Q(
        n108067), .QN(n103271) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25285 ), .CK(Clk), .RN(n106437), .Q(
        n108068), .QN(n102672) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25253 ), .CK(Clk), .RN(n106437), .Q(
        n108069), .QN(n102101) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25221 ), .CK(Clk), .RN(n106437), .Q(
        n108070) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25189 ), .CK(Clk), .RN(n106437), .Q(n70601) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25157 ), .CK(Clk), .RN(n106437), .Q(
        n108071) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25093 ), .CK(Clk), .RN(n106437), .Q(
        n108072) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25061 ), .CK(Clk), .RN(n106437), .Q(n70605), .QN(n104610) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25029 ), .CK(Clk), .RN(n106437), .Q(
        n108073) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24997 ), .CK(Clk), .RN(n106488), .Q(
        n108074), .QN(n100598) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24965 ), .CK(Clk), .RN(n106473), .Q(
        n108075) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24933 ), .CK(Clk), .RN(n106377), .Q(n70609) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24901 ), .CK(Clk), .RN(n106478), .Q(
        n108076), .QN(n101154) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24869 ), .CK(Clk), .RN(n106402), .Q(
        n108077) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24837 ), .CK(Clk), .RN(n106453), .Q(
        n108078) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24805 ), .CK(Clk), .RN(n106413), .Q(n70613) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24773 ), .CK(Clk), .RN(Rst), .Q(n108079)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24709 ), .CK(Clk), .RN(n106454), .Q(
        n108080) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24677 ), .CK(Clk), .RN(n106379), .Q(
        n108081), .QN(n103267) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24645 ), .CK(Clk), .RN(n106499), .Q(n70618) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24613 ), .CK(Clk), .RN(n106501), .Q(n70619) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24549 ), .CK(Clk), .RN(n106500), .Q(
        n108082) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24517 ), .CK(Clk), .RN(n106499), .Q(
        n108083), .QN(n102665) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24485 ), .CK(Clk), .RN(n106419), .Q(n70623), .QN(n104631) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24453 ), .CK(Clk), .RN(n106436), .Q(
        n108084) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24421 ), .CK(Clk), .RN(Rst), .Q(n108085)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24389 ), .CK(Clk), .RN(Rst), .Q(n108086)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24357 ), .CK(Clk), .RN(n106498), .Q(
        n108087) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24325 ), .CK(Clk), .RN(n106497), .Q(
        n108088) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24293 ), .CK(Clk), .RN(n106503), .Q(
        n108089), .QN(n103265) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24261 ), .CK(Clk), .RN(n106502), .Q(
        n108090) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24165 ), .CK(Clk), .RN(n106444), .Q(
        n108091) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24133 ), .CK(Clk), .RN(n106444), .Q(
        n108092) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24069 ), .CK(Clk), .RN(n106444), .Q(
        n108093), .QN(n103829) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24037 ), .CK(Clk), .RN(n106444), .Q(n70637) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24005 ), .CK(Clk), .RN(n106444), .Q(
        n108094), .QN(n102663) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23973 ), .CK(Clk), .RN(n106444), .Q(n70639) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23941 ), .CK(Clk), .RN(n106444), .Q(
        n108095) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23909 ), .CK(Clk), .RN(n106444), .Q(
        n108096), .QN(n103263) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23877 ), .CK(Clk), .RN(n106444), .Q(
        n108097) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23813 ), .CK(Clk), .RN(Rst), .Q(n108098)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23781 ), .CK(Clk), .RN(Rst), .Q(n108099), 
        .QN(n101026) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23749 ), .CK(Clk), .RN(n106492), .Q(
        n108100) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23717 ), .CK(Clk), .RN(Rst), .Q(n70647) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23685 ), .CK(Clk), .RN(Rst), .Q(n108101)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23653 ), .CK(Clk), .RN(Rst), .Q(n70649) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23621 ), .CK(Clk), .RN(Rst), .Q(n108102)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23589 ), .CK(Clk), .RN(Rst), .Q(n108103)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23557 ), .CK(Clk), .RN(Rst), .Q(n70652) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23525 ), .CK(Clk), .RN(n106372), .Q(
        n108104) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][26]  ( .D(n104054), 
        .CK(Clk), .RN(Rst), .Q(n70654) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23461 ), .CK(Clk), .RN(Rst), .Q(n70655) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23429 ), .CK(Clk), .RN(n106375), .Q(n70656) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23397 ), .CK(Clk), .RN(n106371), .Q(
        n108105) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23365 ), .CK(Clk), .RN(n106382), .Q(n70658) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23333 ), .CK(Clk), .RN(n106498), .Q(
        n108106) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23301 ), .CK(Clk), .RN(Rst), .Q(n108107)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23269 ), .CK(Clk), .RN(n106381), .Q(
        n108108), .QN(n103261) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23237 ), .CK(Clk), .RN(n106469), .Q(
        n108109) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23205 ), .CK(Clk), .RN(Rst), .Q(n108110)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23141 ), .CK(Clk), .RN(n106381), .Q(
        n108111) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23109 ), .CK(Clk), .RN(Rst), .Q(n108112)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23077 ), .CK(Clk), .RN(Rst), .Q(n108113)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23045 ), .CK(Clk), .RN(Rst), .Q(n108114)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23013 ), .CK(Clk), .RN(Rst), .Q(n108115)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22981 ), .CK(Clk), .RN(Rst), .Q(n108116)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22949 ), .CK(Clk), .RN(Rst), .Q(n70671) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22917 ), .CK(Clk), .RN(n106492), .Q(n70672) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22885 ), .CK(Clk), .RN(Rst), .Q(n108117)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22853 ), .CK(Clk), .RN(Rst), .Q(n108118)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22821 ), .CK(Clk), .RN(Rst), .Q(n70675) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22789 ), .CK(Clk), .RN(Rst), .Q(n108119)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22757 ), .CK(Clk), .RN(Rst), .Q(n70677) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22725 ), .CK(Clk), .RN(Rst), .Q(n108120)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22693 ), .CK(Clk), .RN(Rst), .Q(n108121)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22661 ), .CK(Clk), .RN(Rst), .Q(n108122)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22629 ), .CK(Clk), .RN(Rst), .Q(n108123)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22597 ), .CK(Clk), .RN(Rst), .Q(n108124)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][26]  ( .D(n104262), 
        .CK(Clk), .RN(Rst), .Q(n108126) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25957 ), .CK(Clk), .RN(Rst), .Q(n108127)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25989 ), .CK(Clk), .RN(Rst), .Q(n108128)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26021 ), .CK(Clk), .RN(Rst), .Q(n108129)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26053 ), .CK(Clk), .RN(Rst), .Q(n108130)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26085 ), .CK(Clk), .RN(Rst), .Q(n108131)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26149 ), .CK(Clk), .RN(n106454), .Q(
        n108133), .QN(n102105) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][26]  ( .D(n104245), 
        .CK(Clk), .RN(n106395), .Q(n70693) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26213 ), .CK(Clk), .RN(Rst), .Q(n70694) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26245 ), .CK(Clk), .RN(n106377), .Q(
        n108134) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26277 ), .CK(Clk), .RN(Rst), .Q(n70696) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26309 ), .CK(Clk), .RN(Rst), .Q(n108135)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26341 ), .CK(Clk), .RN(n106448), .Q(
        n108136) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26373 ), .CK(Clk), .RN(n106445), .Q(
        n108137) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26405 ), .CK(Clk), .RN(n106498), .Q(
        n108138) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26437 ), .CK(Clk), .RN(Rst), .Q(n108139)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26469 ), .CK(Clk), .RN(Rst), .Q(n108140)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26501 ), .CK(Clk), .RN(Rst), .Q(n108141), 
        .QN(n103837) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26533 ), .CK(Clk), .RN(Rst), .Q(n108142)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26597 ), .CK(Clk), .RN(Rst), .Q(n108144)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26629 ), .CK(Clk), .RN(Rst), .Q(n108145)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][26]  ( .D(n106985), 
        .CK(Clk), .RN(Rst), .Q(n108146) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26693 ), .CK(Clk), .RN(Rst), .Q(n108147), 
        .QN(n102673) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26725 ), .CK(Clk), .RN(Rst), .Q(n108148), 
        .QN(n103274) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26757 ), .CK(Clk), .RN(Rst), .Q(n70711), 
        .QN(n104551) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][26]  ( .D(n107016), 
        .CK(Clk), .RN(Rst), .Q(n108149), .QN(n102106) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26853 ), .CK(Clk), .RN(Rst), .Q(n108151), 
        .QN(n103275) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[26]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107088), .Q(
        \DLX_Datapath/next_A_IDEX[26] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[26]  ( .D(n106628), .CK(Clk), .RN(Rst), .Q(
        n108152) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[26]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [26]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [26]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[26]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [26]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [26]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[26]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107054), .Q(
        \DLX_Datapath/next_B_IDEX [26]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[26]  ( .D(n106684), .CK(Clk), .RN(Rst), .Q(
        n70717), .QN(n104666) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[26]  ( .D(n58983), .CK(Clk), .RN(Rst), .Q(
        n108154) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[26]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [26]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [26]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[26]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N171 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [26]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[25]  ( .D(n106917), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [25]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[25]  ( .D(n104335), .CK(Clk), .RN(Rst), .Q(DataAddr[25]), .QN(n58673) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[25]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [25]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [25]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[25]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [25]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [25]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[24]  ( .D(n103916), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [24]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[24]  ( .D(n104336), .CK(Clk), .RN(Rst), .Q(DataAddr[24]), .QN(n58671) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[24]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [24]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [24]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[24]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [24]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [24]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[15]  ( .D(n106903), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [15]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[15]  ( .D(n104337), .CK(Clk), .RN(Rst), .Q(DataAddr[15]), .QN(n58669) );
  DFFR_X2 \DLX_Datapath/PC_reg[15]  ( .D(n60310), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [3]), .QN(n62182) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[15]  ( .D(n106534), .CK(Clk), .RN(Rst), 
        .Q(n108158) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[15]  ( .D(n106657), .CK(Clk), .RN(Rst), 
        .Q(n70726) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[15]  ( .D(n58976), .CK(Clk), .RN(Rst), 
        .Q(n108159), .QN(n59338) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25850 ), .CK(Clk), .RN(Rst), .Q(n70729) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25818 ), .CK(Clk), .RN(Rst), .Q(n108160)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][15]  ( .D(n104217), 
        .CK(Clk), .RN(Rst), .Q(n108161) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25754 ), .CK(Clk), .RN(Rst), .Q(n108162)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25690 ), .CK(Clk), .RN(Rst), .Q(n108163)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25626 ), .CK(Clk), .RN(Rst), .Q(n108164)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25594 ), .CK(Clk), .RN(Rst), .Q(n108165)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25562 ), .CK(Clk), .RN(Rst), .Q(n108166)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25530 ), .CK(Clk), .RN(Rst), .Q(n108167)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25498 ), .CK(Clk), .RN(Rst), .Q(n108168), 
        .QN(n100577) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25466 ), .CK(Clk), .RN(Rst), .Q(n70741) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25434 ), .CK(Clk), .RN(n106445), .Q(
        n108169) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25402 ), .CK(Clk), .RN(Rst), .Q(n108170)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25370 ), .CK(Clk), .RN(n106447), .Q(
        n108171) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][15]  ( .D(n104298), 
        .CK(Clk), .RN(Rst), .Q(n108172) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25306 ), .CK(Clk), .RN(n106446), .Q(
        n108173), .QN(n103060) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25274 ), .CK(Clk), .RN(Rst), .Q(n108174), 
        .QN(n102489) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25242 ), .CK(Clk), .RN(n106426), .Q(
        n108175), .QN(n101921) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25210 ), .CK(Clk), .RN(n106382), .Q(
        n108176) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25178 ), .CK(Clk), .RN(Rst), .Q(n70750) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][15]  ( .D(n104198), 
        .CK(Clk), .RN(Rst), .Q(n108177) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][15]  ( .D(n104287), 
        .CK(Clk), .RN(Rst), .Q(n108178) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25050 ), .CK(Clk), .RN(n106468), .Q(n70754), .QN(n104599) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][15]  ( .D(n104208), 
        .CK(Clk), .RN(n106496), .Q(n108179) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24986 ), .CK(Clk), .RN(n106467), .Q(
        n108180), .QN(n100609) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][15]  ( .D(n104297), 
        .CK(Clk), .RN(Rst), .Q(n108181) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24922 ), .CK(Clk), .RN(n106422), .Q(n70758) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24890 ), .CK(Clk), .RN(n106421), .Q(
        n108182), .QN(n101164) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24858 ), .CK(Clk), .RN(n106420), .Q(
        n108183) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][15]  ( .D(n104156), 
        .CK(Clk), .RN(Rst), .Q(n108184) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24794 ), .CK(Clk), .RN(n106469), .Q(n70762) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][15]  ( .D(n104181), 
        .CK(Clk), .RN(n106498), .Q(n108185) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][15]  ( .D(n104162), 
        .CK(Clk), .RN(n106400), .Q(n108186) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24666 ), .CK(Clk), .RN(n106454), .Q(
        n108187), .QN(n103056) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][15]  ( .D(n104172), 
        .CK(Clk), .RN(n106451), .Q(n70767) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24602 ), .CK(Clk), .RN(n106453), .Q(
        n108188) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24538 ), .CK(Clk), .RN(n106383), .Q(
        n108189) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24506 ), .CK(Clk), .RN(n106452), .Q(
        n108190), .QN(n102482) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24474 ), .CK(Clk), .RN(Rst), .Q(n70772), 
        .QN(n104620) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][15]  ( .D(n104144), 
        .CK(Clk), .RN(n106376), .Q(n108191) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24410 ), .CK(Clk), .RN(Rst), .Q(n108192)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][15]  ( .D(n104192), 
        .CK(Clk), .RN(n106450), .Q(n108193) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24346 ), .CK(Clk), .RN(Rst), .Q(n108194)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][15]  ( .D(n104074), 
        .CK(Clk), .RN(Rst), .Q(n108195) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24282 ), .CK(Clk), .RN(n106405), .Q(
        n108196), .QN(n103053) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24250 ), .CK(Clk), .RN(n106413), .Q(
        n108197) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24218 ), .CK(Clk), .RN(n106439), .Q(
        n108198) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24154 ), .CK(Clk), .RN(n106438), .Q(
        n108199) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][15]  ( .D(n104112), 
        .CK(Clk), .RN(n106434), .Q(n108200) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][15]  ( .D(n104083), 
        .CK(Clk), .RN(n106504), .Q(n108201) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24026 ), .CK(Clk), .RN(n106437), .Q(n70786) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23994 ), .CK(Clk), .RN(n106432), .Q(
        n108202), .QN(n101065) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23962 ), .CK(Clk), .RN(n106433), .Q(
        n108203) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][15]  ( .D(n104093), 
        .CK(Clk), .RN(Rst), .Q(n108204), .QN(n103642) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23898 ), .CK(Clk), .RN(n106444), .Q(
        n108205), .QN(n103051) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][15]  ( .D(n104127), 
        .CK(Clk), .RN(Rst), .Q(n108206) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][15]  ( .D(n104020), 
        .CK(Clk), .RN(n106392), .Q(n108207) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23770 ), .CK(Clk), .RN(n106392), .Q(
        n108208), .QN(n101037) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][15]  ( .D(n104036), 
        .CK(Clk), .RN(n106392), .Q(n108209) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23706 ), .CK(Clk), .RN(n106392), .Q(n70796) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23674 ), .CK(Clk), .RN(n106392), .Q(
        n108210), .QN(n101006) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23642 ), .CK(Clk), .RN(n106392), .Q(n70798) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23610 ), .CK(Clk), .RN(n106392), .Q(
        n108211) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23578 ), .CK(Clk), .RN(n106392), .Q(
        n108212) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][15]  ( .D(n104031), 
        .CK(Clk), .RN(n106392), .Q(n108213), .QN(n103638) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23514 ), .CK(Clk), .RN(n106392), .Q(
        n108214) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][15]  ( .D(n104045), 
        .CK(Clk), .RN(n106392), .Q(n70803) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23450 ), .CK(Clk), .RN(n106391), .Q(n70804) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23418 ), .CK(Clk), .RN(n106391), .Q(
        n108215) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23386 ), .CK(Clk), .RN(n106391), .Q(
        n108216) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][15]  ( .D(n104065), 
        .CK(Clk), .RN(n106391), .Q(n108217) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23322 ), .CK(Clk), .RN(n106391), .Q(
        n108218) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][15]  ( .D(n104005), 
        .CK(Clk), .RN(n106391), .Q(n108219) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23258 ), .CK(Clk), .RN(n106391), .Q(
        n108220), .QN(n103049) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23226 ), .CK(Clk), .RN(n106391), .Q(
        n108221) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23194 ), .CK(Clk), .RN(n106391), .Q(
        n108222) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23162 ), .CK(Clk), .RN(n106391), .Q(
        n108223) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23130 ), .CK(Clk), .RN(n106391), .Q(
        n108224) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23098 ), .CK(Clk), .RN(n106391), .Q(
        n108225) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23066 ), .CK(Clk), .RN(n106390), .Q(
        n108226) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23034 ), .CK(Clk), .RN(n106390), .Q(
        n108227) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23002 ), .CK(Clk), .RN(n106390), .Q(
        n108228) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][15]  ( .D(n104015), 
        .CK(Clk), .RN(n106390), .Q(n108229) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22938 ), .CK(Clk), .RN(n106390), .Q(n70820) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][15]  ( .D(n103997), 
        .CK(Clk), .RN(n106390), .Q(n70821) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22874 ), .CK(Clk), .RN(n106390), .Q(
        n108230) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22842 ), .CK(Clk), .RN(n106390), .Q(
        n108231) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22810 ), .CK(Clk), .RN(n106390), .Q(
        n108232) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22778 ), .CK(Clk), .RN(n106390), .Q(
        n108233) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22746 ), .CK(Clk), .RN(n106390), .Q(n70826) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22714 ), .CK(Clk), .RN(n106390), .Q(
        n108234) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22682 ), .CK(Clk), .RN(Rst), .Q(n108235)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22650 ), .CK(Clk), .RN(Rst), .Q(n108236)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22618 ), .CK(Clk), .RN(n106504), .Q(
        n108237) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22586 ), .CK(Clk), .RN(Rst), .Q(n108238)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25882 ), .CK(Clk), .RN(n106413), .Q(n70833) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][15]  ( .D(n104277), 
        .CK(Clk), .RN(n106434), .Q(n108240) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25946 ), .CK(Clk), .RN(n106438), .Q(
        n108241) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25978 ), .CK(Clk), .RN(n106437), .Q(
        n108242), .QN(n103650) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26010 ), .CK(Clk), .RN(n106432), .Q(
        n108243) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][15]  ( .D(n104231), 
        .CK(Clk), .RN(Rst), .Q(n108244) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26074 ), .CK(Clk), .RN(n106433), .Q(
        n108245) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26106 ), .CK(Clk), .RN(Rst), .Q(n70840) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26138 ), .CK(Clk), .RN(Rst), .Q(n108246), 
        .QN(n101923) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26170 ), .CK(Clk), .RN(n106501), .Q(n70842) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26202 ), .CK(Clk), .RN(n106503), .Q(n70843) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26234 ), .CK(Clk), .RN(n106419), .Q(
        n108247) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26266 ), .CK(Clk), .RN(n106480), .Q(n70845) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][15]  ( .D(n104241), 
        .CK(Clk), .RN(n106458), .Q(n108248) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26330 ), .CK(Clk), .RN(n106491), .Q(
        n108249) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26362 ), .CK(Clk), .RN(n106481), .Q(
        n108250) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26394 ), .CK(Clk), .RN(n106456), .Q(
        n108251) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26458 ), .CK(Clk), .RN(n106455), .Q(
        n108253) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26490 ), .CK(Clk), .RN(n106389), .Q(
        n108254), .QN(n103651) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26522 ), .CK(Clk), .RN(n106389), .Q(
        n108255) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26554 ), .CK(Clk), .RN(n106389), .Q(
        n108256) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26586 ), .CK(Clk), .RN(n106389), .Q(
        n108257) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26618 ), .CK(Clk), .RN(n106389), .Q(
        n108258) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][15]  ( .D(n106974), 
        .CK(Clk), .RN(n106389), .Q(n108259) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26682 ), .CK(Clk), .RN(n106389), .Q(
        n108260), .QN(n102491) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26714 ), .CK(Clk), .RN(n106389), .Q(
        n108261), .QN(n103063) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26746 ), .CK(Clk), .RN(n106389), .Q(n70860), .QN(n104540) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][15]  ( .D(n107005), 
        .CK(Clk), .RN(n106389), .Q(n108262), .QN(n101924) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26842 ), .CK(Clk), .RN(n106389), .Q(
        n108264), .QN(n103064) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[15]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107077), .Q(
        \DLX_Datapath/next_A_IDEX[15] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[15]  ( .D(n106621), .CK(Clk), .RN(n106388), 
        .Q(n108265) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[15]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [15]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[15]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [15]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [15]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[15]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [15]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [15]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[15]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107043), .Q(
        \DLX_Datapath/next_B_IDEX [15]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[15]  ( .D(n106693), .CK(Clk), .RN(n106388), 
        .Q(n70872) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[15]  ( .D(n58974), .CK(Clk), .RN(n106388), 
        .Q(n108270) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[15]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [15]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [15]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[15]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [15]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [15]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[15]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N160 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [15]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[14]  ( .D(n106901), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [14]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[14]  ( .D(n104338), .CK(Clk), .RN(
        n106388), .Q(DataAddr[14]), .QN(n58664) );
  DFFR_X2 \DLX_Datapath/PC_reg[14]  ( .D(n60311), .CK(Clk), .RN(n106388), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [2]), .QN(n62199) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[12]  ( .D(n106537), .CK(Clk), .RN(n106388), .Q(n108276) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[12]  ( .D(n106646), .CK(Clk), .RN(n106388), .Q(n70880) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[12]  ( .D(n58971), .CK(Clk), .RN(n106388), .Q(n108277), .QN(n59335) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[13]  ( .D(n106536), .CK(Clk), .RN(n106388), .Q(n108278) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[13]  ( .D(n106656), .CK(Clk), .RN(n106388), .Q(n70882) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[13]  ( .D(n58970), .CK(Clk), .RN(n106388), .Q(n108279), .QN(n59336) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[14]  ( .D(n106535), .CK(Clk), .RN(n106387), .Q(n108280) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[14]  ( .D(n106636), .CK(Clk), .RN(n106387), .Q(n70884) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[14]  ( .D(n58969), .CK(Clk), .RN(n106387), .Q(n108281), .QN(n59337) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25849 ), .CK(Clk), .RN(n106387), .Q(n70888) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25817 ), .CK(Clk), .RN(n106387), .Q(
        n108283) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25785 ), .CK(Clk), .RN(n106387), .Q(
        n108284) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25753 ), .CK(Clk), .RN(n106387), .Q(
        n108285) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25689 ), .CK(Clk), .RN(n106387), .Q(
        n108286) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25625 ), .CK(Clk), .RN(n106386), .Q(
        n108287) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25593 ), .CK(Clk), .RN(n106386), .Q(
        n108288) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25561 ), .CK(Clk), .RN(n106386), .Q(
        n108289) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25529 ), .CK(Clk), .RN(n106386), .Q(
        n108290) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25497 ), .CK(Clk), .RN(n106386), .Q(
        n108291), .QN(n100578) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25465 ), .CK(Clk), .RN(n106386), .Q(n70900) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25433 ), .CK(Clk), .RN(n106386), .Q(
        n108292) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25401 ), .CK(Clk), .RN(n106386), .Q(
        n108293) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25369 ), .CK(Clk), .RN(n106386), .Q(
        n108294) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25337 ), .CK(Clk), .RN(n106386), .Q(
        n108295) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25305 ), .CK(Clk), .RN(n106386), .Q(
        n108296), .QN(n103040) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25273 ), .CK(Clk), .RN(n106386), .Q(
        n108297), .QN(n102471) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25241 ), .CK(Clk), .RN(n106385), .Q(
        n108298), .QN(n101905) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25209 ), .CK(Clk), .RN(n106385), .Q(
        n108299) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25177 ), .CK(Clk), .RN(n106385), .Q(n70909) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][14]  ( .D(n104200), 
        .CK(Clk), .RN(n106385), .Q(n108300) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25081 ), .CK(Clk), .RN(n106385), .Q(
        n108301) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25049 ), .CK(Clk), .RN(n106385), .Q(n70913), .QN(n104598) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][14]  ( .D(n104207), 
        .CK(Clk), .RN(n106385), .Q(n108302) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24985 ), .CK(Clk), .RN(n106385), .Q(
        n108303), .QN(n100610) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24953 ), .CK(Clk), .RN(n106385), .Q(
        n108304) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24921 ), .CK(Clk), .RN(n106385), .Q(n70917) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24889 ), .CK(Clk), .RN(n106385), .Q(
        n108305), .QN(n101165) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24857 ), .CK(Clk), .RN(n106384), .Q(
        n108306) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24825 ), .CK(Clk), .RN(n106384), .Q(
        n108307) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24793 ), .CK(Clk), .RN(n106384), .Q(n70921) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][14]  ( .D(n104184), 
        .CK(Clk), .RN(n106384), .Q(n108308) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24697 ), .CK(Clk), .RN(n106384), .Q(
        n108309) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24665 ), .CK(Clk), .RN(n106384), .Q(
        n108310), .QN(n103036) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][14]  ( .D(n104174), 
        .CK(Clk), .RN(n106384), .Q(n70926) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24601 ), .CK(Clk), .RN(n106384), .Q(
        n108311) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24537 ), .CK(Clk), .RN(n106384), .Q(
        n108312) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24505 ), .CK(Clk), .RN(n106384), .Q(
        n108313), .QN(n102464) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24473 ), .CK(Clk), .RN(n106379), .Q(n70931), .QN(n104619) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24441 ), .CK(Clk), .RN(Rst), .Q(n108314)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24409 ), .CK(Clk), .RN(n106390), .Q(
        n108315) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24377 ), .CK(Clk), .RN(Rst), .Q(n108316)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24345 ), .CK(Clk), .RN(n106391), .Q(
        n108317) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][14]  ( .D(n104100), 
        .CK(Clk), .RN(n106390), .Q(n108318) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24281 ), .CK(Clk), .RN(n106392), .Q(
        n108319), .QN(n103033) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24249 ), .CK(Clk), .RN(n106393), .Q(
        n108320) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24217 ), .CK(Clk), .RN(n106380), .Q(
        n108321) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24153 ), .CK(Clk), .RN(n106455), .Q(
        n108322) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][14]  ( .D(n104121), 
        .CK(Clk), .RN(Rst), .Q(n108323) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][14]  ( .D(n104082), 
        .CK(Clk), .RN(Rst), .Q(n108324) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24025 ), .CK(Clk), .RN(Rst), .Q(n70945) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23993 ), .CK(Clk), .RN(Rst), .Q(n108325), 
        .QN(n102462) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23961 ), .CK(Clk), .RN(Rst), .Q(n108326)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23929 ), .CK(Clk), .RN(Rst), .Q(n108327), 
        .QN(n103624) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23897 ), .CK(Clk), .RN(Rst), .Q(n108328), 
        .QN(n103031) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23865 ), .CK(Clk), .RN(Rst), .Q(n108329)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][14]  ( .D(n104019), 
        .CK(Clk), .RN(Rst), .Q(n108330) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23769 ), .CK(Clk), .RN(Rst), .Q(n108331), 
        .QN(n101038) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][14]  ( .D(n104037), 
        .CK(Clk), .RN(Rst), .Q(n108332) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23705 ), .CK(Clk), .RN(n106388), .Q(n70955) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23673 ), .CK(Clk), .RN(Rst), .Q(n108333), 
        .QN(n101007) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23641 ), .CK(Clk), .RN(Rst), .Q(n70957) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23609 ), .CK(Clk), .RN(Rst), .Q(n108334)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23577 ), .CK(Clk), .RN(Rst), .Q(n108335)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][14]  ( .D(n104030), 
        .CK(Clk), .RN(Rst), .Q(n108336), .QN(n103620) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23513 ), .CK(Clk), .RN(Rst), .Q(n108337)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][14]  ( .D(n104046), 
        .CK(Clk), .RN(Rst), .Q(n70962) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23449 ), .CK(Clk), .RN(Rst), .Q(n70963) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23417 ), .CK(Clk), .RN(Rst), .Q(n108338)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23385 ), .CK(Clk), .RN(Rst), .Q(n108339)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][14]  ( .D(n104069), 
        .CK(Clk), .RN(Rst), .Q(n108340) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23321 ), .CK(Clk), .RN(n106397), .Q(
        n108341) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23289 ), .CK(Clk), .RN(n106397), .Q(
        n108342) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23257 ), .CK(Clk), .RN(n106397), .Q(
        n108343), .QN(n103029) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23225 ), .CK(Clk), .RN(n106397), .Q(
        n108344) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23193 ), .CK(Clk), .RN(n106397), .Q(
        n108345) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23161 ), .CK(Clk), .RN(n106397), .Q(
        n108346) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23129 ), .CK(Clk), .RN(n106397), .Q(
        n108347) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23097 ), .CK(Clk), .RN(n106397), .Q(
        n108348) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23065 ), .CK(Clk), .RN(n106397), .Q(
        n108349) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23033 ), .CK(Clk), .RN(n106397), .Q(
        n108350) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23001 ), .CK(Clk), .RN(n106397), .Q(
        n108351) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22969 ), .CK(Clk), .RN(n106397), .Q(
        n108352) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22937 ), .CK(Clk), .RN(Rst), .Q(n70979) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22905 ), .CK(Clk), .RN(n106371), .Q(n70980) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22873 ), .CK(Clk), .RN(n106490), .Q(
        n108353) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22841 ), .CK(Clk), .RN(Rst), .Q(n108354)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22809 ), .CK(Clk), .RN(Rst), .Q(n108355)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22777 ), .CK(Clk), .RN(Rst), .Q(n108356)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22745 ), .CK(Clk), .RN(Rst), .Q(n70985) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22713 ), .CK(Clk), .RN(Rst), .Q(n108357)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22681 ), .CK(Clk), .RN(Rst), .Q(n108358)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22649 ), .CK(Clk), .RN(Rst), .Q(n108359)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22617 ), .CK(Clk), .RN(Rst), .Q(n108360)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22585 ), .CK(Clk), .RN(n106371), .Q(
        n108361) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25881 ), .CK(Clk), .RN(n106396), .Q(n70992) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][14]  ( .D(n104269), 
        .CK(Clk), .RN(n106396), .Q(n108363) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25945 ), .CK(Clk), .RN(n106396), .Q(
        n108364) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25977 ), .CK(Clk), .RN(n106396), .Q(
        n108365), .QN(n103632) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26009 ), .CK(Clk), .RN(n106396), .Q(
        n108366) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][14]  ( .D(n104230), 
        .CK(Clk), .RN(n106396), .Q(n108367) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26073 ), .CK(Clk), .RN(n106396), .Q(
        n108368) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26105 ), .CK(Clk), .RN(n106396), .Q(n70999) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26137 ), .CK(Clk), .RN(n106396), .Q(
        n108369), .QN(n101907) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26169 ), .CK(Clk), .RN(n106396), .Q(n71001) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26201 ), .CK(Clk), .RN(n106396), .Q(n71002) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26233 ), .CK(Clk), .RN(n106471), .Q(
        n108370) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26265 ), .CK(Clk), .RN(n106470), .Q(n71004) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][14]  ( .D(n104240), 
        .CK(Clk), .RN(n106396), .Q(n108371) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26329 ), .CK(Clk), .RN(n106397), .Q(
        n108372) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26361 ), .CK(Clk), .RN(n106469), .Q(
        n108373) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26393 ), .CK(Clk), .RN(n106468), .Q(
        n108374) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26457 ), .CK(Clk), .RN(n106467), .Q(
        n108376) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26489 ), .CK(Clk), .RN(n106466), .Q(
        n108377), .QN(n103634) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26521 ), .CK(Clk), .RN(n106465), .Q(
        n108378) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26553 ), .CK(Clk), .RN(n106474), .Q(
        n108379) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26585 ), .CK(Clk), .RN(Rst), .Q(n108380)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26617 ), .CK(Clk), .RN(n106404), .Q(
        n108381) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][14]  ( .D(n106973), 
        .CK(Clk), .RN(n106425), .Q(n108382) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26681 ), .CK(Clk), .RN(Rst), .Q(n108383), 
        .QN(n102473) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26713 ), .CK(Clk), .RN(Rst), .Q(n108384), 
        .QN(n103043) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26745 ), .CK(Clk), .RN(Rst), .Q(n71019), 
        .QN(n104539) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][14]  ( .D(n107004), 
        .CK(Clk), .RN(Rst), .Q(n108385), .QN(n101908) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26841 ), .CK(Clk), .RN(n106371), .Q(
        n108387), .QN(n103044) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[14]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107076), .Q(
        \DLX_Datapath/next_A_IDEX[14] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[14]  ( .D(n106607), .CK(Clk), .RN(Rst), .Q(
        n108388) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[14]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [14]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[14]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [14]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [14]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[14]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [14]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [14]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[14]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107042), .Q(
        \DLX_Datapath/next_B_IDEX [14]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[14]  ( .D(n106671), .CK(Clk), .RN(n106371), 
        .Q(n71026) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[14]  ( .D(n58966), .CK(Clk), .RN(Rst), .Q(
        n108391) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[14]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [14]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [14]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[14]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [14]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [14]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[14]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N159 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [14]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[13]  ( .D(n106899), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [13]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[13]  ( .D(n104339), .CK(Clk), .RN(
        n106418), .Q(DataAddr[13]), .QN(n58656) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25848 ), .CK(Clk), .RN(n106395), .Q(n71033) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25816 ), .CK(Clk), .RN(n106395), .Q(
        n108394) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25784 ), .CK(Clk), .RN(n106395), .Q(
        n108395) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25752 ), .CK(Clk), .RN(n106395), .Q(
        n108396) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25688 ), .CK(Clk), .RN(n106395), .Q(
        n108397) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25624 ), .CK(Clk), .RN(n106395), .Q(
        n108398) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25592 ), .CK(Clk), .RN(n106395), .Q(
        n108399) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25560 ), .CK(Clk), .RN(n106395), .Q(
        n108400) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25528 ), .CK(Clk), .RN(n106394), .Q(
        n108401) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25496 ), .CK(Clk), .RN(n106394), .Q(
        n108402), .QN(n100579) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25464 ), .CK(Clk), .RN(n106394), .Q(n71045) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25432 ), .CK(Clk), .RN(n106394), .Q(
        n108403) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25400 ), .CK(Clk), .RN(n106394), .Q(
        n108404) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25368 ), .CK(Clk), .RN(n106394), .Q(
        n108405) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][13]  ( .D(n104302), 
        .CK(Clk), .RN(n106394), .Q(n108406) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25304 ), .CK(Clk), .RN(n106394), .Q(
        n108407), .QN(n103020) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25272 ), .CK(Clk), .RN(n106394), .Q(
        n108408), .QN(n102451) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25240 ), .CK(Clk), .RN(n106394), .Q(
        n108409), .QN(n101889) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25208 ), .CK(Clk), .RN(n106394), .Q(
        n108410) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25176 ), .CK(Clk), .RN(n106394), .Q(n71054) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25144 ), .CK(Clk), .RN(Rst), .Q(n108411)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][13]  ( .D(n104286), 
        .CK(Clk), .RN(Rst), .Q(n108412) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25048 ), .CK(Clk), .RN(Rst), .Q(n71058), 
        .QN(n104597) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][13]  ( .D(n104209), 
        .CK(Clk), .RN(Rst), .Q(n108413) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24984 ), .CK(Clk), .RN(Rst), .Q(n108414), 
        .QN(n100611) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][13]  ( .D(n104296), 
        .CK(Clk), .RN(n106430), .Q(n108415) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24920 ), .CK(Clk), .RN(Rst), .Q(n71062) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24888 ), .CK(Clk), .RN(n106477), .Q(
        n108416), .QN(n101166) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24856 ), .CK(Clk), .RN(Rst), .Q(n108417)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][13]  ( .D(n104155), 
        .CK(Clk), .RN(Rst), .Q(n108418) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24792 ), .CK(Clk), .RN(Rst), .Q(n71066) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][13]  ( .D(n104182), 
        .CK(Clk), .RN(n106494), .Q(n108419) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24696 ), .CK(Clk), .RN(n106409), .Q(
        n108420) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24664 ), .CK(Clk), .RN(n106411), .Q(
        n108421), .QN(n103016) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24632 ), .CK(Clk), .RN(n106410), .Q(n71071) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24600 ), .CK(Clk), .RN(Rst), .Q(n108422)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24536 ), .CK(Clk), .RN(n106409), .Q(
        n108423) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24504 ), .CK(Clk), .RN(n106411), .Q(
        n108424), .QN(n102444) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24472 ), .CK(Clk), .RN(n106508), .Q(n71076), .QN(n104618) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][13]  ( .D(n104148), 
        .CK(Clk), .RN(n106493), .Q(n108425) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24408 ), .CK(Clk), .RN(n106410), .Q(
        n108426) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][13]  ( .D(n104197), 
        .CK(Clk), .RN(Rst), .Q(n108427) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24344 ), .CK(Clk), .RN(Rst), .Q(n108428)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][13]  ( .D(n104111), 
        .CK(Clk), .RN(Rst), .Q(n108429) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24280 ), .CK(Clk), .RN(Rst), .Q(n108430), 
        .QN(n103013) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24248 ), .CK(Clk), .RN(Rst), .Q(n108431)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24216 ), .CK(Clk), .RN(Rst), .Q(n108432)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24152 ), .CK(Clk), .RN(Rst), .Q(n108433)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][13]  ( .D(n104113), 
        .CK(Clk), .RN(Rst), .Q(n108434) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][13]  ( .D(n104081), 
        .CK(Clk), .RN(Rst), .Q(n108435) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24024 ), .CK(Clk), .RN(Rst), .Q(n71090) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23992 ), .CK(Clk), .RN(Rst), .Q(n108436), 
        .QN(n101066) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23960 ), .CK(Clk), .RN(Rst), .Q(n108437)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][13]  ( .D(n104092), 
        .CK(Clk), .RN(Rst), .Q(n108438), .QN(n103605) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23896 ), .CK(Clk), .RN(Rst), .Q(n108439), 
        .QN(n103011) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][13]  ( .D(n104128), 
        .CK(Clk), .RN(Rst), .Q(n108440) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][13]  ( .D(n104018), 
        .CK(Clk), .RN(Rst), .Q(n108441) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23768 ), .CK(Clk), .RN(n106473), .Q(
        n108442), .QN(n101039) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][13]  ( .D(n104035), 
        .CK(Clk), .RN(Rst), .Q(n108443) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23704 ), .CK(Clk), .RN(Rst), .Q(n71100) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23672 ), .CK(Clk), .RN(Rst), .Q(n108444), 
        .QN(n101008) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23640 ), .CK(Clk), .RN(Rst), .Q(n71102) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23608 ), .CK(Clk), .RN(n106393), .Q(
        n108445) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23576 ), .CK(Clk), .RN(n106393), .Q(
        n108446) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][13]  ( .D(n104029), 
        .CK(Clk), .RN(n106393), .Q(n108447), .QN(n103601) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23512 ), .CK(Clk), .RN(n106393), .Q(
        n108448) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][13]  ( .D(n104044), 
        .CK(Clk), .RN(n106393), .Q(n71107) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23448 ), .CK(Clk), .RN(n106393), .Q(n71108) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23416 ), .CK(Clk), .RN(n106393), .Q(
        n108449) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23384 ), .CK(Clk), .RN(n106393), .Q(
        n108450) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][13]  ( .D(n104066), 
        .CK(Clk), .RN(n106393), .Q(n108451) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23320 ), .CK(Clk), .RN(n106393), .Q(
        n108452) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][13]  ( .D(n104000), 
        .CK(Clk), .RN(n106393), .Q(n108453) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23256 ), .CK(Clk), .RN(n106393), .Q(
        n108454), .QN(n103009) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23224 ), .CK(Clk), .RN(n106395), .Q(
        n108455) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23192 ), .CK(Clk), .RN(Rst), .Q(n108456)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23160 ), .CK(Clk), .RN(Rst), .Q(n108457)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23128 ), .CK(Clk), .RN(Rst), .Q(n108458)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][13]  ( .D(n104011), 
        .CK(Clk), .RN(Rst), .Q(n108459) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23064 ), .CK(Clk), .RN(Rst), .Q(n108460)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23032 ), .CK(Clk), .RN(Rst), .Q(n108461)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23000 ), .CK(Clk), .RN(Rst), .Q(n108462)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][13]  ( .D(n104013), 
        .CK(Clk), .RN(Rst), .Q(n108463) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22936 ), .CK(Clk), .RN(Rst), .Q(n71124) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][13]  ( .D(n103996), 
        .CK(Clk), .RN(Rst), .Q(n71125) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22872 ), .CK(Clk), .RN(Rst), .Q(n108464)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22840 ), .CK(Clk), .RN(Rst), .Q(n108465)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22808 ), .CK(Clk), .RN(Rst), .Q(n108466)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22776 ), .CK(Clk), .RN(Rst), .Q(n108467)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22744 ), .CK(Clk), .RN(Rst), .Q(n71130) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22712 ), .CK(Clk), .RN(Rst), .Q(n108468)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22680 ), .CK(Clk), .RN(Rst), .Q(n108469)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22648 ), .CK(Clk), .RN(Rst), .Q(n108470)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22616 ), .CK(Clk), .RN(Rst), .Q(n108471)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22584 ), .CK(Clk), .RN(Rst), .Q(n108472)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25880 ), .CK(Clk), .RN(Rst), .Q(n71137) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][13]  ( .D(n104275), 
        .CK(Clk), .RN(Rst), .Q(n108474) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25944 ), .CK(Clk), .RN(Rst), .Q(n108475)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25976 ), .CK(Clk), .RN(Rst), .Q(n108476), 
        .QN(n103614) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26008 ), .CK(Clk), .RN(Rst), .Q(n108477)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][13]  ( .D(n104229), 
        .CK(Clk), .RN(Rst), .Q(n108478) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26072 ), .CK(Clk), .RN(Rst), .Q(n108479)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26104 ), .CK(Clk), .RN(Rst), .Q(n71144) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26136 ), .CK(Clk), .RN(Rst), .Q(n108480), 
        .QN(n101891) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26168 ), .CK(Clk), .RN(Rst), .Q(n71146) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26200 ), .CK(Clk), .RN(Rst), .Q(n71147) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26232 ), .CK(Clk), .RN(Rst), .Q(n108481)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26264 ), .CK(Clk), .RN(Rst), .Q(n71149) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][13]  ( .D(n104239), 
        .CK(Clk), .RN(Rst), .Q(n108482) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26328 ), .CK(Clk), .RN(Rst), .Q(n108483)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26360 ), .CK(Clk), .RN(n106376), .Q(
        n108484) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26392 ), .CK(Clk), .RN(n106400), .Q(
        n108485) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26456 ), .CK(Clk), .RN(n106451), .Q(
        n108487) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26488 ), .CK(Clk), .RN(n106450), .Q(
        n108488), .QN(n103616) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26520 ), .CK(Clk), .RN(Rst), .Q(n108489)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26552 ), .CK(Clk), .RN(Rst), .Q(n108490)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26584 ), .CK(Clk), .RN(Rst), .Q(n108491)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26616 ), .CK(Clk), .RN(Rst), .Q(n108492)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][13]  ( .D(n106972), 
        .CK(Clk), .RN(Rst), .Q(n108493) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26680 ), .CK(Clk), .RN(n106487), .Q(
        n108494), .QN(n102453) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26712 ), .CK(Clk), .RN(n106461), .Q(
        n108495), .QN(n103023) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26744 ), .CK(Clk), .RN(n106415), .Q(n71164), .QN(n104538) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][13]  ( .D(n107003), 
        .CK(Clk), .RN(Rst), .Q(n108496), .QN(n101892) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26840 ), .CK(Clk), .RN(Rst), .Q(n108498), 
        .QN(n103024) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[13]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107075), .Q(
        \DLX_Datapath/next_A_IDEX[13] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[13]  ( .D(n106606), .CK(Clk), .RN(n106404), 
        .Q(n108499) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[13]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107041), .Q(
        \DLX_Datapath/next_B_IDEX [13]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[13]  ( .D(n106692), .CK(Clk), .RN(Rst), .Q(
        n71169) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[13]  ( .D(n58963), .CK(Clk), .RN(n106408), 
        .Q(n108500) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[13]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [13]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[11]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N124 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [11]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[11]  ( .D(n106897), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [11]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[11]  ( .D(n104340), .CK(Clk), .RN(
        n106384), .Q(DataAddr[11]), .QN(n58653) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[11]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [11]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [11]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[11]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [11]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [11]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[11]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N156 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [11]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[10]  ( .D(n106895), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [10]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[10]  ( .D(n104341), .CK(Clk), .RN(
        n106374), .Q(DataAddr[10]), .QN(n58651) );
  DFFR_X2 \DLX_Datapath/PC_reg[10]  ( .D(n60315), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [2]), .QN(n104581) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[10]  ( .D(n106539), .CK(Clk), .RN(Rst), 
        .Q(n108508) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[10]  ( .D(n106645), .CK(Clk), .RN(n106427), .Q(n71179) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[10]  ( .D(n58958), .CK(Clk), .RN(n106403), .Q(n108509), .QN(n59333) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25845 ), .CK(Clk), .RN(Rst), .Q(n71182) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25813 ), .CK(Clk), .RN(Rst), .Q(n108511)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][10]  ( .D(n104215), 
        .CK(Clk), .RN(Rst), .Q(n108512) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25749 ), .CK(Clk), .RN(Rst), .Q(n108513)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25685 ), .CK(Clk), .RN(Rst), .Q(n108514)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25621 ), .CK(Clk), .RN(n106428), .Q(
        n108515) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25589 ), .CK(Clk), .RN(n106402), .Q(
        n108516), .QN(n103559) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25557 ), .CK(Clk), .RN(n106443), .Q(
        n108517) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25525 ), .CK(Clk), .RN(n106486), .Q(
        n108518) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25493 ), .CK(Clk), .RN(n106429), .Q(
        n108519), .QN(n100582) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25461 ), .CK(Clk), .RN(n106418), .Q(n71194) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25429 ), .CK(Clk), .RN(n106425), .Q(
        n108520) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25397 ), .CK(Clk), .RN(n106490), .Q(
        n108521) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25365 ), .CK(Clk), .RN(n106488), .Q(
        n108522) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][10]  ( .D(n104301), 
        .CK(Clk), .RN(n106484), .Q(n108523) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25301 ), .CK(Clk), .RN(Rst), .Q(n108524), 
        .QN(n102963) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25269 ), .CK(Clk), .RN(n106441), .Q(
        n108525), .QN(n102393) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25237 ), .CK(Clk), .RN(n106397), .Q(
        n108526), .QN(n101837) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25205 ), .CK(Clk), .RN(n106377), .Q(
        n108527) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25173 ), .CK(Clk), .RN(n106377), .Q(n71203) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][10]  ( .D(n104203), 
        .CK(Clk), .RN(n106377), .Q(n108528) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][10]  ( .D(n104281), 
        .CK(Clk), .RN(n106377), .Q(n108529) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25045 ), .CK(Clk), .RN(n106377), .Q(n71207), .QN(n104594) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][10]  ( .D(n104211), 
        .CK(Clk), .RN(n106377), .Q(n108530) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24981 ), .CK(Clk), .RN(n106377), .Q(
        n108531), .QN(n100614) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][10]  ( .D(n104292), 
        .CK(Clk), .RN(n106377), .Q(n108532) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24917 ), .CK(Clk), .RN(n106377), .Q(n71211) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24885 ), .CK(Clk), .RN(n106377), .Q(
        n108533), .QN(n101169) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24853 ), .CK(Clk), .RN(n106377), .Q(
        n108534) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][10]  ( .D(n104153), 
        .CK(Clk), .RN(n106376), .Q(n108535) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24789 ), .CK(Clk), .RN(n106376), .Q(n71215) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][10]  ( .D(n104185), 
        .CK(Clk), .RN(n106376), .Q(n108536) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][10]  ( .D(n104160), 
        .CK(Clk), .RN(n106376), .Q(n108537) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24661 ), .CK(Clk), .RN(n106376), .Q(
        n108538), .QN(n102959) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][10]  ( .D(n104175), 
        .CK(Clk), .RN(n106376), .Q(n71220) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24597 ), .CK(Clk), .RN(n106376), .Q(
        n108539) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24533 ), .CK(Clk), .RN(n106376), .Q(
        n108540) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24501 ), .CK(Clk), .RN(n106376), .Q(
        n108541), .QN(n102386) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24469 ), .CK(Clk), .RN(n106376), .Q(n71225), .QN(n104647) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][10]  ( .D(n104143), 
        .CK(Clk), .RN(Rst), .Q(n108542) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24405 ), .CK(Clk), .RN(Rst), .Q(n108543)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][10]  ( .D(n104196), 
        .CK(Clk), .RN(Rst), .Q(n108544) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24341 ), .CK(Clk), .RN(Rst), .Q(n108545)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][10]  ( .D(n104101), 
        .CK(Clk), .RN(Rst), .Q(n108546) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24277 ), .CK(Clk), .RN(Rst), .Q(n108547), 
        .QN(n102956) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24245 ), .CK(Clk), .RN(Rst), .Q(n108548)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24213 ), .CK(Clk), .RN(Rst), .Q(n108549)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24149 ), .CK(Clk), .RN(Rst), .Q(n108550)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][10]  ( .D(n104119), 
        .CK(Clk), .RN(Rst), .Q(n108551) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][10]  ( .D(n104076), 
        .CK(Clk), .RN(n106375), .Q(n108552), .QN(n103552) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24021 ), .CK(Clk), .RN(n106375), .Q(n71239) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23989 ), .CK(Clk), .RN(n106375), .Q(
        n108553), .QN(n102384) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23957 ), .CK(Clk), .RN(n106375), .Q(
        n108554) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][10]  ( .D(n104087), 
        .CK(Clk), .RN(n106375), .Q(n108555) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23893 ), .CK(Clk), .RN(n106375), .Q(
        n108556), .QN(n102954) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][10]  ( .D(n104125), 
        .CK(Clk), .RN(n106375), .Q(n108557) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23797 ), .CK(Clk), .RN(n106375), .Q(
        n108558) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23765 ), .CK(Clk), .RN(n106375), .Q(
        n108559), .QN(n101042) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][10]  ( .D(n104038), 
        .CK(Clk), .RN(n106375), .Q(n108560) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23701 ), .CK(Clk), .RN(n106375), .Q(n71249) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23669 ), .CK(Clk), .RN(n106374), .Q(
        n108561) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23637 ), .CK(Clk), .RN(n106374), .Q(n71251) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23605 ), .CK(Clk), .RN(n106374), .Q(
        n108562) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23573 ), .CK(Clk), .RN(n106374), .Q(
        n108563) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][10]  ( .D(n104027), 
        .CK(Clk), .RN(n106374), .Q(n108564), .QN(n103548) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23509 ), .CK(Clk), .RN(n106374), .Q(
        n108565) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][10]  ( .D(n104052), 
        .CK(Clk), .RN(n106374), .Q(n71256) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23445 ), .CK(Clk), .RN(n106374), .Q(n71257) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23413 ), .CK(Clk), .RN(n106374), .Q(
        n108566) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23381 ), .CK(Clk), .RN(n106374), .Q(
        n108567) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][10]  ( .D(n104072), 
        .CK(Clk), .RN(n106374), .Q(n108568) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23317 ), .CK(Clk), .RN(n106374), .Q(
        n108569) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23253 ), .CK(Clk), .RN(n106373), .Q(
        n108570), .QN(n102952) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23221 ), .CK(Clk), .RN(n106373), .Q(
        n108571) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23189 ), .CK(Clk), .RN(n106373), .Q(
        n108572) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23125 ), .CK(Clk), .RN(n106373), .Q(
        n108573) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23093 ), .CK(Clk), .RN(n106373), .Q(
        n108574) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23061 ), .CK(Clk), .RN(n106373), .Q(
        n108575) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23029 ), .CK(Clk), .RN(n106373), .Q(
        n108576) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22997 ), .CK(Clk), .RN(n106373), .Q(
        n108577) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][10]  ( .D(n104014), 
        .CK(Clk), .RN(n106373), .Q(n108578) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22933 ), .CK(Clk), .RN(n106502), .Q(n71273) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][10]  ( .D(n103995), 
        .CK(Clk), .RN(n106383), .Q(n71274) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22869 ), .CK(Clk), .RN(n106383), .Q(
        n108579) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22837 ), .CK(Clk), .RN(n106383), .Q(
        n108580) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22805 ), .CK(Clk), .RN(n106383), .Q(
        n108581) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22773 ), .CK(Clk), .RN(n106383), .Q(
        n108582) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22741 ), .CK(Clk), .RN(n106383), .Q(n71279) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22709 ), .CK(Clk), .RN(n106383), .Q(
        n108583) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22677 ), .CK(Clk), .RN(n106383), .Q(
        n108584) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22645 ), .CK(Clk), .RN(n106383), .Q(
        n108585) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22613 ), .CK(Clk), .RN(n106383), .Q(
        n108586) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22581 ), .CK(Clk), .RN(n106383), .Q(
        n108587) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][10]  ( .D(
        \DLX_Datapath/RegisterFile/N22549 ), .CK(Clk), .RN(Rst), .Q(n71285), 
        .QN(n104521) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25877 ), .CK(Clk), .RN(Rst), .Q(n71286) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][10]  ( .D(n104268), 
        .CK(Clk), .RN(Rst), .Q(n108588) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25941 ), .CK(Clk), .RN(Rst), .Q(n108589)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25973 ), .CK(Clk), .RN(Rst), .Q(n108590)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26005 ), .CK(Clk), .RN(Rst), .Q(n108591)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][10]  ( .D(n104227), 
        .CK(Clk), .RN(Rst), .Q(n108592) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26069 ), .CK(Clk), .RN(Rst), .Q(n108593)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26101 ), .CK(Clk), .RN(Rst), .Q(n71293), 
        .QN(n104615) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26133 ), .CK(Clk), .RN(Rst), .Q(n108594), 
        .QN(n101841) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26165 ), .CK(Clk), .RN(Rst), .Q(n71295) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26197 ), .CK(Clk), .RN(Rst), .Q(n71296) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26229 ), .CK(Clk), .RN(Rst), .Q(n108595)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26261 ), .CK(Clk), .RN(Rst), .Q(n71298) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][10]  ( .D(n104237), 
        .CK(Clk), .RN(Rst), .Q(n108596) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26325 ), .CK(Clk), .RN(Rst), .Q(n108597)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26357 ), .CK(Clk), .RN(Rst), .Q(n108598)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26389 ), .CK(Clk), .RN(Rst), .Q(n108599)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26453 ), .CK(Clk), .RN(Rst), .Q(n108601)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26485 ), .CK(Clk), .RN(Rst), .Q(n108602), 
        .QN(n103562) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26517 ), .CK(Clk), .RN(Rst), .Q(n108603)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26549 ), .CK(Clk), .RN(Rst), .Q(n108604)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26581 ), .CK(Clk), .RN(Rst), .Q(n108605)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26613 ), .CK(Clk), .RN(Rst), .Q(n108606)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][10]  ( .D(n106969), 
        .CK(Clk), .RN(Rst), .Q(n108607) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26677 ), .CK(Clk), .RN(Rst), .Q(n108608), 
        .QN(n102395) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26709 ), .CK(Clk), .RN(Rst), .Q(n108609), 
        .QN(n102966) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26741 ), .CK(Clk), .RN(Rst), .Q(n71313), 
        .QN(n104535) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][10]  ( .D(n107000), 
        .CK(Clk), .RN(Rst), .Q(n108610), .QN(n101842) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26837 ), .CK(Clk), .RN(Rst), .Q(n108612), 
        .QN(n102967) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[10]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107072), .Q(
        \DLX_Datapath/next_A_IDEX[10] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[10]  ( .D(n106605), .CK(Clk), .RN(Rst), .Q(
        n108613) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[10]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [10]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[3]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N116 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [3]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[3]  ( .D(n106885), .GN(n106360), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [3]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[3]  ( .D(n104342), .CK(Clk), .RN(Rst), 
        .Q(DataAddr[3]), .QN(n58647) );
  DFFR_X2 \DLX_Datapath/PC_reg[3]  ( .D(n60322), .CK(Clk), .RN(Rst), .Q(
        PC_out[3]), .QN(net2465244) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[0]  ( .D(n60293), .CK(Clk), .RN(Rst), .Q(
        n108615) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[1]  ( .D(n60292), .CK(Clk), .RN(Rst), .Q(
        n108616) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[2]  ( .D(n60291), .CK(Clk), .RN(n106373), 
        .Q(n108617) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[3]  ( .D(n60290), .CK(Clk), .RN(n106393), 
        .Q(n108618) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[1]  ( .D(n106548), .CK(Clk), .RN(Rst), 
        .Q(n108619), .QN(n100460) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[1]  ( .D(n106642), .CK(Clk), .RN(n106473), 
        .Q(n71325) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[1]  ( .D(n58954), .CK(Clk), .RN(Rst), 
        .Q(n108620), .QN(n100413) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[2]  ( .D(n106547), .CK(Clk), .RN(n106475), 
        .Q(n108621) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[2]  ( .D(n106653), .CK(Clk), .RN(n106457), 
        .Q(n71327) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[2]  ( .D(n58953), .CK(Clk), .RN(Rst), 
        .Q(n108622), .QN(n58643) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[3]  ( .D(n106546), .CK(Clk), .RN(n106392), 
        .Q(n108631) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[3]  ( .D(n106632), .CK(Clk), .RN(n106391), 
        .Q(n71329) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[3]  ( .D(n58952), .CK(Clk), .RN(Rst), 
        .Q(n108632), .QN(n100799) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25838 ), .CK(Clk), .RN(n106382), .Q(n71331) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25806 ), .CK(Clk), .RN(n106382), .Q(
        n108633) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][3]  ( .D(n104219), 
        .CK(Clk), .RN(n106382), .Q(n108634) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25742 ), .CK(Clk), .RN(n106382), .Q(
        n108635) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25678 ), .CK(Clk), .RN(n106382), .Q(
        n108636) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25614 ), .CK(Clk), .RN(n106382), .Q(
        n108637) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25582 ), .CK(Clk), .RN(n106382), .Q(
        n108638) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25550 ), .CK(Clk), .RN(n106382), .Q(
        n108639) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25518 ), .CK(Clk), .RN(n106382), .Q(
        n108640) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25486 ), .CK(Clk), .RN(n106381), .Q(
        n108641), .QN(n100589) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25454 ), .CK(Clk), .RN(n106381), .Q(n71343) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25422 ), .CK(Clk), .RN(n106381), .Q(
        n108642) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25390 ), .CK(Clk), .RN(n106381), .Q(
        n108643) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25358 ), .CK(Clk), .RN(n106381), .Q(
        n108644) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25326 ), .CK(Clk), .RN(n106381), .Q(
        n108645) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25294 ), .CK(Clk), .RN(n106381), .Q(
        n108646), .QN(n102823) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25262 ), .CK(Clk), .RN(n106381), .Q(
        n108647), .QN(n102256) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25230 ), .CK(Clk), .RN(n106381), .Q(
        n108648), .QN(n101715) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25198 ), .CK(Clk), .RN(n106381), .Q(
        n108649) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25166 ), .CK(Clk), .RN(n106381), .Q(n71352) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25134 ), .CK(Clk), .RN(n106380), .Q(
        n108650) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25070 ), .CK(Clk), .RN(n106380), .Q(
        n108651) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25038 ), .CK(Clk), .RN(n106380), .Q(n71356), .QN(n104587) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][3]  ( .D(n104212), 
        .CK(Clk), .RN(n106380), .Q(n108652) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24974 ), .CK(Clk), .RN(n106380), .Q(
        n108653), .QN(n100621) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24942 ), .CK(Clk), .RN(n106380), .Q(
        n108654) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24910 ), .CK(Clk), .RN(n106380), .Q(n71360) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24878 ), .CK(Clk), .RN(n106380), .Q(
        n108655), .QN(n101176) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24846 ), .CK(Clk), .RN(n106380), .Q(
        n108656) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24814 ), .CK(Clk), .RN(n106380), .Q(
        n108657) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24782 ), .CK(Clk), .RN(n106380), .Q(n71364) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][3]  ( .D(n104189), 
        .CK(Clk), .RN(n106379), .Q(n108658) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24686 ), .CK(Clk), .RN(n106379), .Q(
        n108659) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24654 ), .CK(Clk), .RN(n106379), .Q(
        n108660), .QN(n102819) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][3]  ( .D(n104178), 
        .CK(Clk), .RN(n106379), .Q(n71369) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24590 ), .CK(Clk), .RN(n106379), .Q(
        n108661) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24526 ), .CK(Clk), .RN(n106379), .Q(
        n108662) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24494 ), .CK(Clk), .RN(n106379), .Q(
        n108663), .QN(n102249) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24462 ), .CK(Clk), .RN(n106379), .Q(n71374), .QN(n104640) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24430 ), .CK(Clk), .RN(n106379), .Q(
        n108664) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24398 ), .CK(Clk), .RN(n106379), .Q(
        n108665) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][3]  ( .D(n104193), 
        .CK(Clk), .RN(n106378), .Q(n108666) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24334 ), .CK(Clk), .RN(n106378), .Q(
        n108667) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24302 ), .CK(Clk), .RN(n106378), .Q(
        n108668) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24270 ), .CK(Clk), .RN(n106378), .Q(
        n108669), .QN(n102816) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24238 ), .CK(Clk), .RN(n106378), .Q(
        n108670) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24206 ), .CK(Clk), .RN(n106378), .Q(
        n108671) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24142 ), .CK(Clk), .RN(n106378), .Q(
        n108672) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24110 ), .CK(Clk), .RN(n106378), .Q(
        n108673) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24046 ), .CK(Clk), .RN(n106378), .Q(
        n108674) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24014 ), .CK(Clk), .RN(n106378), .Q(n71388) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23982 ), .CK(Clk), .RN(Rst), .Q(n108675), 
        .QN(n102247) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23950 ), .CK(Clk), .RN(Rst), .Q(n108676)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23918 ), .CK(Clk), .RN(Rst), .Q(n108677), 
        .QN(n103418) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23886 ), .CK(Clk), .RN(Rst), .Q(n108678), 
        .QN(n102814) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23854 ), .CK(Clk), .RN(Rst), .Q(n108679)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23790 ), .CK(Clk), .RN(Rst), .Q(n108680)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23758 ), .CK(Clk), .RN(Rst), .Q(n108681), 
        .QN(n101049) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23726 ), .CK(Clk), .RN(Rst), .Q(n108682)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23694 ), .CK(Clk), .RN(Rst), .Q(n71398) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23662 ), .CK(Clk), .RN(Rst), .Q(n108683), 
        .QN(n101017) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23630 ), .CK(Clk), .RN(Rst), .Q(n71400) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23598 ), .CK(Clk), .RN(Rst), .Q(n108684)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23566 ), .CK(Clk), .RN(Rst), .Q(n108685)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23534 ), .CK(Clk), .RN(Rst), .Q(n108686), 
        .QN(n103414) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23502 ), .CK(Clk), .RN(Rst), .Q(n108687)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][3]  ( .D(n104058), 
        .CK(Clk), .RN(n106420), .Q(n71405) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23438 ), .CK(Clk), .RN(n106492), .Q(n71406) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23406 ), .CK(Clk), .RN(Rst), .Q(n108688)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23374 ), .CK(Clk), .RN(Rst), .Q(n108689)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][3]  ( .D(n104073), 
        .CK(Clk), .RN(n106372), .Q(n108690) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23310 ), .CK(Clk), .RN(Rst), .Q(n108691)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23278 ), .CK(Clk), .RN(n106442), .Q(
        n108692) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23246 ), .CK(Clk), .RN(Rst), .Q(n108693), 
        .QN(n102812) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23214 ), .CK(Clk), .RN(Rst), .Q(n108694)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23182 ), .CK(Clk), .RN(n106506), .Q(
        n108695) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23150 ), .CK(Clk), .RN(Rst), .Q(n108696)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23118 ), .CK(Clk), .RN(Rst), .Q(n108697)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23086 ), .CK(Clk), .RN(Rst), .Q(n108698)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23054 ), .CK(Clk), .RN(n106493), .Q(
        n108699) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23022 ), .CK(Clk), .RN(Rst), .Q(n108700)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22990 ), .CK(Clk), .RN(Rst), .Q(n108701)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22958 ), .CK(Clk), .RN(Rst), .Q(n108702)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22926 ), .CK(Clk), .RN(n106494), .Q(n71422) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22894 ), .CK(Clk), .RN(Rst), .Q(n71423) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22862 ), .CK(Clk), .RN(Rst), .Q(n108703)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22830 ), .CK(Clk), .RN(n106381), .Q(
        n108704) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22798 ), .CK(Clk), .RN(n106383), .Q(
        n108705) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22766 ), .CK(Clk), .RN(Rst), .Q(n108706)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22734 ), .CK(Clk), .RN(Rst), .Q(n71428) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22670 ), .CK(Clk), .RN(Rst), .Q(n108707)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22638 ), .CK(Clk), .RN(Rst), .Q(n108708)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22606 ), .CK(Clk), .RN(Rst), .Q(n108709)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22574 ), .CK(Clk), .RN(Rst), .Q(n108710)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22542 ), .CK(Clk), .RN(Rst), .Q(n71434), 
        .QN(n104515) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25870 ), .CK(Clk), .RN(Rst), .Q(n71435) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][3]  ( .D(n104253), 
        .CK(Clk), .RN(Rst), .Q(n108711) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25934 ), .CK(Clk), .RN(Rst), .Q(n108712)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25966 ), .CK(Clk), .RN(Rst), .Q(n108713), 
        .QN(n103427) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25998 ), .CK(Clk), .RN(n106422), .Q(
        n108714) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][3]  ( .D(n104235), 
        .CK(Clk), .RN(n106422), .Q(n108715) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26062 ), .CK(Clk), .RN(n106422), .Q(
        n108716) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26094 ), .CK(Clk), .RN(n106422), .Q(n71442) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26126 ), .CK(Clk), .RN(n106422), .Q(
        n108717), .QN(n101719) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26158 ), .CK(Clk), .RN(n106422), .Q(n71444) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26190 ), .CK(Clk), .RN(n106422), .Q(n71445) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26222 ), .CK(Clk), .RN(n106422), .Q(
        n108718) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26254 ), .CK(Clk), .RN(n106422), .Q(n71447) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26286 ), .CK(Clk), .RN(n106422), .Q(
        n108719) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26318 ), .CK(Clk), .RN(n106422), .Q(
        n108720) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26350 ), .CK(Clk), .RN(n106422), .Q(
        n108721) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26382 ), .CK(Clk), .RN(n106421), .Q(
        n108722) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26446 ), .CK(Clk), .RN(n106421), .Q(
        n108724) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26478 ), .CK(Clk), .RN(n106421), .Q(
        n108725), .QN(n103429) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26510 ), .CK(Clk), .RN(n106421), .Q(
        n108726) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26542 ), .CK(Clk), .RN(n106421), .Q(
        n108727) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26574 ), .CK(Clk), .RN(n106421), .Q(
        n108728) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26606 ), .CK(Clk), .RN(n106421), .Q(
        n108729) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][3]  ( .D(n106962), 
        .CK(Clk), .RN(n106421), .Q(n108730) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26670 ), .CK(Clk), .RN(n106421), .Q(
        n108731), .QN(n102258) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26702 ), .CK(Clk), .RN(n106421), .Q(
        n108732), .QN(n102826) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26734 ), .CK(Clk), .RN(n106421), .Q(n71462), .QN(n104530) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][3]  ( .D(n106993), 
        .CK(Clk), .RN(n106420), .Q(n108733), .QN(n101720) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26830 ), .CK(Clk), .RN(n106420), .Q(
        n108735), .QN(n102827) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[3]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107065), .Q(
        \DLX_Datapath/next_A_IDEX[3] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[3]  ( .D(n106601), .CK(Clk), .RN(n106420), 
        .Q(n108736) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[3]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [3]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[3]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [3]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [3]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[3]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [3]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [3]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[3]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107031), .Q(
        \DLX_Datapath/next_B_IDEX [3]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[3]  ( .D(n106665), .CK(Clk), .RN(n106420), 
        .Q(n71469) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[3]  ( .D(n58948), .CK(Clk), .RN(n106420), 
        .Q(n108739) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[3]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [3]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [3]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[3]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [3]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [3]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_shf_reg[3]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [3]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/B_shf [3]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[3]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N148 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [3]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[0]  ( .D(n104359), .GN(n60159), 
        .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [0]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[1]  ( .D(n106881), .GN(n106360), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [1]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[1]  ( .D(n104343), .CK(Clk), .RN(
        n106420), .Q(DataAddr[1]), .QN(n58635) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25836 ), .CK(Clk), .RN(n106420), .Q(n71482) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25804 ), .CK(Clk), .RN(n106420), .Q(
        n108748) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][1]  ( .D(n104218), 
        .CK(Clk), .RN(n106420), .Q(n108749) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25740 ), .CK(Clk), .RN(n106420), .Q(
        n108750) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25676 ), .CK(Clk), .RN(Rst), .Q(n108751)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25612 ), .CK(Clk), .RN(Rst), .Q(n108752)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25580 ), .CK(Clk), .RN(Rst), .Q(n108753)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25548 ), .CK(Clk), .RN(Rst), .Q(n108754)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25516 ), .CK(Clk), .RN(Rst), .Q(n108755)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25484 ), .CK(Clk), .RN(n106467), .Q(
        n108756), .QN(n100591) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25452 ), .CK(Clk), .RN(n106468), .Q(n71494) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25420 ), .CK(Clk), .RN(n106469), .Q(
        n108757) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25388 ), .CK(Clk), .RN(n106397), .Q(
        n108758) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25356 ), .CK(Clk), .RN(n106429), .Q(
        n108759) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][1]  ( .D(n104310), 
        .CK(Clk), .RN(n106419), .Q(n108760) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25292 ), .CK(Clk), .RN(n106419), .Q(
        n108761), .QN(n102783) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25260 ), .CK(Clk), .RN(n106419), .Q(
        n108762), .QN(n102217) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25228 ), .CK(Clk), .RN(n106419), .Q(
        n108763), .QN(n101679) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25196 ), .CK(Clk), .RN(n106419), .Q(
        n108764) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25164 ), .CK(Clk), .RN(n106419), .Q(n71503) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25132 ), .CK(Clk), .RN(n106419), .Q(
        n108765) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][1]  ( .D(n104280), 
        .CK(Clk), .RN(n106419), .Q(n108766) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25036 ), .CK(Clk), .RN(n106419), .Q(n71507), .QN(n104585) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][1]  ( .D(n104214), 
        .CK(Clk), .RN(n106419), .Q(n108767) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24972 ), .CK(Clk), .RN(n106419), .Q(
        n108768), .QN(n100623) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][1]  ( .D(n104289), 
        .CK(Clk), .RN(n106418), .Q(n108769) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24908 ), .CK(Clk), .RN(n106418), .Q(n71511) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24876 ), .CK(Clk), .RN(n106418), .Q(
        n108770), .QN(n101178) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24844 ), .CK(Clk), .RN(n106418), .Q(
        n108771) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24812 ), .CK(Clk), .RN(n106418), .Q(
        n108772) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24780 ), .CK(Clk), .RN(n106418), .Q(n71515) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][1]  ( .D(n104187), 
        .CK(Clk), .RN(n106418), .Q(n108773) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][1]  ( .D(n104166), 
        .CK(Clk), .RN(n106418), .Q(n108774) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24652 ), .CK(Clk), .RN(n106418), .Q(
        n108775), .QN(n102779) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][1]  ( .D(n104179), 
        .CK(Clk), .RN(n106418), .Q(n71520) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24588 ), .CK(Clk), .RN(n106417), .Q(
        n108776) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24524 ), .CK(Clk), .RN(n106417), .Q(
        n108777) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24492 ), .CK(Clk), .RN(n106417), .Q(
        n108778), .QN(n102210) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24460 ), .CK(Clk), .RN(n106417), .Q(n71525), .QN(n104638) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][1]  ( .D(n104142), 
        .CK(Clk), .RN(n106417), .Q(n108779) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24396 ), .CK(Clk), .RN(n106417), .Q(
        n108780) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][1]  ( .D(n104191), 
        .CK(Clk), .RN(n106417), .Q(n108781) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24332 ), .CK(Clk), .RN(n106417), .Q(
        n108782) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][1]  ( .D(n104109), 
        .CK(Clk), .RN(n106417), .Q(n108783) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24268 ), .CK(Clk), .RN(n106417), .Q(
        n108784), .QN(n102776) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24236 ), .CK(Clk), .RN(n106417), .Q(
        n108785) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24204 ), .CK(Clk), .RN(Rst), .Q(n108786)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24140 ), .CK(Clk), .RN(Rst), .Q(n108787)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][1]  ( .D(n104118), 
        .CK(Clk), .RN(Rst), .Q(n108788) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][1]  ( .D(n104085), 
        .CK(Clk), .RN(Rst), .Q(n108789) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24012 ), .CK(Clk), .RN(Rst), .Q(n71539) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23980 ), .CK(Clk), .RN(Rst), .Q(n108790), 
        .QN(n102208) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23948 ), .CK(Clk), .RN(Rst), .Q(n108791)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][1]  ( .D(n104097), 
        .CK(Clk), .RN(Rst), .Q(n108792), .QN(n103378) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23884 ), .CK(Clk), .RN(Rst), .Q(n108793), 
        .QN(n102774) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][1]  ( .D(n104130), 
        .CK(Clk), .RN(Rst), .Q(n108794) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][1]  ( .D(n104023), 
        .CK(Clk), .RN(n106416), .Q(n108795) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23756 ), .CK(Clk), .RN(n106416), .Q(
        n108796), .QN(n101051) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][1]  ( .D(n104042), 
        .CK(Clk), .RN(n106416), .Q(n108797) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23692 ), .CK(Clk), .RN(n106416), .Q(n71549) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23660 ), .CK(Clk), .RN(n106416), .Q(
        n108798), .QN(n101019) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23628 ), .CK(Clk), .RN(n106416), .Q(n71551) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23596 ), .CK(Clk), .RN(n106416), .Q(
        n108799) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23564 ), .CK(Clk), .RN(n106416), .Q(
        n108800) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][1]  ( .D(n104032), 
        .CK(Clk), .RN(n106416), .Q(n108801), .QN(n103374) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23500 ), .CK(Clk), .RN(n106416), .Q(
        n108802) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][1]  ( .D(n104059), 
        .CK(Clk), .RN(n106416), .Q(n71556) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23436 ), .CK(Clk), .RN(n106415), .Q(n71557) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23404 ), .CK(Clk), .RN(n106415), .Q(
        n108803) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23372 ), .CK(Clk), .RN(n106415), .Q(
        n108804) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][1]  ( .D(n104071), 
        .CK(Clk), .RN(n106415), .Q(n108805) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23308 ), .CK(Clk), .RN(n106415), .Q(
        n108806) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][1]  ( .D(n104003), 
        .CK(Clk), .RN(n106415), .Q(n108807) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23244 ), .CK(Clk), .RN(n106415), .Q(
        n108808), .QN(n102772) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23212 ), .CK(Clk), .RN(n106415), .Q(
        n108809) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23180 ), .CK(Clk), .RN(n106415), .Q(
        n108810) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23148 ), .CK(Clk), .RN(n106415), .Q(
        n108811) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23116 ), .CK(Clk), .RN(n106415), .Q(
        n108812) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23084 ), .CK(Clk), .RN(n106415), .Q(
        n108813) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23052 ), .CK(Clk), .RN(n106414), .Q(
        n108814) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23020 ), .CK(Clk), .RN(n106414), .Q(
        n108815) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22988 ), .CK(Clk), .RN(n106414), .Q(
        n108816) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][1]  ( .D(n104017), 
        .CK(Clk), .RN(n106414), .Q(n108817) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22924 ), .CK(Clk), .RN(n106414), .Q(n71573) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][1]  ( .D(n103998), 
        .CK(Clk), .RN(n106414), .Q(n71574) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22860 ), .CK(Clk), .RN(n106414), .Q(
        n108818) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22828 ), .CK(Clk), .RN(n106414), .Q(
        n108819) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22796 ), .CK(Clk), .RN(n106414), .Q(
        n108820) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22764 ), .CK(Clk), .RN(n106414), .Q(
        n108821) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22732 ), .CK(Clk), .RN(n106414), .Q(n71579) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22700 ), .CK(Clk), .RN(n106414), .Q(
        n108822) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22668 ), .CK(Clk), .RN(Rst), .Q(n108823)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][1]  ( .D(n103955), 
        .CK(Clk), .RN(Rst), .Q(n108824) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22604 ), .CK(Clk), .RN(Rst), .Q(n108825)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22572 ), .CK(Clk), .RN(Rst), .Q(n108826)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][1]  ( .D(
        \DLX_Datapath/RegisterFile/N22540 ), .CK(Clk), .RN(Rst), .Q(n71585), 
        .QN(n104513) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25868 ), .CK(Clk), .RN(Rst), .Q(n71586) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][1]  ( .D(n104256), 
        .CK(Clk), .RN(Rst), .Q(n108827) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25932 ), .CK(Clk), .RN(Rst), .Q(n108828)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25964 ), .CK(Clk), .RN(Rst), .Q(n108829), 
        .QN(n103387) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25996 ), .CK(Clk), .RN(Rst), .Q(n108830)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][1]  ( .D(n104233), 
        .CK(Clk), .RN(Rst), .Q(n108831) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26060 ), .CK(Clk), .RN(Rst), .Q(n108832)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26092 ), .CK(Clk), .RN(n106418), .Q(n71593) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26124 ), .CK(Clk), .RN(Rst), .Q(n108833), 
        .QN(n101683) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26156 ), .CK(Clk), .RN(n106423), .Q(n71595) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26188 ), .CK(Clk), .RN(Rst), .Q(n71596) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26220 ), .CK(Clk), .RN(n106424), .Q(
        n108834) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26252 ), .CK(Clk), .RN(Rst), .Q(n71598) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26284 ), .CK(Clk), .RN(n106474), .Q(
        n108835) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26316 ), .CK(Clk), .RN(n106441), .Q(
        n108836) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26348 ), .CK(Clk), .RN(n106420), .Q(
        n108837) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26380 ), .CK(Clk), .RN(n106421), .Q(
        n108838) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26444 ), .CK(Clk), .RN(n106422), .Q(
        n108840) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26476 ), .CK(Clk), .RN(Rst), .Q(n108841), 
        .QN(n103389) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26508 ), .CK(Clk), .RN(Rst), .Q(n108842)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26540 ), .CK(Clk), .RN(Rst), .Q(n108843)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26572 ), .CK(Clk), .RN(Rst), .Q(n108844)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26604 ), .CK(Clk), .RN(Rst), .Q(n108845)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][1]  ( .D(n106960), 
        .CK(Clk), .RN(Rst), .Q(n108846) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26668 ), .CK(Clk), .RN(Rst), .Q(n108847), 
        .QN(n102219) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26700 ), .CK(Clk), .RN(Rst), .Q(n108848), 
        .QN(n102786) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26732 ), .CK(Clk), .RN(Rst), .Q(n71613), 
        .QN(n104529) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][1]  ( .D(n106991), 
        .CK(Clk), .RN(Rst), .Q(n108849), .QN(n101684) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26828 ), .CK(Clk), .RN(Rst), .Q(n108851), 
        .QN(n102787) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[1]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107063), .Q(
        \DLX_Datapath/next_A_IDEX[1] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[1]  ( .D(n106600), .CK(Clk), .RN(n106428), 
        .Q(n108853) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[1]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107029), .Q(
        \DLX_Datapath/next_B_IDEX [1]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[1]  ( .D(n106675), .CK(Clk), .RN(n106428), 
        .Q(n71618) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[1]  ( .D(n58945), .CK(Clk), .RN(n106428), 
        .Q(n108854) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[1]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [1]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[1]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [1]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [1]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[1]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [1]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [1]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[1]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [1]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [1]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[0]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N113 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [0]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[1]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N114 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [1]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[1]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [1]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [1]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_shf_reg[1]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [1]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/B_shf [1]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[1]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N146 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [1]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[1]  ( .D(n107575), .GN(n60159), 
        .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [1]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[2]  ( .D(n106883), .GN(n106360), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [2]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[2]  ( .D(n104344), .CK(Clk), .RN(
        n106428), .Q(DataAddr[2]), .QN(n58632) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25837 ), .CK(Clk), .RN(n106428), .Q(n71626) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25805 ), .CK(Clk), .RN(n106428), .Q(
        n108860) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][2]  ( .D(n104220), 
        .CK(Clk), .RN(n106428), .Q(n108861) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25741 ), .CK(Clk), .RN(n106428), .Q(
        n108862) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25677 ), .CK(Clk), .RN(n106428), .Q(
        n108863) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25613 ), .CK(Clk), .RN(n106476), .Q(
        n108864) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25581 ), .CK(Clk), .RN(n106417), .Q(
        n108865) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25549 ), .CK(Clk), .RN(Rst), .Q(n108866)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25517 ), .CK(Clk), .RN(n106416), .Q(
        n108867) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25485 ), .CK(Clk), .RN(n106415), .Q(
        n108868), .QN(n100590) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25453 ), .CK(Clk), .RN(n106414), .Q(n71638) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25421 ), .CK(Clk), .RN(Rst), .Q(n108869)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25389 ), .CK(Clk), .RN(n106413), .Q(
        n108870) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25357 ), .CK(Clk), .RN(n106507), .Q(
        n108871) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25325 ), .CK(Clk), .RN(n106412), .Q(
        n108872) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25293 ), .CK(Clk), .RN(n106411), .Q(
        n108873), .QN(n102803) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25261 ), .CK(Clk), .RN(n106395), .Q(
        n108874), .QN(n102237) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25229 ), .CK(Clk), .RN(n106427), .Q(
        n108875), .QN(n101697) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25197 ), .CK(Clk), .RN(n106427), .Q(
        n108876) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25165 ), .CK(Clk), .RN(n106427), .Q(n71647) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25133 ), .CK(Clk), .RN(n106427), .Q(
        n108877) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25069 ), .CK(Clk), .RN(n106427), .Q(
        n108878) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25037 ), .CK(Clk), .RN(n106427), .Q(n71651), .QN(n104586) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][2]  ( .D(n104205), 
        .CK(Clk), .RN(n106427), .Q(n108879) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24973 ), .CK(Clk), .RN(n106427), .Q(
        n108880), .QN(n100622) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24941 ), .CK(Clk), .RN(n106427), .Q(
        n108881) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24909 ), .CK(Clk), .RN(n106427), .Q(n71655) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24877 ), .CK(Clk), .RN(n106427), .Q(
        n108882), .QN(n101177) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24845 ), .CK(Clk), .RN(Rst), .Q(n108883)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24813 ), .CK(Clk), .RN(Rst), .Q(n108884)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24781 ), .CK(Clk), .RN(Rst), .Q(n71659) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24749 ), .CK(Clk), .RN(Rst), .Q(n108885)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24685 ), .CK(Clk), .RN(Rst), .Q(n108886)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24653 ), .CK(Clk), .RN(Rst), .Q(n108887), 
        .QN(n102799) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][2]  ( .D(n104171), 
        .CK(Clk), .RN(Rst), .Q(n71664) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24589 ), .CK(Clk), .RN(Rst), .Q(n108888)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24525 ), .CK(Clk), .RN(Rst), .Q(n108889)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24493 ), .CK(Clk), .RN(Rst), .Q(n108890), 
        .QN(n102230) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24461 ), .CK(Clk), .RN(n106426), .Q(n71669), .QN(n104639) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24429 ), .CK(Clk), .RN(n106426), .Q(
        n108891) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24397 ), .CK(Clk), .RN(n106426), .Q(
        n108892) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24365 ), .CK(Clk), .RN(n106426), .Q(
        n108893) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24333 ), .CK(Clk), .RN(n106426), .Q(
        n108894) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24301 ), .CK(Clk), .RN(n106426), .Q(
        n108895) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24269 ), .CK(Clk), .RN(n106426), .Q(
        n108896), .QN(n102796) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24237 ), .CK(Clk), .RN(n106426), .Q(
        n108897) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24205 ), .CK(Clk), .RN(n106426), .Q(
        n108898) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24141 ), .CK(Clk), .RN(n106426), .Q(
        n108899) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][2]  ( .D(n104114), 
        .CK(Clk), .RN(n106425), .Q(n108900) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24045 ), .CK(Clk), .RN(n106425), .Q(
        n108901) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24013 ), .CK(Clk), .RN(n106425), .Q(n71683) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23981 ), .CK(Clk), .RN(n106425), .Q(
        n108902), .QN(n102228) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23949 ), .CK(Clk), .RN(n106425), .Q(
        n108903) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23917 ), .CK(Clk), .RN(n106425), .Q(
        n108904), .QN(n103398) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23885 ), .CK(Clk), .RN(n106425), .Q(
        n108905), .QN(n102794) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][2]  ( .D(n104123), 
        .CK(Clk), .RN(n106425), .Q(n108906) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23789 ), .CK(Clk), .RN(n106425), .Q(
        n108907) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23757 ), .CK(Clk), .RN(n106425), .Q(
        n108908), .QN(n101050) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23725 ), .CK(Clk), .RN(n106471), .Q(
        n108909) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23693 ), .CK(Clk), .RN(n106435), .Q(n71693) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23661 ), .CK(Clk), .RN(n106396), .Q(
        n108910), .QN(n101018) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23629 ), .CK(Clk), .RN(n106440), .Q(n71695) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23597 ), .CK(Clk), .RN(n106470), .Q(
        n108911) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23565 ), .CK(Clk), .RN(n106489), .Q(
        n108912) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23533 ), .CK(Clk), .RN(Rst), .Q(n108913), 
        .QN(n103394) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23501 ), .CK(Clk), .RN(n106442), .Q(
        n108914) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23469 ), .CK(Clk), .RN(Rst), .Q(n71700) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23437 ), .CK(Clk), .RN(n106464), .Q(n71701) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23405 ), .CK(Clk), .RN(n106463), .Q(
        n108915) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23373 ), .CK(Clk), .RN(n106462), .Q(
        n108916) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23341 ), .CK(Clk), .RN(Rst), .Q(n108917)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23309 ), .CK(Clk), .RN(Rst), .Q(n108918)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23277 ), .CK(Clk), .RN(Rst), .Q(n108919)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23245 ), .CK(Clk), .RN(Rst), .Q(n108920), 
        .QN(n102792) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23213 ), .CK(Clk), .RN(Rst), .Q(n108921)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23181 ), .CK(Clk), .RN(Rst), .Q(n108922)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23149 ), .CK(Clk), .RN(Rst), .Q(n108923)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23117 ), .CK(Clk), .RN(Rst), .Q(n108924)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23085 ), .CK(Clk), .RN(Rst), .Q(n108925)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23053 ), .CK(Clk), .RN(Rst), .Q(n108926)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23021 ), .CK(Clk), .RN(Rst), .Q(n108927)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22989 ), .CK(Clk), .RN(Rst), .Q(n108928)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22957 ), .CK(Clk), .RN(n106424), .Q(
        n108929) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22925 ), .CK(Clk), .RN(n106424), .Q(n71717) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22893 ), .CK(Clk), .RN(n106424), .Q(n71718) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22861 ), .CK(Clk), .RN(n106424), .Q(
        n108930) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22829 ), .CK(Clk), .RN(n106424), .Q(
        n108931) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22797 ), .CK(Clk), .RN(n106424), .Q(
        n108932) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22765 ), .CK(Clk), .RN(n106424), .Q(
        n108933) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22733 ), .CK(Clk), .RN(n106424), .Q(n71723) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22701 ), .CK(Clk), .RN(n106424), .Q(
        n108934) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22669 ), .CK(Clk), .RN(n106424), .Q(
        n108935) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22637 ), .CK(Clk), .RN(n106424), .Q(
        n108936) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22605 ), .CK(Clk), .RN(n106424), .Q(
        n108937) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][2]  ( .D(n104323), 
        .CK(Clk), .RN(Rst), .Q(n108938) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][2]  ( .D(
        \DLX_Datapath/RegisterFile/N22541 ), .CK(Clk), .RN(Rst), .Q(n71729), 
        .QN(n104514) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25869 ), .CK(Clk), .RN(Rst), .Q(n71730) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][2]  ( .D(n104254), 
        .CK(Clk), .RN(Rst), .Q(n108939) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25933 ), .CK(Clk), .RN(Rst), .Q(n108940)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][2]  ( .D(n104316), 
        .CK(Clk), .RN(Rst), .Q(n108941), .QN(n103407) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25997 ), .CK(Clk), .RN(Rst), .Q(n108942)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][2]  ( .D(n104234), 
        .CK(Clk), .RN(Rst), .Q(n108943) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26061 ), .CK(Clk), .RN(Rst), .Q(n108944)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26093 ), .CK(Clk), .RN(Rst), .Q(n71737) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26125 ), .CK(Clk), .RN(Rst), .Q(n108945), 
        .QN(n101701) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26157 ), .CK(Clk), .RN(Rst), .Q(n71739) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26189 ), .CK(Clk), .RN(n106423), .Q(n71740) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26221 ), .CK(Clk), .RN(n106423), .Q(
        n108946) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26253 ), .CK(Clk), .RN(n106423), .Q(n71742) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26285 ), .CK(Clk), .RN(n106423), .Q(
        n108947) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26317 ), .CK(Clk), .RN(n106423), .Q(
        n108948) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26349 ), .CK(Clk), .RN(n106423), .Q(
        n108949) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26381 ), .CK(Clk), .RN(n106423), .Q(
        n108950) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26445 ), .CK(Clk), .RN(n106423), .Q(
        n108952) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26477 ), .CK(Clk), .RN(n106423), .Q(
        n108953), .QN(n103409) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26509 ), .CK(Clk), .RN(n106423), .Q(
        n108954) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26541 ), .CK(Clk), .RN(n106423), .Q(
        n108955) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26573 ), .CK(Clk), .RN(n106426), .Q(
        n108956) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26605 ), .CK(Clk), .RN(n106404), .Q(
        n108957) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][2]  ( .D(n106961), 
        .CK(Clk), .RN(n106404), .Q(n108958) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26669 ), .CK(Clk), .RN(n106404), .Q(
        n108959), .QN(n102239) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26701 ), .CK(Clk), .RN(n106404), .Q(
        n108960), .QN(n102806) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][2]  ( .D(n104320), 
        .CK(Clk), .RN(n106404), .Q(n71757), .QN(n104527) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][2]  ( .D(n106992), 
        .CK(Clk), .RN(n106404), .Q(n108961), .QN(n101702) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26829 ), .CK(Clk), .RN(n106404), .Q(
        n108963), .QN(n102807) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[2]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107064), .Q(
        \DLX_Datapath/next_A_IDEX[2] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[2]  ( .D(n106615), .CK(Clk), .RN(n106404), 
        .Q(n108964) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[2]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107030), .Q(
        \DLX_Datapath/next_B_IDEX [2]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[2]  ( .D(n106664), .CK(Clk), .RN(n106404), 
        .Q(n71762) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[2]  ( .D(n58942), .CK(Clk), .RN(n106404), 
        .Q(n108965) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[2]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [2]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[2]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [2]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [2]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[2]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [2]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [2]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[2]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [2]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [2]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[2]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N115 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [2]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[2]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [2]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [2]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_shf_reg[2]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [2]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/B_shf [2]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[2]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N147 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [2]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[2]  ( .D(n107576), .GN(n60159), 
        .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [2]) );
  DFFR_X2 \DLX_Datapath/PC_IFID_reg[3]  ( .D(n60226), .CK(Clk), .RN(n106404), 
        .Q(n108971), .QN(n59422) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[3]  ( .D(n107577), .GN(n60159), 
        .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [3]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[7]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N120 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [7]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[7]  ( .D(n106891), .GN(n106360), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [7]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[7]  ( .D(n104345), .CK(Clk), .RN(
        n106403), .Q(DataAddr[7]), .QN(n58629) );
  DFFR_X2 \DLX_Datapath/PC_reg[7]  ( .D(n60318), .CK(Clk), .RN(n106403), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [3]), .QN(n62183) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[7]  ( .D(n106542), .CK(Clk), .RN(n106403), 
        .Q(n108972) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[7]  ( .D(n106644), .CK(Clk), .RN(n106403), 
        .Q(n71772) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[7]  ( .D(n58939), .CK(Clk), .RN(n106403), 
        .Q(n108973), .QN(n59330) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25842 ), .CK(Clk), .RN(n106403), .Q(n71775) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25810 ), .CK(Clk), .RN(n106403), .Q(
        n108976) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25778 ), .CK(Clk), .RN(n106403), .Q(
        n108977) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25746 ), .CK(Clk), .RN(n106403), .Q(
        n108978) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25682 ), .CK(Clk), .RN(n106402), .Q(
        n108979) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25618 ), .CK(Clk), .RN(n106402), .Q(
        n108980) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25586 ), .CK(Clk), .RN(n106402), .Q(
        n108981) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25554 ), .CK(Clk), .RN(n106402), .Q(
        n108982) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25522 ), .CK(Clk), .RN(n106402), .Q(
        n108983) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25490 ), .CK(Clk), .RN(n106402), .Q(
        n108984), .QN(n100585) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25458 ), .CK(Clk), .RN(n106402), .Q(n71787) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25426 ), .CK(Clk), .RN(n106402), .Q(
        n108985) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25394 ), .CK(Clk), .RN(n106402), .Q(
        n108986) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25362 ), .CK(Clk), .RN(n106402), .Q(
        n108987) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25330 ), .CK(Clk), .RN(n106402), .Q(
        n108988) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25298 ), .CK(Clk), .RN(n106401), .Q(
        n108989), .QN(n102903) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25266 ), .CK(Clk), .RN(n106401), .Q(
        n108990), .QN(n102335) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25234 ), .CK(Clk), .RN(n106401), .Q(
        n108991), .QN(n101785) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25202 ), .CK(Clk), .RN(n106401), .Q(
        n108992) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25170 ), .CK(Clk), .RN(n106401), .Q(n71796) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25138 ), .CK(Clk), .RN(n106401), .Q(
        n108993) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25074 ), .CK(Clk), .RN(n106401), .Q(
        n108994) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25042 ), .CK(Clk), .RN(n106401), .Q(n71800), .QN(n104591) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25010 ), .CK(Clk), .RN(n106401), .Q(
        n108995) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24978 ), .CK(Clk), .RN(n106401), .Q(
        n108996), .QN(n100617) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24946 ), .CK(Clk), .RN(n106401), .Q(
        n108997) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24914 ), .CK(Clk), .RN(n106400), .Q(n71804) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24882 ), .CK(Clk), .RN(n106400), .Q(
        n108998), .QN(n101172) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24850 ), .CK(Clk), .RN(n106400), .Q(
        n108999) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24818 ), .CK(Clk), .RN(n106400), .Q(
        n109000) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24786 ), .CK(Clk), .RN(n106400), .Q(n71808) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24754 ), .CK(Clk), .RN(n106400), .Q(
        n109001) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24690 ), .CK(Clk), .RN(n106400), .Q(
        n109002) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24658 ), .CK(Clk), .RN(n106400), .Q(
        n109003), .QN(n102899) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][7]  ( .D(n104176), 
        .CK(Clk), .RN(n106400), .Q(n71813) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24594 ), .CK(Clk), .RN(n106400), .Q(
        n109004) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24530 ), .CK(Clk), .RN(Rst), .Q(n109005)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24498 ), .CK(Clk), .RN(Rst), .Q(n109006), 
        .QN(n102328) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24466 ), .CK(Clk), .RN(Rst), .Q(n71818), 
        .QN(n104644) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24434 ), .CK(Clk), .RN(Rst), .Q(n109007)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24402 ), .CK(Clk), .RN(Rst), .Q(n109008)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24370 ), .CK(Clk), .RN(Rst), .Q(n109009)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24338 ), .CK(Clk), .RN(Rst), .Q(n109010)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24306 ), .CK(Clk), .RN(Rst), .Q(n109011)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24274 ), .CK(Clk), .RN(Rst), .Q(n109012), 
        .QN(n102896) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24242 ), .CK(Clk), .RN(Rst), .Q(n109013)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24210 ), .CK(Clk), .RN(Rst), .Q(n109014)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24146 ), .CK(Clk), .RN(n106399), .Q(
        n109015) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24114 ), .CK(Clk), .RN(n106399), .Q(
        n109016) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24050 ), .CK(Clk), .RN(n106399), .Q(
        n109017) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24018 ), .CK(Clk), .RN(n106399), .Q(n71832) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23986 ), .CK(Clk), .RN(n106399), .Q(
        n109018), .QN(n102326) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23954 ), .CK(Clk), .RN(n106399), .Q(
        n109019) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23922 ), .CK(Clk), .RN(n106399), .Q(
        n109020), .QN(n103496) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23890 ), .CK(Clk), .RN(n106399), .Q(
        n109021), .QN(n102894) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23858 ), .CK(Clk), .RN(n106399), .Q(
        n109022) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23794 ), .CK(Clk), .RN(n106475), .Q(
        n109023) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23762 ), .CK(Clk), .RN(n106393), .Q(
        n109024), .QN(n101045) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23730 ), .CK(Clk), .RN(n106392), .Q(
        n109025) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23698 ), .CK(Clk), .RN(n106391), .Q(n71842) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23666 ), .CK(Clk), .RN(n106390), .Q(
        n109026), .QN(n101014) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23634 ), .CK(Clk), .RN(n106405), .Q(n71844) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23602 ), .CK(Clk), .RN(Rst), .Q(n109027)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23570 ), .CK(Clk), .RN(n106389), .Q(
        n109028) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23538 ), .CK(Clk), .RN(n106388), .Q(
        n109029), .QN(n103492) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23506 ), .CK(Clk), .RN(n106403), .Q(
        n109030) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23474 ), .CK(Clk), .RN(n106410), .Q(n71849) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23442 ), .CK(Clk), .RN(Rst), .Q(n71850) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23410 ), .CK(Clk), .RN(Rst), .Q(n109031)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23378 ), .CK(Clk), .RN(Rst), .Q(n109032)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23346 ), .CK(Clk), .RN(Rst), .Q(n109033)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23314 ), .CK(Clk), .RN(Rst), .Q(n109034)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23282 ), .CK(Clk), .RN(Rst), .Q(n109035)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23250 ), .CK(Clk), .RN(Rst), .Q(n109036), 
        .QN(n102892) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23218 ), .CK(Clk), .RN(Rst), .Q(n109037)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23186 ), .CK(Clk), .RN(Rst), .Q(n109038)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23154 ), .CK(Clk), .RN(Rst), .Q(n109039)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23122 ), .CK(Clk), .RN(Rst), .Q(n109040)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23090 ), .CK(Clk), .RN(Rst), .Q(n109041)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23058 ), .CK(Clk), .RN(Rst), .Q(n109042)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23026 ), .CK(Clk), .RN(n106398), .Q(
        n109043) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22994 ), .CK(Clk), .RN(n106398), .Q(
        n109044) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22962 ), .CK(Clk), .RN(n106398), .Q(
        n109045) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22930 ), .CK(Clk), .RN(n106398), .Q(n71866) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22898 ), .CK(Clk), .RN(n106398), .Q(n71867) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22866 ), .CK(Clk), .RN(n106398), .Q(
        n109046) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22834 ), .CK(Clk), .RN(n106398), .Q(
        n109047) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22802 ), .CK(Clk), .RN(n106398), .Q(
        n109048) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22770 ), .CK(Clk), .RN(n106398), .Q(
        n109049) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22738 ), .CK(Clk), .RN(n106398), .Q(n71872) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22706 ), .CK(Clk), .RN(n106398), .Q(
        n109050) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22674 ), .CK(Clk), .RN(n106398), .Q(
        n109051) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22642 ), .CK(Clk), .RN(Rst), .Q(n109052)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][7]  ( .D(
        \DLX_Datapath/RegisterFile/N22610 ), .CK(Clk), .RN(Rst), .Q(n109053), 
        .QN(n101624) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][7]  ( .D(n104324), 
        .CK(Clk), .RN(Rst), .Q(n109054), .QN(n102318) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25874 ), .CK(Clk), .RN(Rst), .Q(n71879) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][7]  ( .D(n104255), 
        .CK(Clk), .RN(Rst), .Q(n109056) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25938 ), .CK(Clk), .RN(Rst), .Q(n109057)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25970 ), .CK(Clk), .RN(Rst), .Q(n109058), 
        .QN(n103505) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26002 ), .CK(Clk), .RN(Rst), .Q(n109059)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26034 ), .CK(Clk), .RN(Rst), .Q(n109060)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26066 ), .CK(Clk), .RN(Rst), .Q(n109061)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26098 ), .CK(Clk), .RN(Rst), .Q(n71886) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26130 ), .CK(Clk), .RN(Rst), .Q(n109062), 
        .QN(n101789) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26162 ), .CK(Clk), .RN(Rst), .Q(n71888) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26194 ), .CK(Clk), .RN(Rst), .Q(n71889) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26226 ), .CK(Clk), .RN(Rst), .Q(n109063)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26258 ), .CK(Clk), .RN(Rst), .Q(n71891) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26290 ), .CK(Clk), .RN(Rst), .Q(n109064)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26322 ), .CK(Clk), .RN(Rst), .Q(n109065)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26354 ), .CK(Clk), .RN(Rst), .Q(n109066)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26386 ), .CK(Clk), .RN(Rst), .Q(n109067)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26450 ), .CK(Clk), .RN(Rst), .Q(n109069)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26482 ), .CK(Clk), .RN(Rst), .Q(n109070), 
        .QN(n103507) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26514 ), .CK(Clk), .RN(Rst), .Q(n109071)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26546 ), .CK(Clk), .RN(Rst), .Q(n109072)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26578 ), .CK(Clk), .RN(Rst), .Q(n109073)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26610 ), .CK(Clk), .RN(Rst), .Q(n109074)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][7]  ( .D(n106966), 
        .CK(Clk), .RN(Rst), .Q(n109075) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26674 ), .CK(Clk), .RN(Rst), .Q(n109076), 
        .QN(n102337) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26706 ), .CK(Clk), .RN(Rst), .Q(n109077), 
        .QN(n102906) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26738 ), .CK(Clk), .RN(Rst), .Q(n71906), 
        .QN(n104533) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][7]  ( .D(n106997), 
        .CK(Clk), .RN(Rst), .Q(n109078), .QN(n101790) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26834 ), .CK(Clk), .RN(Rst), .Q(n109080), 
        .QN(n102907) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[7]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107069), .Q(
        \DLX_Datapath/next_A_IDEX[7] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[7]  ( .D(n106603), .CK(Clk), .RN(Rst), .Q(
        n109081) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[7]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [7]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[7]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [7]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [7]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[7]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [7]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [7]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[7]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107035), .Q(
        \DLX_Datapath/next_B_IDEX [7]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[7]  ( .D(n106689), .CK(Clk), .RN(n106399), 
        .Q(n71913) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[7]  ( .D(n58937), .CK(Clk), .RN(n106413), 
        .Q(n109084) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[7]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [7]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [7]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[7]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [7]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [7]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[7]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N152 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [7]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[4]  ( .D(n104360), .GN(n60159), 
        .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [4]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[5]  ( .D(n107612), .GN(n60159), 
        .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [5]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[6]  ( .D(n106889), .GN(n106360), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [6]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[6]  ( .D(n104346), .CK(Clk), .RN(
        n106413), .Q(DataAddr[6]), .QN(n58624) );
  DFFR_X2 \DLX_Datapath/PC_reg[6]  ( .D(n60319), .CK(Clk), .RN(n106413), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [2]), .QN(n62200) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[4]  ( .D(n106545), .CK(Clk), .RN(n106413), 
        .Q(n109092) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[4]  ( .D(n106654), .CK(Clk), .RN(n106413), 
        .Q(n71922) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[4]  ( .D(n58934), .CK(Clk), .RN(n106413), 
        .Q(n109093), .QN(n59327) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[5]  ( .D(n106544), .CK(Clk), .RN(n106413), 
        .Q(n109094) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[5]  ( .D(n106643), .CK(Clk), .RN(n106413), 
        .Q(n71924) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[5]  ( .D(n58933), .CK(Clk), .RN(n106413), 
        .Q(n109095), .QN(n59328) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[6]  ( .D(n106543), .CK(Clk), .RN(n106413), 
        .Q(n109096) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[6]  ( .D(n106633), .CK(Clk), .RN(n106413), 
        .Q(n71926) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[6]  ( .D(n58932), .CK(Clk), .RN(n106485), 
        .Q(n109097), .QN(n59329) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25839 ), .CK(Clk), .RN(n106401), .Q(n71929) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25807 ), .CK(Clk), .RN(n106466), .Q(
        n109098) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25775 ), .CK(Clk), .RN(n106465), .Q(
        n109099) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25743 ), .CK(Clk), .RN(Rst), .Q(n109100)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25679 ), .CK(Clk), .RN(Rst), .Q(n109101)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25615 ), .CK(Clk), .RN(Rst), .Q(n109102)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25583 ), .CK(Clk), .RN(n106460), .Q(
        n109103) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25551 ), .CK(Clk), .RN(n106398), .Q(
        n109104) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25519 ), .CK(Clk), .RN(n106412), .Q(
        n109105) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25487 ), .CK(Clk), .RN(n106412), .Q(
        n109106), .QN(n100588) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25455 ), .CK(Clk), .RN(n106412), .Q(n71941) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25423 ), .CK(Clk), .RN(n106412), .Q(
        n109107) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25391 ), .CK(Clk), .RN(n106412), .Q(
        n109108) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25359 ), .CK(Clk), .RN(n106412), .Q(
        n109109) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25327 ), .CK(Clk), .RN(n106412), .Q(
        n109110) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25295 ), .CK(Clk), .RN(n106412), .Q(
        n109111), .QN(n102843) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25263 ), .CK(Clk), .RN(n106412), .Q(
        n109112), .QN(n102276) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25231 ), .CK(Clk), .RN(n106412), .Q(
        n109113), .QN(n101733) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25199 ), .CK(Clk), .RN(n106412), .Q(
        n109114) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25167 ), .CK(Clk), .RN(n106412), .Q(n71950) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25135 ), .CK(Clk), .RN(n106411), .Q(
        n109115) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25071 ), .CK(Clk), .RN(n106411), .Q(
        n109116) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25039 ), .CK(Clk), .RN(n106411), .Q(n71954), .QN(n104588) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25007 ), .CK(Clk), .RN(n106411), .Q(
        n109117) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24975 ), .CK(Clk), .RN(n106411), .Q(
        n109118), .QN(n100620) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24943 ), .CK(Clk), .RN(n106411), .Q(
        n109119) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24911 ), .CK(Clk), .RN(n106411), .Q(n71958) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24879 ), .CK(Clk), .RN(n106411), .Q(
        n109120), .QN(n101175) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24847 ), .CK(Clk), .RN(n106411), .Q(
        n109121) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24815 ), .CK(Clk), .RN(n106411), .Q(
        n109122) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24783 ), .CK(Clk), .RN(n106411), .Q(n71962) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24751 ), .CK(Clk), .RN(n106410), .Q(
        n109123) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24687 ), .CK(Clk), .RN(n106410), .Q(
        n109124) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24655 ), .CK(Clk), .RN(n106410), .Q(
        n109125), .QN(n102839) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][4]  ( .D(n104173), 
        .CK(Clk), .RN(n106410), .Q(n71967) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24591 ), .CK(Clk), .RN(n106410), .Q(
        n109126) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24527 ), .CK(Clk), .RN(n106410), .Q(
        n109127) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24495 ), .CK(Clk), .RN(n106410), .Q(
        n109128), .QN(n102269) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24463 ), .CK(Clk), .RN(n106410), .Q(n71972), .QN(n104641) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24431 ), .CK(Clk), .RN(n106410), .Q(
        n109129) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24399 ), .CK(Clk), .RN(n106410), .Q(
        n109130) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][4]  ( .D(n104194), 
        .CK(Clk), .RN(n106409), .Q(n109131) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24335 ), .CK(Clk), .RN(n106409), .Q(
        n109132) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24303 ), .CK(Clk), .RN(n106409), .Q(
        n109133) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24271 ), .CK(Clk), .RN(n106409), .Q(
        n109134), .QN(n102836) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24239 ), .CK(Clk), .RN(n106409), .Q(
        n109135) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24207 ), .CK(Clk), .RN(n106409), .Q(
        n109136) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24143 ), .CK(Clk), .RN(n106409), .Q(
        n109137) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][4]  ( .D(n104115), 
        .CK(Clk), .RN(n106409), .Q(n109138) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24047 ), .CK(Clk), .RN(n106409), .Q(
        n109139) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24015 ), .CK(Clk), .RN(n106409), .Q(n71986) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23983 ), .CK(Clk), .RN(n106408), .Q(
        n109140), .QN(n102267) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23951 ), .CK(Clk), .RN(n106408), .Q(
        n109141) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23919 ), .CK(Clk), .RN(n106408), .Q(
        n109142), .QN(n103438) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23887 ), .CK(Clk), .RN(n106408), .Q(
        n109143), .QN(n102834) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][4]  ( .D(n104122), 
        .CK(Clk), .RN(n106408), .Q(n109144) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23791 ), .CK(Clk), .RN(n106408), .Q(
        n109145) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23759 ), .CK(Clk), .RN(n106408), .Q(
        n109146), .QN(n101048) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23727 ), .CK(Clk), .RN(n106408), .Q(
        n109147) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23695 ), .CK(Clk), .RN(n106408), .Q(n71996) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23663 ), .CK(Clk), .RN(n106408), .Q(n71997), .QN(n104649) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23631 ), .CK(Clk), .RN(n106407), .Q(n71998) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23599 ), .CK(Clk), .RN(n106407), .Q(
        n109148) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23567 ), .CK(Clk), .RN(n106407), .Q(
        n109149) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23535 ), .CK(Clk), .RN(n106407), .Q(
        n109150), .QN(n103434) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23503 ), .CK(Clk), .RN(n106407), .Q(
        n109151) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23471 ), .CK(Clk), .RN(n106407), .Q(n72003) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23439 ), .CK(Clk), .RN(n106407), .Q(n72004) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23407 ), .CK(Clk), .RN(n106407), .Q(
        n109152) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23375 ), .CK(Clk), .RN(n106407), .Q(
        n109153) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23343 ), .CK(Clk), .RN(n106407), .Q(
        n109154) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23311 ), .CK(Clk), .RN(n106407), .Q(
        n109155) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23279 ), .CK(Clk), .RN(n106407), .Q(
        n109156) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23247 ), .CK(Clk), .RN(Rst), .Q(n109157), 
        .QN(n102832) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23215 ), .CK(Clk), .RN(Rst), .Q(n109158)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23183 ), .CK(Clk), .RN(Rst), .Q(n109159)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23151 ), .CK(Clk), .RN(Rst), .Q(n109160)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23119 ), .CK(Clk), .RN(Rst), .Q(n109161)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23087 ), .CK(Clk), .RN(Rst), .Q(n109162)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23055 ), .CK(Clk), .RN(Rst), .Q(n109163)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23023 ), .CK(Clk), .RN(Rst), .Q(n109164)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22991 ), .CK(Clk), .RN(Rst), .Q(n109165)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22959 ), .CK(Clk), .RN(Rst), .Q(n109166)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22927 ), .CK(Clk), .RN(Rst), .Q(n72020) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22895 ), .CK(Clk), .RN(Rst), .Q(n72021) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22863 ), .CK(Clk), .RN(Rst), .Q(n109167)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22831 ), .CK(Clk), .RN(Rst), .Q(n109168)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22799 ), .CK(Clk), .RN(Rst), .Q(n109169)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22767 ), .CK(Clk), .RN(Rst), .Q(n109170)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22735 ), .CK(Clk), .RN(Rst), .Q(n72026) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22703 ), .CK(Clk), .RN(Rst), .Q(n109171)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22671 ), .CK(Clk), .RN(Rst), .Q(n109172)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22639 ), .CK(Clk), .RN(Rst), .Q(n109173)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22607 ), .CK(Clk), .RN(Rst), .Q(n109174)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22575 ), .CK(Clk), .RN(Rst), .Q(n109175)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][4]  ( .D(
        \DLX_Datapath/RegisterFile/N22543 ), .CK(Clk), .RN(Rst), .Q(n72032), 
        .QN(n104516) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25871 ), .CK(Clk), .RN(Rst), .Q(n72033) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][4]  ( .D(n104257), 
        .CK(Clk), .RN(n106406), .Q(n109176) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25935 ), .CK(Clk), .RN(n106406), .Q(
        n109177) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25967 ), .CK(Clk), .RN(n106406), .Q(
        n109178), .QN(n103447) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25999 ), .CK(Clk), .RN(n106406), .Q(
        n109179) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26031 ), .CK(Clk), .RN(n106406), .Q(
        n109180) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26063 ), .CK(Clk), .RN(n106406), .Q(
        n109181) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26095 ), .CK(Clk), .RN(n106406), .Q(n72040) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26127 ), .CK(Clk), .RN(n106406), .Q(
        n109182), .QN(n101737) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26159 ), .CK(Clk), .RN(n106406), .Q(n72042) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26191 ), .CK(Clk), .RN(n106406), .Q(n72043) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26223 ), .CK(Clk), .RN(n106406), .Q(
        n109183) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26255 ), .CK(Clk), .RN(n106406), .Q(n72045) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26287 ), .CK(Clk), .RN(Rst), .Q(n109184)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26319 ), .CK(Clk), .RN(Rst), .Q(n109185)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26351 ), .CK(Clk), .RN(Rst), .Q(n109186)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26383 ), .CK(Clk), .RN(Rst), .Q(n109187)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26447 ), .CK(Clk), .RN(Rst), .Q(n109189)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26479 ), .CK(Clk), .RN(Rst), .Q(n109190), 
        .QN(n103449) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26511 ), .CK(Clk), .RN(Rst), .Q(n109191)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26543 ), .CK(Clk), .RN(Rst), .Q(n109192)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26575 ), .CK(Clk), .RN(Rst), .Q(n109193)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26607 ), .CK(Clk), .RN(Rst), .Q(n109194)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][4]  ( .D(n106963), 
        .CK(Clk), .RN(Rst), .Q(n109195) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26671 ), .CK(Clk), .RN(n106405), .Q(
        n109196), .QN(n102278) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26703 ), .CK(Clk), .RN(n106405), .Q(
        n109197), .QN(n102846) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26735 ), .CK(Clk), .RN(n106405), .Q(n72060), .QN(n104531) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][4]  ( .D(n106994), 
        .CK(Clk), .RN(n106405), .Q(n109198), .QN(n101738) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26831 ), .CK(Clk), .RN(n106405), .Q(
        n109200), .QN(n102847) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[4]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107066), .Q(
        \DLX_Datapath/next_A_IDEX[4] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[4]  ( .D(n106616), .CK(Clk), .RN(n106405), 
        .Q(n109201) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[4]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107032), .Q(
        \DLX_Datapath/next_B_IDEX [4]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[4]  ( .D(n106666), .CK(Clk), .RN(n106405), 
        .Q(n72065) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[4]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [4]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [4]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[4]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [4]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [4]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_shf_reg[4]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [4]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/B_shf [4]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[4]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N149 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [4]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[4]  ( .D(n103921), .GN(n106360), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [4]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[4]  ( .D(n104347), .CK(Clk), .RN(
        n106405), .Q(DataAddr[4]), .QN(n58618) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[4]  ( .D(n58928), .CK(Clk), .RN(n106405), 
        .Q(n109203) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[4]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [4]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[4]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [4]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [4]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[4]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [4]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [4]) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25840 ), .CK(Clk), .RN(n106405), .Q(n72073) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25808 ), .CK(Clk), .RN(n106408), .Q(
        n109206) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25776 ), .CK(Clk), .RN(n106413), .Q(
        n109207) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25744 ), .CK(Clk), .RN(n106425), .Q(
        n109208) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25680 ), .CK(Clk), .RN(n106488), .Q(
        n109209) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25616 ), .CK(Clk), .RN(n106488), .Q(
        n109210) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25584 ), .CK(Clk), .RN(n106488), .Q(
        n109211) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25552 ), .CK(Clk), .RN(n106488), .Q(
        n109212) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25520 ), .CK(Clk), .RN(n106488), .Q(
        n109213) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25488 ), .CK(Clk), .RN(Rst), .Q(n109214), 
        .QN(n100587) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25456 ), .CK(Clk), .RN(Rst), .Q(n72085) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25424 ), .CK(Clk), .RN(Rst), .Q(n109215)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25392 ), .CK(Clk), .RN(Rst), .Q(n109216)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25360 ), .CK(Clk), .RN(Rst), .Q(n109217)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25328 ), .CK(Clk), .RN(Rst), .Q(n109218)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25296 ), .CK(Clk), .RN(Rst), .Q(n109219), 
        .QN(n102863) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25264 ), .CK(Clk), .RN(Rst), .Q(n109220), 
        .QN(n102295) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25232 ), .CK(Clk), .RN(Rst), .Q(n109221), 
        .QN(n101751) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25200 ), .CK(Clk), .RN(Rst), .Q(n109222)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25168 ), .CK(Clk), .RN(Rst), .Q(n72094) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25136 ), .CK(Clk), .RN(Rst), .Q(n109223)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25072 ), .CK(Clk), .RN(Rst), .Q(n109224)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25040 ), .CK(Clk), .RN(Rst), .Q(n72098), 
        .QN(n104589) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25008 ), .CK(Clk), .RN(Rst), .Q(n109225)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24976 ), .CK(Clk), .RN(Rst), .Q(n109226), 
        .QN(n100619) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24944 ), .CK(Clk), .RN(Rst), .Q(n109227)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24912 ), .CK(Clk), .RN(Rst), .Q(n72102) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24880 ), .CK(Clk), .RN(Rst), .Q(n109228), 
        .QN(n101174) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24848 ), .CK(Clk), .RN(Rst), .Q(n109229)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24816 ), .CK(Clk), .RN(Rst), .Q(n109230)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24784 ), .CK(Clk), .RN(Rst), .Q(n72106) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24752 ), .CK(Clk), .RN(Rst), .Q(n109231)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24688 ), .CK(Clk), .RN(n106420), .Q(
        n109232) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24656 ), .CK(Clk), .RN(Rst), .Q(n109233), 
        .QN(n102859) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24624 ), .CK(Clk), .RN(Rst), .Q(n72111) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24592 ), .CK(Clk), .RN(Rst), .Q(n109234)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24528 ), .CK(Clk), .RN(Rst), .Q(n109235)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24496 ), .CK(Clk), .RN(Rst), .Q(n109236), 
        .QN(n102288) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24464 ), .CK(Clk), .RN(n106480), .Q(n72116), .QN(n104642) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24432 ), .CK(Clk), .RN(n106491), .Q(
        n109237) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24400 ), .CK(Clk), .RN(n106481), .Q(
        n109238) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24368 ), .CK(Clk), .RN(Rst), .Q(n109239)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24336 ), .CK(Clk), .RN(n106400), .Q(
        n109240) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24304 ), .CK(Clk), .RN(n106435), .Q(
        n109241) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24272 ), .CK(Clk), .RN(Rst), .Q(n109242), 
        .QN(n102856) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24240 ), .CK(Clk), .RN(n106454), .Q(
        n109243) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24208 ), .CK(Clk), .RN(n106453), .Q(
        n109244) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24144 ), .CK(Clk), .RN(Rst), .Q(n109245)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][5]  ( .D(n104120), 
        .CK(Clk), .RN(n106442), .Q(n109246) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24048 ), .CK(Clk), .RN(n106459), .Q(
        n109247) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24016 ), .CK(Clk), .RN(n106452), .Q(n72130) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23984 ), .CK(Clk), .RN(Rst), .Q(n109248), 
        .QN(n102286) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23952 ), .CK(Clk), .RN(n106487), .Q(
        n109249) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23920 ), .CK(Clk), .RN(n106487), .Q(
        n109250), .QN(n103458) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23888 ), .CK(Clk), .RN(n106487), .Q(
        n109251), .QN(n102854) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23856 ), .CK(Clk), .RN(n106487), .Q(
        n109252) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23792 ), .CK(Clk), .RN(n106487), .Q(
        n109253) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23760 ), .CK(Clk), .RN(n106487), .Q(
        n109254), .QN(n101047) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23728 ), .CK(Clk), .RN(n106487), .Q(
        n109255) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23696 ), .CK(Clk), .RN(n106487), .Q(n72140) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23664 ), .CK(Clk), .RN(n106487), .Q(
        n109256), .QN(n101016) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23632 ), .CK(Clk), .RN(n106487), .Q(n72142) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23600 ), .CK(Clk), .RN(n106487), .Q(
        n109257) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23568 ), .CK(Clk), .RN(Rst), .Q(n109258)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23536 ), .CK(Clk), .RN(n106410), .Q(
        n109259), .QN(n103454) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23504 ), .CK(Clk), .RN(Rst), .Q(n109260)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23472 ), .CK(Clk), .RN(Rst), .Q(n72147) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23440 ), .CK(Clk), .RN(Rst), .Q(n72148) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23408 ), .CK(Clk), .RN(Rst), .Q(n109261)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23376 ), .CK(Clk), .RN(n106479), .Q(
        n109262) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23344 ), .CK(Clk), .RN(Rst), .Q(n109263)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23312 ), .CK(Clk), .RN(Rst), .Q(n109264)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23280 ), .CK(Clk), .RN(n106382), .Q(
        n109265) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23248 ), .CK(Clk), .RN(n106489), .Q(
        n109266), .QN(n102852) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23216 ), .CK(Clk), .RN(Rst), .Q(n109267)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23184 ), .CK(Clk), .RN(n106460), .Q(
        n109268) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23152 ), .CK(Clk), .RN(n106429), .Q(
        n109269) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23120 ), .CK(Clk), .RN(n106485), .Q(
        n109270) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23088 ), .CK(Clk), .RN(n106482), .Q(
        n109271) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23056 ), .CK(Clk), .RN(n106401), .Q(
        n109272) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23024 ), .CK(Clk), .RN(n106483), .Q(
        n109273) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22992 ), .CK(Clk), .RN(n106398), .Q(
        n109274) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22960 ), .CK(Clk), .RN(n106443), .Q(
        n109275) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22928 ), .CK(Clk), .RN(n106465), .Q(n72164) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22896 ), .CK(Clk), .RN(n106486), .Q(n72165) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22864 ), .CK(Clk), .RN(n106466), .Q(
        n109276) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22832 ), .CK(Clk), .RN(n106473), .Q(
        n109277) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22800 ), .CK(Clk), .RN(Rst), .Q(n109278)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22768 ), .CK(Clk), .RN(Rst), .Q(n109279)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22736 ), .CK(Clk), .RN(n106373), .Q(n72170) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22672 ), .CK(Clk), .RN(n106472), .Q(
        n109280) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22640 ), .CK(Clk), .RN(n106475), .Q(
        n109281) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22608 ), .CK(Clk), .RN(n106471), .Q(
        n109282) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22576 ), .CK(Clk), .RN(n106470), .Q(
        n109283) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22544 ), .CK(Clk), .RN(Rst), .Q(n72176), 
        .QN(n104517) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][5]  ( .D(n104258), 
        .CK(Clk), .RN(n106457), .Q(n109284) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25936 ), .CK(Clk), .RN(Rst), .Q(n109285)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25968 ), .CK(Clk), .RN(Rst), .Q(n109286), 
        .QN(n103467) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26000 ), .CK(Clk), .RN(Rst), .Q(n109287)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][5]  ( .D(n104236), 
        .CK(Clk), .RN(n106481), .Q(n109288) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26064 ), .CK(Clk), .RN(Rst), .Q(n109289)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26096 ), .CK(Clk), .RN(Rst), .Q(n72184) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26128 ), .CK(Clk), .RN(Rst), .Q(n109290), 
        .QN(n101755) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26160 ), .CK(Clk), .RN(Rst), .Q(n72186) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26192 ), .CK(Clk), .RN(Rst), .Q(n72187) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26224 ), .CK(Clk), .RN(Rst), .Q(n109291)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26256 ), .CK(Clk), .RN(n106480), .Q(n72189) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26288 ), .CK(Clk), .RN(n106491), .Q(
        n109292) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26320 ), .CK(Clk), .RN(n106427), .Q(
        n109293) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26352 ), .CK(Clk), .RN(Rst), .Q(n109294)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26384 ), .CK(Clk), .RN(Rst), .Q(n109295)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26448 ), .CK(Clk), .RN(Rst), .Q(n109297)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26480 ), .CK(Clk), .RN(n106372), .Q(
        n109298), .QN(n103469) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26512 ), .CK(Clk), .RN(Rst), .Q(n109299)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26544 ), .CK(Clk), .RN(Rst), .Q(n109300)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26576 ), .CK(Clk), .RN(n106508), .Q(
        n109301) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26608 ), .CK(Clk), .RN(Rst), .Q(n109302)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][5]  ( .D(n106964), 
        .CK(Clk), .RN(Rst), .Q(n109303) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26672 ), .CK(Clk), .RN(Rst), .Q(n109304), 
        .QN(n102297) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26704 ), .CK(Clk), .RN(Rst), .Q(n109305), 
        .QN(n102866) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26736 ), .CK(Clk), .RN(n106409), .Q(n72204), .QN(n104532) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][5]  ( .D(n106995), 
        .CK(Clk), .RN(Rst), .Q(n109306), .QN(n101756) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26832 ), .CK(Clk), .RN(Rst), .Q(n109308), 
        .QN(n102867) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[5]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107067), .Q(
        \DLX_Datapath/next_A_IDEX[5] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[5]  ( .D(n106602), .CK(Clk), .RN(n106395), 
        .Q(n109309) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[5]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107033), .Q(
        \DLX_Datapath/next_B_IDEX [5]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[5]  ( .D(n106676), .CK(Clk), .RN(Rst), .Q(
        n72209) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[5]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [5]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [5]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[4]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N117 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [4]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[5]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [5]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [5]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[5]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N150 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [5]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[5]  ( .D(n106887), .GN(n106360), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [5]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[5]  ( .D(n104348), .CK(Clk), .RN(Rst), 
        .Q(DataAddr[5]), .QN(n58614) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[5]  ( .D(n58924), .CK(Clk), .RN(Rst), .Q(
        n109312) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[5]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [5]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[5]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [5]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [5]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[5]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [5]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [5]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[5]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N118 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [5]) );
  DFFR_X2 \DLX_Datapath/PC_reg[5]  ( .D(n60320), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [1]), .QN(n62201) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[4]  ( .D(n103949), .CK(Clk), .RN(Rst), .Q(
        n109316) );
  DFFR_X2 \DLX_Datapath/PC_reg[4]  ( .D(n60321), .CK(Clk), .RN(n106419), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [0]), .QN(net2465400)
         );
  DFFR_X2 \DLX_Datapath/PC_IFID_reg[4]  ( .D(n60225), .CK(Clk), .RN(n106392), 
        .Q(n109317), .QN(n59423) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[9][0]  ( .D(n60180), .CK(
        Clk), .RN(n106458), .Q(n109318) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[1][0]  ( .D(n60164), .CK(
        Clk), .RN(Rst), .Q(n109319) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[17][0]  ( .D(n60196), 
        .CK(Clk), .RN(n106393), .Q(n109320) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[5]  ( .D(n103933), .CK(Clk), .RN(n106409), 
        .Q(n109321) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[6]  ( .D(n103934), .CK(Clk), .RN(n106406), 
        .Q(n109322) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[7]  ( .D(n103935), .CK(Clk), .RN(n106427), 
        .Q(n109323) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25841 ), .CK(Clk), .RN(Rst), .Q(n72224) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25809 ), .CK(Clk), .RN(n106405), .Q(
        n109324) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25777 ), .CK(Clk), .RN(n106404), .Q(
        n109325) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25745 ), .CK(Clk), .RN(n106403), .Q(
        n109326) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25681 ), .CK(Clk), .RN(n106402), .Q(
        n109327) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25617 ), .CK(Clk), .RN(n106438), .Q(
        n109328) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25585 ), .CK(Clk), .RN(n106437), .Q(
        n109329) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25553 ), .CK(Clk), .RN(n106484), .Q(
        n109330) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25521 ), .CK(Clk), .RN(Rst), .Q(n109331)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25489 ), .CK(Clk), .RN(Rst), .Q(n109332), 
        .QN(n100586) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25457 ), .CK(Clk), .RN(Rst), .Q(n72236) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25425 ), .CK(Clk), .RN(Rst), .Q(n109333)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25393 ), .CK(Clk), .RN(Rst), .Q(n109334)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25361 ), .CK(Clk), .RN(n106476), .Q(
        n109335) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][6]  ( .D(n104300), 
        .CK(Clk), .RN(n106414), .Q(n109336) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25297 ), .CK(Clk), .RN(n106417), .Q(
        n109337), .QN(n102883) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25265 ), .CK(Clk), .RN(Rst), .Q(n109338), 
        .QN(n102315) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25233 ), .CK(Clk), .RN(Rst), .Q(n109339), 
        .QN(n101769) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25201 ), .CK(Clk), .RN(n106416), .Q(
        n109340) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25169 ), .CK(Clk), .RN(n106477), .Q(n72245) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25137 ), .CK(Clk), .RN(n106428), .Q(
        n109341) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][6]  ( .D(n104284), 
        .CK(Clk), .RN(n106415), .Q(n109342) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25041 ), .CK(Clk), .RN(n106402), .Q(n72249), .QN(n104590) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25009 ), .CK(Clk), .RN(Rst), .Q(n109343)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24977 ), .CK(Clk), .RN(n106433), .Q(
        n109344), .QN(n100618) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][6]  ( .D(n104290), 
        .CK(Clk), .RN(n106437), .Q(n109345) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24913 ), .CK(Clk), .RN(n106432), .Q(n72253) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24881 ), .CK(Clk), .RN(n106485), .Q(
        n109346), .QN(n101173) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24849 ), .CK(Clk), .RN(Rst), .Q(n109347)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][6]  ( .D(n104152), 
        .CK(Clk), .RN(n106438), .Q(n109348) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24785 ), .CK(Clk), .RN(Rst), .Q(n72257) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24753 ), .CK(Clk), .RN(n106439), .Q(
        n109349) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24689 ), .CK(Clk), .RN(Rst), .Q(n109350)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24657 ), .CK(Clk), .RN(Rst), .Q(n109351), 
        .QN(n102879) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24625 ), .CK(Clk), .RN(Rst), .Q(n72262) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24593 ), .CK(Clk), .RN(Rst), .Q(n109352)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24529 ), .CK(Clk), .RN(Rst), .Q(n109353)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24497 ), .CK(Clk), .RN(Rst), .Q(n109354), 
        .QN(n102308) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24465 ), .CK(Clk), .RN(Rst), .Q(n72267), 
        .QN(n104643) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][6]  ( .D(n104147), 
        .CK(Clk), .RN(Rst), .Q(n109355) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24401 ), .CK(Clk), .RN(Rst), .Q(n109356)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][6]  ( .D(n104195), 
        .CK(Clk), .RN(Rst), .Q(n109357) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24337 ), .CK(Clk), .RN(Rst), .Q(n109358)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][6]  ( .D(n104110), 
        .CK(Clk), .RN(Rst), .Q(n109359) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24273 ), .CK(Clk), .RN(Rst), .Q(n109360), 
        .QN(n102876) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24241 ), .CK(Clk), .RN(Rst), .Q(n109361)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24209 ), .CK(Clk), .RN(Rst), .Q(n109362)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24145 ), .CK(Clk), .RN(n106495), .Q(
        n109363) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][6]  ( .D(n104116), 
        .CK(Clk), .RN(Rst), .Q(n109364) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][6]  ( .D(n104075), 
        .CK(Clk), .RN(n106444), .Q(n109365) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24017 ), .CK(Clk), .RN(Rst), .Q(n72281) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23985 ), .CK(Clk), .RN(Rst), .Q(n109366), 
        .QN(n102306) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23953 ), .CK(Clk), .RN(Rst), .Q(n109367)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][6]  ( .D(n104086), 
        .CK(Clk), .RN(Rst), .Q(n109368), .QN(n103477) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23889 ), .CK(Clk), .RN(n106371), .Q(
        n109369), .QN(n102874) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][6]  ( .D(n104124), 
        .CK(Clk), .RN(Rst), .Q(n109370) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23793 ), .CK(Clk), .RN(Rst), .Q(n109371)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23761 ), .CK(Clk), .RN(Rst), .Q(n109372), 
        .QN(n101046) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23729 ), .CK(Clk), .RN(Rst), .Q(n109373)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23697 ), .CK(Clk), .RN(Rst), .Q(n72291) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23665 ), .CK(Clk), .RN(Rst), .Q(n109374), 
        .QN(n101015) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23633 ), .CK(Clk), .RN(Rst), .Q(n72293) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23601 ), .CK(Clk), .RN(Rst), .Q(n109375)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23569 ), .CK(Clk), .RN(Rst), .Q(n109376)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][6]  ( .D(n104026), 
        .CK(Clk), .RN(Rst), .Q(n109377), .QN(n103473) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23505 ), .CK(Clk), .RN(Rst), .Q(n109378)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23473 ), .CK(Clk), .RN(Rst), .Q(n72298) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23441 ), .CK(Clk), .RN(Rst), .Q(n72299) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23409 ), .CK(Clk), .RN(Rst), .Q(n109379)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23377 ), .CK(Clk), .RN(Rst), .Q(n109380)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][6]  ( .D(n104060), 
        .CK(Clk), .RN(Rst), .Q(n109381) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23313 ), .CK(Clk), .RN(Rst), .Q(n109382)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][6]  ( .D(n103999), 
        .CK(Clk), .RN(Rst), .Q(n109383) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23249 ), .CK(Clk), .RN(Rst), .Q(n109384), 
        .QN(n102872) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23217 ), .CK(Clk), .RN(Rst), .Q(n109385)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23185 ), .CK(Clk), .RN(Rst), .Q(n109386)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23153 ), .CK(Clk), .RN(Rst), .Q(n109387)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23121 ), .CK(Clk), .RN(Rst), .Q(n109388)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23089 ), .CK(Clk), .RN(Rst), .Q(n109389)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23057 ), .CK(Clk), .RN(Rst), .Q(n109390)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][6]  ( .D(n103991), 
        .CK(Clk), .RN(Rst), .Q(n109391) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22993 ), .CK(Clk), .RN(Rst), .Q(n109392)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22961 ), .CK(Clk), .RN(Rst), .Q(n109393)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22929 ), .CK(Clk), .RN(Rst), .Q(n72315) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][6]  ( .D(n103994), 
        .CK(Clk), .RN(Rst), .Q(n72316) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22865 ), .CK(Clk), .RN(Rst), .Q(n109394)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22833 ), .CK(Clk), .RN(Rst), .Q(n109395)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22801 ), .CK(Clk), .RN(Rst), .Q(n109396)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22769 ), .CK(Clk), .RN(Rst), .Q(n109397)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22737 ), .CK(Clk), .RN(Rst), .Q(n72321) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22705 ), .CK(Clk), .RN(n106491), .Q(
        n109398) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22673 ), .CK(Clk), .RN(n106491), .Q(
        n109399) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22641 ), .CK(Clk), .RN(n106491), .Q(
        n109400) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22609 ), .CK(Clk), .RN(n106491), .Q(
        n109401) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22577 ), .CK(Clk), .RN(n106491), .Q(
        n109402) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][6]  ( .D(
        \DLX_Datapath/RegisterFile/N22545 ), .CK(Clk), .RN(n106491), .Q(n72327), .QN(n104518) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25873 ), .CK(Clk), .RN(n106491), .Q(n72328) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][6]  ( .D(n104260), 
        .CK(Clk), .RN(n106491), .Q(n109403) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25937 ), .CK(Clk), .RN(n106491), .Q(
        n109404) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][6]  ( .D(n104317), 
        .CK(Clk), .RN(n106491), .Q(n109405), .QN(n103486) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26001 ), .CK(Clk), .RN(n106491), .Q(
        n109406) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26033 ), .CK(Clk), .RN(n106491), .Q(
        n109407) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26065 ), .CK(Clk), .RN(Rst), .Q(n109408)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26097 ), .CK(Clk), .RN(n106440), .Q(n72335) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26129 ), .CK(Clk), .RN(n106442), .Q(
        n109409), .QN(n101771) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26161 ), .CK(Clk), .RN(n106441), .Q(n72337) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26193 ), .CK(Clk), .RN(n106484), .Q(n72338) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26225 ), .CK(Clk), .RN(n106443), .Q(
        n109410) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26257 ), .CK(Clk), .RN(n106486), .Q(n72340) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26289 ), .CK(Clk), .RN(n106429), .Q(
        n109411) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26321 ), .CK(Clk), .RN(n106482), .Q(
        n109412) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26353 ), .CK(Clk), .RN(n106483), .Q(
        n109413) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26385 ), .CK(Clk), .RN(n106485), .Q(
        n109414) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26449 ), .CK(Clk), .RN(Rst), .Q(n109416)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26481 ), .CK(Clk), .RN(Rst), .Q(n109417), 
        .QN(n103488) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26513 ), .CK(Clk), .RN(Rst), .Q(n109418)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26545 ), .CK(Clk), .RN(Rst), .Q(n109419)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26577 ), .CK(Clk), .RN(Rst), .Q(n109420)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26609 ), .CK(Clk), .RN(Rst), .Q(n109421)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][6]  ( .D(n106965), 
        .CK(Clk), .RN(Rst), .Q(n109422) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26673 ), .CK(Clk), .RN(Rst), .Q(n109423), 
        .QN(n102317) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26705 ), .CK(Clk), .RN(Rst), .Q(n109424), 
        .QN(n102886) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][6]  ( .D(n104321), 
        .CK(Clk), .RN(Rst), .Q(n72355), .QN(n104526) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][6]  ( .D(n106996), 
        .CK(Clk), .RN(Rst), .Q(n109425), .QN(n101772) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26833 ), .CK(Clk), .RN(n106490), .Q(
        n109427), .QN(n102887) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[6]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107068), .Q(
        \DLX_Datapath/next_A_IDEX[6] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[6]  ( .D(n106617), .CK(Clk), .RN(n106490), 
        .Q(n109428) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[6]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [6]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[6]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [6]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [6]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[6]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [6]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [6]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[6]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107034), .Q(
        \DLX_Datapath/next_B_IDEX [6]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[6]  ( .D(n106667), .CK(Clk), .RN(n106490), 
        .Q(n72362) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[6]  ( .D(n58922), .CK(Clk), .RN(n106490), 
        .Q(n109431) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[6]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [6]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [6]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[6]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N119 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [6]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[6]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(\DLX_Datapath/MUX_HDU_ALUInB [6]), .Q(\DLX_Datapath/ArithLogUnit/B_log [6]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[6]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N151 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [6]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[6]  ( .D(n107613), .GN(n60159), 
        .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [6]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[7]  ( .D(n107614), .GN(n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [7]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[8]  ( .D(n104361), .GN(n60159), 
        .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [8]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[9]  ( .D(n106893), .GN(n106360), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [9]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[9]  ( .D(n104349), .CK(Clk), .RN(
        n106490), .Q(DataAddr[9]), .QN(n58609) );
  DFFR_X2 \DLX_Datapath/PC_reg[9]  ( .D(n60316), .CK(Clk), .RN(n106490), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [1]), .QN(n104502) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[8]  ( .D(n106541), .CK(Clk), .RN(n106490), 
        .Q(n109435) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[8]  ( .D(n106634), .CK(Clk), .RN(n106490), 
        .Q(n72370) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[8]  ( .D(n58919), .CK(Clk), .RN(n106490), 
        .Q(n109436), .QN(n59331) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[9]  ( .D(n106540), .CK(Clk), .RN(n106490), 
        .Q(n109437) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[9]  ( .D(n106655), .CK(Clk), .RN(n106490), 
        .Q(n72372) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[9]  ( .D(n58918), .CK(Clk), .RN(n106490), 
        .Q(n109438), .QN(n59332) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25843 ), .CK(Clk), .RN(n106489), .Q(n72375) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25811 ), .CK(Clk), .RN(n106489), .Q(
        n109439) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25779 ), .CK(Clk), .RN(n106489), .Q(
        n109440) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25747 ), .CK(Clk), .RN(n106489), .Q(
        n109441) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25683 ), .CK(Clk), .RN(n106489), .Q(
        n109442) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25619 ), .CK(Clk), .RN(n106489), .Q(
        n109443) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25587 ), .CK(Clk), .RN(n106489), .Q(
        n109444) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25555 ), .CK(Clk), .RN(n106489), .Q(
        n109445) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25523 ), .CK(Clk), .RN(n106489), .Q(
        n109446) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25491 ), .CK(Clk), .RN(n106488), .Q(
        n109447), .QN(n100584) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25459 ), .CK(Clk), .RN(n106488), .Q(n72387) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25427 ), .CK(Clk), .RN(n106488), .Q(
        n109448) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25395 ), .CK(Clk), .RN(n106488), .Q(
        n109449) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25363 ), .CK(Clk), .RN(n106488), .Q(
        n109450) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][8]  ( .D(n104303), 
        .CK(Clk), .RN(n106488), .Q(n109451) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25299 ), .CK(Clk), .RN(Rst), .Q(n109452), 
        .QN(n102923) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25267 ), .CK(Clk), .RN(Rst), .Q(n109453), 
        .QN(n102355) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25235 ), .CK(Clk), .RN(Rst), .Q(n109454), 
        .QN(n101803) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25203 ), .CK(Clk), .RN(Rst), .Q(n109455)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25171 ), .CK(Clk), .RN(Rst), .Q(n72396) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25139 ), .CK(Clk), .RN(n106507), .Q(
        n109456) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][8]  ( .D(n104285), 
        .CK(Clk), .RN(Rst), .Q(n109457) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25043 ), .CK(Clk), .RN(Rst), .Q(n72400), 
        .QN(n104592) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25011 ), .CK(Clk), .RN(Rst), .Q(n109458)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24979 ), .CK(Clk), .RN(Rst), .Q(n109459), 
        .QN(n100616) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][8]  ( .D(n104291), 
        .CK(Clk), .RN(Rst), .Q(n109460) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24915 ), .CK(Clk), .RN(Rst), .Q(n72404) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24883 ), .CK(Clk), .RN(Rst), .Q(n109461), 
        .QN(n101171) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24851 ), .CK(Clk), .RN(Rst), .Q(n109462)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24819 ), .CK(Clk), .RN(Rst), .Q(n109463)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24787 ), .CK(Clk), .RN(Rst), .Q(n72408) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][8]  ( .D(n104180), 
        .CK(Clk), .RN(Rst), .Q(n109464) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][8]  ( .D(n104159), 
        .CK(Clk), .RN(Rst), .Q(n109465) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24659 ), .CK(Clk), .RN(n106482), .Q(
        n109466), .QN(n102919) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][8]  ( .D(n104177), 
        .CK(Clk), .RN(n106482), .Q(n72413) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24595 ), .CK(Clk), .RN(n106482), .Q(
        n109467) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24531 ), .CK(Clk), .RN(n106482), .Q(
        n109468) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24499 ), .CK(Clk), .RN(n106482), .Q(
        n109469), .QN(n102348) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24467 ), .CK(Clk), .RN(n106482), .Q(n72418), .QN(n104645) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24435 ), .CK(Clk), .RN(n106482), .Q(
        n109470) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24403 ), .CK(Clk), .RN(n106482), .Q(
        n109471) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24371 ), .CK(Clk), .RN(n106482), .Q(
        n109472) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24339 ), .CK(Clk), .RN(n106482), .Q(
        n109473) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24307 ), .CK(Clk), .RN(n106482), .Q(
        n109474) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24275 ), .CK(Clk), .RN(Rst), .Q(n109475), 
        .QN(n102916) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24243 ), .CK(Clk), .RN(Rst), .Q(n109476)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24211 ), .CK(Clk), .RN(Rst), .Q(n109477)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24147 ), .CK(Clk), .RN(Rst), .Q(n109478)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24115 ), .CK(Clk), .RN(Rst), .Q(n109479)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24051 ), .CK(Clk), .RN(Rst), .Q(n109480)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24019 ), .CK(Clk), .RN(Rst), .Q(n72432) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23987 ), .CK(Clk), .RN(Rst), .Q(n109481), 
        .QN(n102346) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23955 ), .CK(Clk), .RN(Rst), .Q(n109482)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23923 ), .CK(Clk), .RN(Rst), .Q(n109483), 
        .QN(n103515) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23891 ), .CK(Clk), .RN(n106481), .Q(
        n109484), .QN(n102914) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23859 ), .CK(Clk), .RN(n106481), .Q(
        n109485) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23795 ), .CK(Clk), .RN(n106481), .Q(
        n109486) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23763 ), .CK(Clk), .RN(n106481), .Q(
        n109487), .QN(n101044) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23731 ), .CK(Clk), .RN(n106481), .Q(
        n109488) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23699 ), .CK(Clk), .RN(n106481), .Q(n72442) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23667 ), .CK(Clk), .RN(n106481), .Q(
        n109489), .QN(n101013) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23635 ), .CK(Clk), .RN(n106481), .Q(n72444) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23603 ), .CK(Clk), .RN(n106481), .Q(
        n109490) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23571 ), .CK(Clk), .RN(n106481), .Q(
        n109491) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23539 ), .CK(Clk), .RN(n106481), .Q(
        n109492), .QN(n103511) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23507 ), .CK(Clk), .RN(Rst), .Q(n109493)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][8]  ( .D(n104047), 
        .CK(Clk), .RN(Rst), .Q(n72449) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23443 ), .CK(Clk), .RN(Rst), .Q(n72450) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23411 ), .CK(Clk), .RN(Rst), .Q(n109494)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23379 ), .CK(Clk), .RN(Rst), .Q(n109495)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23347 ), .CK(Clk), .RN(Rst), .Q(n109496)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23315 ), .CK(Clk), .RN(Rst), .Q(n109497)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23283 ), .CK(Clk), .RN(Rst), .Q(n109498)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23251 ), .CK(Clk), .RN(Rst), .Q(n109499), 
        .QN(n102912) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23219 ), .CK(Clk), .RN(Rst), .Q(n109500)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23187 ), .CK(Clk), .RN(Rst), .Q(n109501)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23155 ), .CK(Clk), .RN(Rst), .Q(n109502)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23123 ), .CK(Clk), .RN(Rst), .Q(n109503)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23091 ), .CK(Clk), .RN(Rst), .Q(n109504)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23059 ), .CK(Clk), .RN(Rst), .Q(n109505)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23027 ), .CK(Clk), .RN(Rst), .Q(n109506)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22995 ), .CK(Clk), .RN(Rst), .Q(n109507)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22963 ), .CK(Clk), .RN(Rst), .Q(n109508)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22931 ), .CK(Clk), .RN(Rst), .Q(n72466) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22899 ), .CK(Clk), .RN(Rst), .Q(n72467) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22867 ), .CK(Clk), .RN(Rst), .Q(n109509)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22835 ), .CK(Clk), .RN(Rst), .Q(n109510)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22803 ), .CK(Clk), .RN(Rst), .Q(n109511)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22771 ), .CK(Clk), .RN(Rst), .Q(n109512)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22739 ), .CK(Clk), .RN(Rst), .Q(n72472) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22707 ), .CK(Clk), .RN(Rst), .Q(n109513)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22675 ), .CK(Clk), .RN(Rst), .Q(n109514)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22643 ), .CK(Clk), .RN(Rst), .Q(n109515)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22611 ), .CK(Clk), .RN(Rst), .Q(n109516)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22579 ), .CK(Clk), .RN(Rst), .Q(n109517)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][8]  ( .D(
        \DLX_Datapath/RegisterFile/N22547 ), .CK(Clk), .RN(Rst), .Q(n72478), 
        .QN(n104519) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25875 ), .CK(Clk), .RN(Rst), .Q(n72479) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][8]  ( .D(n104273), 
        .CK(Clk), .RN(Rst), .Q(n109518) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25939 ), .CK(Clk), .RN(Rst), .Q(n109519)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25971 ), .CK(Clk), .RN(Rst), .Q(n109520), 
        .QN(n103524) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26003 ), .CK(Clk), .RN(n106480), .Q(
        n109521) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][8]  ( .D(n104226), 
        .CK(Clk), .RN(n106480), .Q(n109522) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26067 ), .CK(Clk), .RN(n106480), .Q(
        n109523) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26099 ), .CK(Clk), .RN(n106480), .Q(n72486) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26131 ), .CK(Clk), .RN(n106480), .Q(
        n109524), .QN(n101805) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26163 ), .CK(Clk), .RN(n106480), .Q(n72488) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26195 ), .CK(Clk), .RN(n106480), .Q(n72489) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26227 ), .CK(Clk), .RN(n106480), .Q(
        n109525) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26259 ), .CK(Clk), .RN(n106480), .Q(n72491) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26291 ), .CK(Clk), .RN(n106480), .Q(
        n109526) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26323 ), .CK(Clk), .RN(n106480), .Q(
        n109527) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26355 ), .CK(Clk), .RN(n106480), .Q(
        n109528) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26387 ), .CK(Clk), .RN(Rst), .Q(n109529)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26451 ), .CK(Clk), .RN(Rst), .Q(n109531)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26483 ), .CK(Clk), .RN(Rst), .Q(n109532), 
        .QN(n103526) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26515 ), .CK(Clk), .RN(Rst), .Q(n109533)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26547 ), .CK(Clk), .RN(Rst), .Q(n109534)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26579 ), .CK(Clk), .RN(Rst), .Q(n109535)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26611 ), .CK(Clk), .RN(Rst), .Q(n109536)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][8]  ( .D(n106967), 
        .CK(Clk), .RN(Rst), .Q(n109537) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26675 ), .CK(Clk), .RN(Rst), .Q(n109538), 
        .QN(n102357) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26707 ), .CK(Clk), .RN(Rst), .Q(n109539), 
        .QN(n102926) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26739 ), .CK(Clk), .RN(Rst), .Q(n72506), 
        .QN(n104534) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][8]  ( .D(n106998), 
        .CK(Clk), .RN(n106479), .Q(n109540), .QN(n101806) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26835 ), .CK(Clk), .RN(n106479), .Q(
        n109542), .QN(n102927) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[8]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107070), .Q(
        \DLX_Datapath/next_A_IDEX[8] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[8]  ( .D(n106618), .CK(Clk), .RN(n106479), 
        .Q(n109543) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[8]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107036), .Q(
        \DLX_Datapath/next_B_IDEX [8]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[8]  ( .D(n106668), .CK(Clk), .RN(n106479), 
        .Q(n72511) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[8]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [8]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [8]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[8]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [8]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [8]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[8]  ( .D(n103920), .GN(n60158), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [8]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[8]  ( .D(n104350), .CK(Clk), .RN(
        n106479), .Q(DataAddr[8]), .QN(n58604) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[8]  ( .D(n58914), .CK(Clk), .RN(n106479), 
        .Q(n109544) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[8]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [8]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[8]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [8]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [8]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[8]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [8]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [8]) );
  DFFR_X2 \DLX_Datapath/PC_reg[8]  ( .D(n60317), .CK(Clk), .RN(n106479), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [0]), .QN(n62202) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[8]  ( .D(n103945), .CK(Clk), .RN(n106479), 
        .Q(n109547) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[9]  ( .D(n103950), .CK(Clk), .RN(n106479), 
        .Q(n109548) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[10]  ( .D(n103936), .CK(Clk), .RN(n106479), 
        .Q(n109549) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25846 ), .CK(Clk), .RN(Rst), .Q(n72523) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25814 ), .CK(Clk), .RN(Rst), .Q(n109550)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25782 ), .CK(Clk), .RN(Rst), .Q(n109551)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25750 ), .CK(Clk), .RN(Rst), .Q(n109552)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25686 ), .CK(Clk), .RN(Rst), .Q(n109553)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25622 ), .CK(Clk), .RN(Rst), .Q(n109554)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25590 ), .CK(Clk), .RN(Rst), .Q(n109555)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25558 ), .CK(Clk), .RN(Rst), .Q(n109556)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25526 ), .CK(Clk), .RN(Rst), .Q(n109557)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25494 ), .CK(Clk), .RN(Rst), .Q(n109558), 
        .QN(n100581) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25462 ), .CK(Clk), .RN(n106431), .Q(n72535) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25430 ), .CK(Clk), .RN(Rst), .Q(n109559)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25398 ), .CK(Clk), .RN(Rst), .Q(n109560)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25366 ), .CK(Clk), .RN(Rst), .Q(n109561)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25334 ), .CK(Clk), .RN(Rst), .Q(n109562)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25302 ), .CK(Clk), .RN(Rst), .Q(n109563), 
        .QN(n102980) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25270 ), .CK(Clk), .RN(Rst), .Q(n109564), 
        .QN(n102413) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25238 ), .CK(Clk), .RN(Rst), .Q(n109565), 
        .QN(n101855) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25206 ), .CK(Clk), .RN(Rst), .Q(n109566)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25174 ), .CK(Clk), .RN(n106463), .Q(n72544) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25142 ), .CK(Clk), .RN(n106462), .Q(
        n109567) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25078 ), .CK(Clk), .RN(n106429), .Q(
        n109568) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25046 ), .CK(Clk), .RN(n106485), .Q(n72548), .QN(n104595) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25014 ), .CK(Clk), .RN(n106479), .Q(
        n109569) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24982 ), .CK(Clk), .RN(n106489), .Q(
        n109570), .QN(n100613) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24950 ), .CK(Clk), .RN(Rst), .Q(n109571)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24918 ), .CK(Clk), .RN(n106433), .Q(n72552) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24886 ), .CK(Clk), .RN(n106432), .Q(
        n109572), .QN(n101168) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24854 ), .CK(Clk), .RN(n106460), .Q(
        n109573) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24822 ), .CK(Clk), .RN(Rst), .Q(n109574)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24790 ), .CK(Clk), .RN(Rst), .Q(n72556) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24758 ), .CK(Clk), .RN(Rst), .Q(n109575)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24694 ), .CK(Clk), .RN(Rst), .Q(n109576)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24662 ), .CK(Clk), .RN(Rst), .Q(n109577), 
        .QN(n101150) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24630 ), .CK(Clk), .RN(Rst), .Q(n72561) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24598 ), .CK(Clk), .RN(Rst), .Q(n109578)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24534 ), .CK(Clk), .RN(Rst), .Q(n109579)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24502 ), .CK(Clk), .RN(Rst), .Q(n109580), 
        .QN(n102406) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24470 ), .CK(Clk), .RN(Rst), .Q(n72566), 
        .QN(n104616) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24438 ), .CK(Clk), .RN(Rst), .Q(n109581)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24406 ), .CK(Clk), .RN(n106434), .Q(
        n109582) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24374 ), .CK(Clk), .RN(Rst), .Q(n109583)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24342 ), .CK(Clk), .RN(Rst), .Q(n109584)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24310 ), .CK(Clk), .RN(Rst), .Q(n109585)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24278 ), .CK(Clk), .RN(Rst), .Q(n109586), 
        .QN(n102975) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24246 ), .CK(Clk), .RN(Rst), .Q(n109587)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24214 ), .CK(Clk), .RN(Rst), .Q(n109588)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24150 ), .CK(Clk), .RN(Rst), .Q(n109589)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24118 ), .CK(Clk), .RN(Rst), .Q(n109590)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24054 ), .CK(Clk), .RN(n106430), .Q(
        n109591) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24022 ), .CK(Clk), .RN(Rst), .Q(n72580) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23990 ), .CK(Clk), .RN(Rst), .Q(n109592), 
        .QN(n102404) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23958 ), .CK(Clk), .RN(n106486), .Q(
        n109593) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23926 ), .CK(Clk), .RN(n106486), .Q(
        n109594), .QN(n103569) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23894 ), .CK(Clk), .RN(n106486), .Q(
        n109595), .QN(n102973) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23862 ), .CK(Clk), .RN(n106486), .Q(
        n109596) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23798 ), .CK(Clk), .RN(n106486), .Q(
        n109597) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23766 ), .CK(Clk), .RN(n106486), .Q(
        n109598), .QN(n101041) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][11]  ( .D(n104039), 
        .CK(Clk), .RN(n106486), .Q(n109599) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23702 ), .CK(Clk), .RN(n106486), .Q(n72590) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23670 ), .CK(Clk), .RN(n106486), .Q(
        n109600), .QN(n101010) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23638 ), .CK(Clk), .RN(n106486), .Q(n72592) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23606 ), .CK(Clk), .RN(n106486), .Q(
        n109601) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23574 ), .CK(Clk), .RN(n106499), .Q(
        n109602) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23542 ), .CK(Clk), .RN(Rst), .Q(n109603), 
        .QN(n103566) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23510 ), .CK(Clk), .RN(Rst), .Q(n109604)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][11]  ( .D(n104048), 
        .CK(Clk), .RN(n106444), .Q(n72597) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23446 ), .CK(Clk), .RN(n106492), .Q(n72598) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23414 ), .CK(Clk), .RN(Rst), .Q(n109605)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23382 ), .CK(Clk), .RN(Rst), .Q(n72600) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][11]  ( .D(n104064), 
        .CK(Clk), .RN(Rst), .Q(n109606) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23318 ), .CK(Clk), .RN(n106434), .Q(
        n109607) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23254 ), .CK(Clk), .RN(n106496), .Q(
        n109608), .QN(n102971) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23222 ), .CK(Clk), .RN(Rst), .Q(n109609)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23190 ), .CK(Clk), .RN(Rst), .Q(n109610)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23126 ), .CK(Clk), .RN(Rst), .Q(n109611)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][11]  ( .D(n104008), 
        .CK(Clk), .RN(n106494), .Q(n109612) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23062 ), .CK(Clk), .RN(n106415), .Q(
        n109613) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23030 ), .CK(Clk), .RN(n106495), .Q(
        n109614) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22998 ), .CK(Clk), .RN(n106426), .Q(
        n109615) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22966 ), .CK(Clk), .RN(n106460), .Q(
        n109616) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22934 ), .CK(Clk), .RN(Rst), .Q(n72614) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22902 ), .CK(Clk), .RN(Rst), .Q(n72615) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22870 ), .CK(Clk), .RN(n106493), .Q(
        n109617) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22838 ), .CK(Clk), .RN(Rst), .Q(n109618)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22806 ), .CK(Clk), .RN(n106461), .Q(
        n109619) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22774 ), .CK(Clk), .RN(n106399), .Q(
        n109620) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22742 ), .CK(Clk), .RN(Rst), .Q(n72620) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22710 ), .CK(Clk), .RN(Rst), .Q(n109621)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22678 ), .CK(Clk), .RN(n106394), .Q(
        n109622) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22646 ), .CK(Clk), .RN(Rst), .Q(n109623)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22614 ), .CK(Clk), .RN(Rst), .Q(n109624)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22582 ), .CK(Clk), .RN(n106478), .Q(
        n109625) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][11]  ( .D(
        \DLX_Datapath/RegisterFile/N22550 ), .CK(Clk), .RN(n106477), .Q(n72626), .QN(n104522) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25878 ), .CK(Clk), .RN(n106451), .Q(n72627) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][11]  ( .D(n104276), 
        .CK(Clk), .RN(n106450), .Q(n109626) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25942 ), .CK(Clk), .RN(n106506), .Q(
        n109627) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25974 ), .CK(Clk), .RN(Rst), .Q(n109628), 
        .QN(n103578) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26006 ), .CK(Clk), .RN(Rst), .Q(n109629)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26038 ), .CK(Clk), .RN(n106505), .Q(
        n109630) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26070 ), .CK(Clk), .RN(Rst), .Q(n109631)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26102 ), .CK(Clk), .RN(n106407), .Q(n72634) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26134 ), .CK(Clk), .RN(n106504), .Q(
        n109632), .QN(n101857) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26166 ), .CK(Clk), .RN(Rst), .Q(n72636) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26198 ), .CK(Clk), .RN(n106453), .Q(n72637) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26230 ), .CK(Clk), .RN(n106452), .Q(
        n109633) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26262 ), .CK(Clk), .RN(Rst), .Q(n72639) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26294 ), .CK(Clk), .RN(Rst), .Q(n109634)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26326 ), .CK(Clk), .RN(Rst), .Q(n109635)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26358 ), .CK(Clk), .RN(Rst), .Q(n109636)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26390 ), .CK(Clk), .RN(Rst), .Q(n109637)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26454 ), .CK(Clk), .RN(Rst), .Q(n109639)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26486 ), .CK(Clk), .RN(Rst), .Q(n109640), 
        .QN(n103579) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26518 ), .CK(Clk), .RN(Rst), .Q(n109641)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26550 ), .CK(Clk), .RN(Rst), .Q(n109642)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26582 ), .CK(Clk), .RN(Rst), .Q(n109643)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26614 ), .CK(Clk), .RN(Rst), .Q(n109644)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][11]  ( .D(n106970), 
        .CK(Clk), .RN(Rst), .Q(n109645) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26678 ), .CK(Clk), .RN(Rst), .Q(n109646), 
        .QN(n102415) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26710 ), .CK(Clk), .RN(n106485), .Q(
        n109647), .QN(n102983) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26742 ), .CK(Clk), .RN(n106485), .Q(n72654), .QN(n104536) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][11]  ( .D(n107001), 
        .CK(Clk), .RN(n106485), .Q(n109648), .QN(n101858) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26838 ), .CK(Clk), .RN(n106485), .Q(
        n109650), .QN(n102984) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[11]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107073), .Q(
        \DLX_Datapath/next_A_IDEX[11] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[11]  ( .D(n106619), .CK(Clk), .RN(n106485), 
        .Q(n109651) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[11]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [11]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[11]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [11]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [11]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[11]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [11]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [11]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[11]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107039), .Q(
        \DLX_Datapath/next_B_IDEX [11]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[11]  ( .D(n106691), .CK(Clk), .RN(n106485), 
        .Q(n72661) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[11]  ( .D(n58912), .CK(Clk), .RN(n106485), 
        .Q(n109654) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25844 ), .CK(Clk), .RN(n106485), .Q(n72665) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25812 ), .CK(Clk), .RN(n106485), .Q(
        n109655) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25780 ), .CK(Clk), .RN(n106485), .Q(
        n109656) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25748 ), .CK(Clk), .RN(n106484), .Q(
        n109657) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25684 ), .CK(Clk), .RN(n106484), .Q(
        n109658) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25620 ), .CK(Clk), .RN(n106484), .Q(
        n109659) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25588 ), .CK(Clk), .RN(n106484), .Q(
        n109660) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25556 ), .CK(Clk), .RN(n106484), .Q(
        n109661) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25524 ), .CK(Clk), .RN(n106484), .Q(
        n109662) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25492 ), .CK(Clk), .RN(n106484), .Q(
        n109663), .QN(n100583) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25460 ), .CK(Clk), .RN(n106484), .Q(n72677) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25428 ), .CK(Clk), .RN(n106484), .Q(
        n109664) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25396 ), .CK(Clk), .RN(n106484), .Q(
        n109665) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25364 ), .CK(Clk), .RN(n106483), .Q(
        n109666) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][9]  ( .D(n104304), 
        .CK(Clk), .RN(n106483), .Q(n109667) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25300 ), .CK(Clk), .RN(n106483), .Q(
        n109668), .QN(n102943) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25268 ), .CK(Clk), .RN(n106483), .Q(
        n109669), .QN(n102373) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25236 ), .CK(Clk), .RN(n106483), .Q(
        n109670), .QN(n101819) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25204 ), .CK(Clk), .RN(n106483), .Q(
        n109671) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25172 ), .CK(Clk), .RN(n106483), .Q(n72686) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][9]  ( .D(n104199), 
        .CK(Clk), .RN(n106483), .Q(n109672) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25076 ), .CK(Clk), .RN(n106483), .Q(
        n109673) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25044 ), .CK(Clk), .RN(n106483), .Q(n72690), .QN(n104593) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25012 ), .CK(Clk), .RN(n106483), .Q(
        n109674) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24980 ), .CK(Clk), .RN(Rst), .Q(n109675), 
        .QN(n100615) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24948 ), .CK(Clk), .RN(Rst), .Q(n109676)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24916 ), .CK(Clk), .RN(Rst), .Q(n72694) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24884 ), .CK(Clk), .RN(Rst), .Q(n109677), 
        .QN(n101170) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24852 ), .CK(Clk), .RN(Rst), .Q(n109678)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24820 ), .CK(Clk), .RN(Rst), .Q(n109679)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24788 ), .CK(Clk), .RN(Rst), .Q(n72698) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][9]  ( .D(n104183), 
        .CK(Clk), .RN(Rst), .Q(n109680) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][9]  ( .D(n104167), 
        .CK(Clk), .RN(Rst), .Q(n109681) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24660 ), .CK(Clk), .RN(Rst), .Q(n109682), 
        .QN(n102939) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24628 ), .CK(Clk), .RN(Rst), .Q(n72703) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24596 ), .CK(Clk), .RN(Rst), .Q(n109683)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24532 ), .CK(Clk), .RN(Rst), .Q(n109684)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24500 ), .CK(Clk), .RN(n106396), .Q(
        n109685), .QN(n102366) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24468 ), .CK(Clk), .RN(Rst), .Q(n72708), 
        .QN(n104646) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24436 ), .CK(Clk), .RN(n106478), .Q(
        n109686) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24404 ), .CK(Clk), .RN(n106439), .Q(
        n109687) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24372 ), .CK(Clk), .RN(Rst), .Q(n109688)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24340 ), .CK(Clk), .RN(Rst), .Q(n109689)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24308 ), .CK(Clk), .RN(Rst), .Q(n109690)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24276 ), .CK(Clk), .RN(Rst), .Q(n109691), 
        .QN(n102936) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24244 ), .CK(Clk), .RN(Rst), .Q(n109692)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24212 ), .CK(Clk), .RN(Rst), .Q(n109693)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24148 ), .CK(Clk), .RN(Rst), .Q(n109694)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24116 ), .CK(Clk), .RN(Rst), .Q(n109695)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24052 ), .CK(Clk), .RN(Rst), .Q(n109696)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24020 ), .CK(Clk), .RN(Rst), .Q(n72722) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23988 ), .CK(Clk), .RN(Rst), .Q(n109697), 
        .QN(n101067) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23956 ), .CK(Clk), .RN(n106505), .Q(
        n109698) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23924 ), .CK(Clk), .RN(n106505), .Q(
        n109699), .QN(n103533) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23892 ), .CK(Clk), .RN(n106505), .Q(
        n109700), .QN(n102934) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23860 ), .CK(Clk), .RN(n106505), .Q(
        n109701) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][9]  ( .D(n104024), 
        .CK(Clk), .RN(n106505), .Q(n109702) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23764 ), .CK(Clk), .RN(n106505), .Q(
        n109703), .QN(n101043) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23732 ), .CK(Clk), .RN(n106505), .Q(
        n109704) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23700 ), .CK(Clk), .RN(n106505), .Q(n72732) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23668 ), .CK(Clk), .RN(n106505), .Q(
        n109705), .QN(n101012) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23636 ), .CK(Clk), .RN(n106505), .Q(n72734) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23604 ), .CK(Clk), .RN(n106505), .Q(
        n109706) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23572 ), .CK(Clk), .RN(Rst), .Q(n109707)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][9]  ( .D(n104033), 
        .CK(Clk), .RN(Rst), .Q(n109708), .QN(n103530) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23508 ), .CK(Clk), .RN(Rst), .Q(n109709)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23476 ), .CK(Clk), .RN(Rst), .Q(n72739) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23444 ), .CK(Clk), .RN(Rst), .Q(n72740) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23412 ), .CK(Clk), .RN(n106498), .Q(
        n109710) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23380 ), .CK(Clk), .RN(n106499), .Q(
        n109711) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][9]  ( .D(n104061), 
        .CK(Clk), .RN(Rst), .Q(n109712) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23316 ), .CK(Clk), .RN(n106500), .Q(
        n109713) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23252 ), .CK(Clk), .RN(n106496), .Q(
        n109714), .QN(n102932) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23220 ), .CK(Clk), .RN(n106424), .Q(
        n109715) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23188 ), .CK(Clk), .RN(n106478), .Q(
        n109716) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23156 ), .CK(Clk), .RN(Rst), .Q(n109717)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23124 ), .CK(Clk), .RN(n106394), .Q(
        n109718) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23092 ), .CK(Clk), .RN(n106420), .Q(
        n109719) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23060 ), .CK(Clk), .RN(n106402), .Q(
        n109720) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23028 ), .CK(Clk), .RN(Rst), .Q(n109721)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22996 ), .CK(Clk), .RN(n106477), .Q(
        n109722) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22964 ), .CK(Clk), .RN(Rst), .Q(n109723)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22932 ), .CK(Clk), .RN(n106476), .Q(n72756) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22900 ), .CK(Clk), .RN(n106428), .Q(n72757) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22868 ), .CK(Clk), .RN(Rst), .Q(n109724)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22836 ), .CK(Clk), .RN(n106427), .Q(
        n109725) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22804 ), .CK(Clk), .RN(n106504), .Q(
        n109726) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22772 ), .CK(Clk), .RN(n106504), .Q(
        n109727) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22740 ), .CK(Clk), .RN(n106504), .Q(n72762) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22708 ), .CK(Clk), .RN(n106504), .Q(
        n109728) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22676 ), .CK(Clk), .RN(n106504), .Q(
        n109729) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22644 ), .CK(Clk), .RN(n106504), .Q(
        n109730) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22612 ), .CK(Clk), .RN(n106504), .Q(
        n109731) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22580 ), .CK(Clk), .RN(n106504), .Q(
        n109732) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][9]  ( .D(
        \DLX_Datapath/RegisterFile/N22548 ), .CK(Clk), .RN(n106504), .Q(n72768), .QN(n104520) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][9]  ( .D(n104271), 
        .CK(Clk), .RN(n106504), .Q(n109733) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25940 ), .CK(Clk), .RN(n106504), .Q(
        n109734) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25972 ), .CK(Clk), .RN(Rst), .Q(n109735), 
        .QN(n103542) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26004 ), .CK(Clk), .RN(Rst), .Q(n109736)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26036 ), .CK(Clk), .RN(Rst), .Q(n109737)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26068 ), .CK(Clk), .RN(Rst), .Q(n109738)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26100 ), .CK(Clk), .RN(n106505), .Q(n72776) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26132 ), .CK(Clk), .RN(n106507), .Q(
        n109739), .QN(n101823) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26164 ), .CK(Clk), .RN(n106508), .Q(n72778) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26196 ), .CK(Clk), .RN(Rst), .Q(n72779) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26228 ), .CK(Clk), .RN(Rst), .Q(n109740)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26260 ), .CK(Clk), .RN(n106488), .Q(n72781) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26292 ), .CK(Clk), .RN(Rst), .Q(n109741)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26324 ), .CK(Clk), .RN(Rst), .Q(n109742)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26356 ), .CK(Clk), .RN(n106500), .Q(
        n109743) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26388 ), .CK(Clk), .RN(n106499), .Q(
        n109744) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26452 ), .CK(Clk), .RN(Rst), .Q(n109746)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26484 ), .CK(Clk), .RN(n106436), .Q(
        n109747), .QN(n103544) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26516 ), .CK(Clk), .RN(Rst), .Q(n109748)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26548 ), .CK(Clk), .RN(n106503), .Q(
        n109749) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26580 ), .CK(Clk), .RN(Rst), .Q(n109750)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26612 ), .CK(Clk), .RN(n106498), .Q(
        n109751) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][9]  ( .D(n106968), 
        .CK(Clk), .RN(n106497), .Q(n109752) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26676 ), .CK(Clk), .RN(n106496), .Q(
        n109753), .QN(n102375) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26708 ), .CK(Clk), .RN(n106461), .Q(
        n109754), .QN(n102946) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][9]  ( .D(n104322), 
        .CK(Clk), .RN(n106394), .Q(n72796), .QN(n104525) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][9]  ( .D(n106999), 
        .CK(Clk), .RN(n106399), .Q(n109755), .QN(n101824) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26836 ), .CK(Clk), .RN(Rst), .Q(n109757), 
        .QN(n102947) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[9]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107071), .Q(
        \DLX_Datapath/next_A_IDEX[9] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[9]  ( .D(n106604), .CK(Clk), .RN(Rst), .Q(
        n109758) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_mul_reg[9]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [9]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[9]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [9]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [9]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[9]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [9]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [9]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[9]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107037), .Q(
        \DLX_Datapath/next_B_IDEX [9]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[9]  ( .D(n106690), .CK(Clk), .RN(Rst), .Q(
        n72803) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[9]  ( .D(n58910), .CK(Clk), .RN(Rst), .Q(
        n109761) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[9]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [9]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [9]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[9]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [9]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [9]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[9]  ( .D(n107606), .GN(n60159), 
        .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [9]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[8]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N153 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [8]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[9]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N154 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [9]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[8]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N121 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [8]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[9]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N122 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [9]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[10]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [10]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [10]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[10]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [10]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [10]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[10]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107038), .Q(
        \DLX_Datapath/next_B_IDEX [10]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[10]  ( .D(n106669), .CK(Clk), .RN(n106450), 
        .Q(n72808) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[10]  ( .D(n58909), .CK(Clk), .RN(n106451), 
        .Q(n109766) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[10]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [10]), .GN(n105900), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [10]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[10]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N123 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [10]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[12]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N157 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [12]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[10]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [10]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [10]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[10]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N155 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [10]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[10]  ( .D(n107607), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [10]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[11]  ( .D(n107608), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [11]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[12]  ( .D(n104362), .GN(n60159), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [12]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[13]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [13]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [13]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[13]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [13]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [13]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/B_mul_reg[13]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInB [13]), .GN(n105899), .Q(
        \DLX_Datapath/ArithLogUnit/B_mul [13]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[12]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N125 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [12]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[13]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N126 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [13]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[14]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N127 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [14]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[31]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(n106876), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [31]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[29]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(n106841), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [29]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[29]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N174 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [29]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[28]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N173 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [28]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[26]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N139 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [26]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[15]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N128 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [15]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[13]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [13]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [13]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[13]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N158 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [13]) );
  DFFR_X2 \DLX_Datapath/PC_reg[13]  ( .D(n60312), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [1]), .QN(n62194) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[12]  ( .D(n103946), .CK(Clk), .RN(Rst), 
        .Q(n109774) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[13]  ( .D(n103951), .CK(Clk), .RN(n106474), 
        .Q(n109775) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[14]  ( .D(n103937), .CK(Clk), .RN(Rst), 
        .Q(n109776) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[15]  ( .D(n103938), .CK(Clk), .RN(Rst), 
        .Q(n109777) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[13]  ( .D(n107601), .GN(n60159), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [13]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[14]  ( .D(n107602), .GN(n60159), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [14]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[15]  ( .D(n107603), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [15]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[19]  ( .D(n106909), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [19]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[19]  ( .D(n104351), .CK(Clk), .RN(Rst), .Q(DataAddr[19]), .QN(n58596) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[19]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [19]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [19]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[19]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N164 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [19]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[18]  ( .D(n106907), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [18]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[18]  ( .D(n104352), .CK(Clk), .RN(
        n106423), .Q(DataAddr[18]), .QN(n58594) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[18]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [18]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [18]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[18]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N163 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [18]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[16]  ( .D(n104363), .GN(n60159), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [16]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[17]  ( .D(n106905), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [17]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[17]  ( .D(n104353), .CK(Clk), .RN(
        n106424), .Q(DataAddr[17]), .QN(n58592) );
  DFFR_X2 \DLX_Datapath/PC_reg[17]  ( .D(n60308), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [1]), .QN(n59472) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[18]  ( .D(n106531), .CK(Clk), .RN(Rst), 
        .Q(n109783) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[18]  ( .D(n106648), .CK(Clk), .RN(Rst), 
        .Q(n72830) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[18]  ( .D(n58902), .CK(Clk), .RN(Rst), 
        .Q(n109784), .QN(n59341) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25851 ), .CK(Clk), .RN(n106503), .Q(n72833) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25819 ), .CK(Clk), .RN(n106503), .Q(
        n109786) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25787 ), .CK(Clk), .RN(n106503), .Q(
        n109787) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25755 ), .CK(Clk), .RN(n106503), .Q(
        n109788) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25691 ), .CK(Clk), .RN(n106503), .Q(
        n109789) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25627 ), .CK(Clk), .RN(n106503), .Q(
        n109790) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25595 ), .CK(Clk), .RN(n106503), .Q(
        n109791) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25563 ), .CK(Clk), .RN(n106503), .Q(
        n109792) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25531 ), .CK(Clk), .RN(n106503), .Q(
        n109793) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25499 ), .CK(Clk), .RN(n106503), .Q(
        n109794), .QN(n100576) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25467 ), .CK(Clk), .RN(n106502), .Q(n72845) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25435 ), .CK(Clk), .RN(n106502), .Q(
        n109795) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25403 ), .CK(Clk), .RN(n106502), .Q(
        n109796) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25371 ), .CK(Clk), .RN(n106502), .Q(
        n109797) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25339 ), .CK(Clk), .RN(n106502), .Q(
        n109798) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25307 ), .CK(Clk), .RN(n106502), .Q(
        n109799), .QN(n103080) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25275 ), .CK(Clk), .RN(n106502), .Q(
        n109800), .QN(n102507) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25243 ), .CK(Clk), .RN(n106502), .Q(
        n109801), .QN(n101937) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25211 ), .CK(Clk), .RN(n106502), .Q(
        n109802) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25179 ), .CK(Clk), .RN(n106502), .Q(n72854) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25147 ), .CK(Clk), .RN(n106502), .Q(
        n109803) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25083 ), .CK(Clk), .RN(n106501), .Q(
        n109804) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25051 ), .CK(Clk), .RN(n106501), .Q(n72858), .QN(n104600) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25019 ), .CK(Clk), .RN(n106501), .Q(
        n109805) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24987 ), .CK(Clk), .RN(n106501), .Q(
        n109806), .QN(n100608) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24955 ), .CK(Clk), .RN(n106501), .Q(
        n109807) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24923 ), .CK(Clk), .RN(n106501), .Q(n72862) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24891 ), .CK(Clk), .RN(n106501), .Q(
        n109808), .QN(n101163) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24859 ), .CK(Clk), .RN(n106501), .Q(
        n109809) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24827 ), .CK(Clk), .RN(n106501), .Q(
        n109810) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24795 ), .CK(Clk), .RN(n106501), .Q(n72866) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24763 ), .CK(Clk), .RN(n106501), .Q(
        n109811) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24699 ), .CK(Clk), .RN(n106500), .Q(
        n109812) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24667 ), .CK(Clk), .RN(n106500), .Q(
        n109813), .QN(n103076) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24635 ), .CK(Clk), .RN(n106500), .Q(n72871) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24603 ), .CK(Clk), .RN(n106500), .Q(
        n109814) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24539 ), .CK(Clk), .RN(n106500), .Q(
        n109815) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24507 ), .CK(Clk), .RN(n106500), .Q(
        n109816), .QN(n102500) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24475 ), .CK(Clk), .RN(n106500), .Q(n72876), .QN(n104621) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24443 ), .CK(Clk), .RN(n106500), .Q(
        n109817) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24411 ), .CK(Clk), .RN(n106500), .Q(
        n109818) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24379 ), .CK(Clk), .RN(n106500), .Q(
        n109819) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24347 ), .CK(Clk), .RN(n106500), .Q(
        n109820) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24315 ), .CK(Clk), .RN(n106499), .Q(
        n109821) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24283 ), .CK(Clk), .RN(n106501), .Q(
        n109822), .QN(n103073) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24251 ), .CK(Clk), .RN(Rst), .Q(n109823)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24219 ), .CK(Clk), .RN(Rst), .Q(n109824)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24155 ), .CK(Clk), .RN(Rst), .Q(n109825)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24123 ), .CK(Clk), .RN(Rst), .Q(n109826)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24059 ), .CK(Clk), .RN(Rst), .Q(n109827)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24027 ), .CK(Clk), .RN(Rst), .Q(n72890) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23995 ), .CK(Clk), .RN(Rst), .Q(n109828), 
        .QN(n101064) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23963 ), .CK(Clk), .RN(Rst), .Q(n109829)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23931 ), .CK(Clk), .RN(Rst), .Q(n109830), 
        .QN(n103659) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23899 ), .CK(Clk), .RN(Rst), .Q(n109831), 
        .QN(n103071) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23867 ), .CK(Clk), .RN(Rst), .Q(n109832)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23803 ), .CK(Clk), .RN(n106495), .Q(
        n109833) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23771 ), .CK(Clk), .RN(Rst), .Q(n109834), 
        .QN(n101036) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23739 ), .CK(Clk), .RN(Rst), .Q(n109835)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23707 ), .CK(Clk), .RN(Rst), .Q(n72900) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23675 ), .CK(Clk), .RN(Rst), .Q(n109836), 
        .QN(n101005) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23643 ), .CK(Clk), .RN(Rst), .Q(n72902) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23611 ), .CK(Clk), .RN(n106371), .Q(
        n109837) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23579 ), .CK(Clk), .RN(Rst), .Q(n109838)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23547 ), .CK(Clk), .RN(Rst), .Q(n109839), 
        .QN(n103655) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23515 ), .CK(Clk), .RN(Rst), .Q(n109840)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][16]  ( .D(n104049), 
        .CK(Clk), .RN(Rst), .Q(n72907) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23451 ), .CK(Clk), .RN(n106495), .Q(n72908) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23419 ), .CK(Clk), .RN(Rst), .Q(n109841)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23387 ), .CK(Clk), .RN(n106475), .Q(
        n109842) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23355 ), .CK(Clk), .RN(Rst), .Q(n109843)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23323 ), .CK(Clk), .RN(Rst), .Q(n109844)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23291 ), .CK(Clk), .RN(Rst), .Q(n109845)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23259 ), .CK(Clk), .RN(Rst), .Q(n109846), 
        .QN(n103069) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23227 ), .CK(Clk), .RN(Rst), .Q(n109847)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23195 ), .CK(Clk), .RN(Rst), .Q(n109848)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23163 ), .CK(Clk), .RN(Rst), .Q(n109849)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23131 ), .CK(Clk), .RN(Rst), .Q(n109850)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23099 ), .CK(Clk), .RN(n106463), .Q(
        n109851) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23067 ), .CK(Clk), .RN(Rst), .Q(n109852)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23035 ), .CK(Clk), .RN(n106462), .Q(
        n109853) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23003 ), .CK(Clk), .RN(Rst), .Q(n109854)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22971 ), .CK(Clk), .RN(n106426), .Q(
        n109855) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22939 ), .CK(Clk), .RN(Rst), .Q(n72924) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22907 ), .CK(Clk), .RN(Rst), .Q(n72925) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22875 ), .CK(Clk), .RN(Rst), .Q(n109856)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22843 ), .CK(Clk), .RN(Rst), .Q(n109857)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22811 ), .CK(Clk), .RN(Rst), .Q(n109858)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22779 ), .CK(Clk), .RN(Rst), .Q(n109859)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22747 ), .CK(Clk), .RN(Rst), .Q(n72930) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22715 ), .CK(Clk), .RN(Rst), .Q(n109860)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22683 ), .CK(Clk), .RN(Rst), .Q(n109861)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22651 ), .CK(Clk), .RN(Rst), .Q(n109862)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22619 ), .CK(Clk), .RN(Rst), .Q(n109863)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22587 ), .CK(Clk), .RN(Rst), .Q(n109864)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25883 ), .CK(Clk), .RN(Rst), .Q(n72937) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][16]  ( .D(n104274), 
        .CK(Clk), .RN(Rst), .Q(n109866) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25947 ), .CK(Clk), .RN(Rst), .Q(n109867)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25979 ), .CK(Clk), .RN(Rst), .Q(n109868), 
        .QN(n103667) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26011 ), .CK(Clk), .RN(Rst), .Q(n109869)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26043 ), .CK(Clk), .RN(Rst), .Q(n109870)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26075 ), .CK(Clk), .RN(Rst), .Q(n109871)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26107 ), .CK(Clk), .RN(Rst), .Q(n72944) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26139 ), .CK(Clk), .RN(Rst), .Q(n109872), 
        .QN(n101939) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26171 ), .CK(Clk), .RN(Rst), .Q(n72946) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26203 ), .CK(Clk), .RN(Rst), .Q(n72947) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26235 ), .CK(Clk), .RN(Rst), .Q(n109873)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26267 ), .CK(Clk), .RN(Rst), .Q(n72949) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26299 ), .CK(Clk), .RN(Rst), .Q(n109874)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26331 ), .CK(Clk), .RN(Rst), .Q(n109875)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26363 ), .CK(Clk), .RN(Rst), .Q(n109876)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26395 ), .CK(Clk), .RN(Rst), .Q(n109877)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26459 ), .CK(Clk), .RN(Rst), .Q(n109879)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26491 ), .CK(Clk), .RN(Rst), .Q(n109880), 
        .QN(n103669) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26523 ), .CK(Clk), .RN(Rst), .Q(n109881)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26555 ), .CK(Clk), .RN(Rst), .Q(n109882)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26587 ), .CK(Clk), .RN(Rst), .Q(n109883)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26619 ), .CK(Clk), .RN(Rst), .Q(n109884)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][16]  ( .D(n106975), 
        .CK(Clk), .RN(Rst), .Q(n109885) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26683 ), .CK(Clk), .RN(Rst), .Q(n109886), 
        .QN(n102509) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26715 ), .CK(Clk), .RN(Rst), .Q(n109887), 
        .QN(n103083) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26747 ), .CK(Clk), .RN(Rst), .Q(n72964), 
        .QN(n104541) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][16]  ( .D(n107006), 
        .CK(Clk), .RN(Rst), .Q(n109888), .QN(n101940) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26843 ), .CK(Clk), .RN(Rst), .Q(n109890), 
        .QN(n103084) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[16]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107078), .Q(
        \DLX_Datapath/next_A_IDEX[16] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[16]  ( .D(n106608), .CK(Clk), .RN(Rst), .Q(
        n109891) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[16]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107044), .Q(
        \DLX_Datapath/next_B_IDEX [16]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[16]  ( .D(n106672), .CK(Clk), .RN(Rst), .Q(
        n72969), .QN(n104656) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[16]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [16]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [16]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[16]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N161 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [16]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[16]  ( .D(n103918), .GN(n60158), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [16]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[16]  ( .D(n104354), .CK(Clk), .RN(
        n106507), .Q(DataAddr[16]), .QN(n58588) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[16]  ( .D(n58898), .CK(Clk), .RN(n106507), 
        .Q(n109895) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[16]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [16]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [16]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[16]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [16]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [16]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[16]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N129 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [16]) );
  DFFR_X2 \DLX_Datapath/PC_reg[16]  ( .D(n60309), .CK(Clk), .RN(n106507), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [0]), .QN(n59471) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[16]  ( .D(n103952), .CK(Clk), .RN(n106507), 
        .Q(n109897) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[17]  ( .D(n103939), .CK(Clk), .RN(n106507), 
        .Q(n109898) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[16]  ( .D(n106533), .CK(Clk), .RN(n106507), .Q(n109899) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[16]  ( .D(n106647), .CK(Clk), .RN(n106507), .Q(n72978) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[16]  ( .D(n58897), .CK(Clk), .RN(n106507), .Q(n109900), .QN(n59339) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[17]  ( .D(n106532), .CK(Clk), .RN(n106507), .Q(n109901) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[17]  ( .D(n106637), .CK(Clk), .RN(n106507), .Q(n72980) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[17]  ( .D(n58896), .CK(Clk), .RN(n106507), .Q(n109902), .QN(n59340) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25852 ), .CK(Clk), .RN(Rst), .Q(n72983) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25820 ), .CK(Clk), .RN(Rst), .Q(n109904)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25788 ), .CK(Clk), .RN(Rst), .Q(n109905)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25756 ), .CK(Clk), .RN(n106495), .Q(
        n109906) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25692 ), .CK(Clk), .RN(Rst), .Q(n109907)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25628 ), .CK(Clk), .RN(Rst), .Q(n109908)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25596 ), .CK(Clk), .RN(Rst), .Q(n109909)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25564 ), .CK(Clk), .RN(Rst), .Q(n109910)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25532 ), .CK(Clk), .RN(Rst), .Q(n109911)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25500 ), .CK(Clk), .RN(Rst), .Q(n109912), 
        .QN(n100575) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25468 ), .CK(Clk), .RN(Rst), .Q(n72995) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25436 ), .CK(Clk), .RN(Rst), .Q(n109913)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25404 ), .CK(Clk), .RN(Rst), .Q(n109914)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25372 ), .CK(Clk), .RN(Rst), .Q(n109915)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25340 ), .CK(Clk), .RN(Rst), .Q(n109916)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25308 ), .CK(Clk), .RN(Rst), .Q(n109917), 
        .QN(n103100) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25276 ), .CK(Clk), .RN(Rst), .Q(n109918), 
        .QN(n102526) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25244 ), .CK(Clk), .RN(Rst), .Q(n109919), 
        .QN(n101953) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25212 ), .CK(Clk), .RN(Rst), .Q(n109920)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25180 ), .CK(Clk), .RN(Rst), .Q(n73004) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25148 ), .CK(Clk), .RN(Rst), .Q(n109921)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25084 ), .CK(Clk), .RN(n106506), .Q(
        n109922) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25052 ), .CK(Clk), .RN(n106506), .Q(n73008), .QN(n104601) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25020 ), .CK(Clk), .RN(n106506), .Q(
        n109923) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24988 ), .CK(Clk), .RN(n106506), .Q(
        n109924), .QN(n100607) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24956 ), .CK(Clk), .RN(n106506), .Q(
        n109925) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24924 ), .CK(Clk), .RN(n106506), .Q(n73012) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24892 ), .CK(Clk), .RN(n106506), .Q(
        n109926), .QN(n101162) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24860 ), .CK(Clk), .RN(n106506), .Q(
        n109927) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24828 ), .CK(Clk), .RN(n106506), .Q(
        n109928) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24796 ), .CK(Clk), .RN(n106506), .Q(n73016) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24700 ), .CK(Clk), .RN(Rst), .Q(n109929)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24668 ), .CK(Clk), .RN(Rst), .Q(n109930), 
        .QN(n103096) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24636 ), .CK(Clk), .RN(Rst), .Q(n73021) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24604 ), .CK(Clk), .RN(Rst), .Q(n109931)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24540 ), .CK(Clk), .RN(Rst), .Q(n109932)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24508 ), .CK(Clk), .RN(Rst), .Q(n109933), 
        .QN(n102520) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24476 ), .CK(Clk), .RN(Rst), .Q(n73026), 
        .QN(n104622) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24444 ), .CK(Clk), .RN(Rst), .Q(n109934)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24412 ), .CK(Clk), .RN(Rst), .Q(n109935)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24380 ), .CK(Clk), .RN(Rst), .Q(n109936)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24348 ), .CK(Clk), .RN(n106493), .Q(
        n109937) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24316 ), .CK(Clk), .RN(n106493), .Q(
        n109938) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24284 ), .CK(Clk), .RN(n106493), .Q(
        n109939), .QN(n103093) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24252 ), .CK(Clk), .RN(n106493), .Q(
        n109940) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24220 ), .CK(Clk), .RN(n106493), .Q(
        n109941) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24156 ), .CK(Clk), .RN(n106493), .Q(
        n109942) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24124 ), .CK(Clk), .RN(n106493), .Q(
        n109943) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24060 ), .CK(Clk), .RN(n106506), .Q(
        n109944) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24028 ), .CK(Clk), .RN(Rst), .Q(n73040) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23996 ), .CK(Clk), .RN(Rst), .Q(n109945), 
        .QN(n102518) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23964 ), .CK(Clk), .RN(Rst), .Q(n109946)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23932 ), .CK(Clk), .RN(Rst), .Q(n109947), 
        .QN(n103677) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23900 ), .CK(Clk), .RN(Rst), .Q(n109948), 
        .QN(n103091) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23868 ), .CK(Clk), .RN(n106507), .Q(
        n109949) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][17]  ( .D(n104021), 
        .CK(Clk), .RN(Rst), .Q(n109950) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23772 ), .CK(Clk), .RN(Rst), .Q(n109951), 
        .QN(n101035) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23740 ), .CK(Clk), .RN(Rst), .Q(n109952)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23708 ), .CK(Clk), .RN(n106406), .Q(n73050) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23676 ), .CK(Clk), .RN(n106371), .Q(
        n109953), .QN(n101004) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23644 ), .CK(Clk), .RN(Rst), .Q(n73052) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23612 ), .CK(Clk), .RN(Rst), .Q(n109954)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23580 ), .CK(Clk), .RN(Rst), .Q(n109955)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23548 ), .CK(Clk), .RN(Rst), .Q(n109956), 
        .QN(n103673) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23516 ), .CK(Clk), .RN(Rst), .Q(n109957)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][17]  ( .D(n104050), 
        .CK(Clk), .RN(Rst), .Q(n73057) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23452 ), .CK(Clk), .RN(n106448), .Q(n73058) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23420 ), .CK(Clk), .RN(Rst), .Q(n109958)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23388 ), .CK(Clk), .RN(n106427), .Q(
        n109959) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23356 ), .CK(Clk), .RN(Rst), .Q(n109960)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23324 ), .CK(Clk), .RN(n106436), .Q(
        n109961) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23292 ), .CK(Clk), .RN(n106465), .Q(
        n109962) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23260 ), .CK(Clk), .RN(n106472), .Q(
        n109963), .QN(n103089) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23228 ), .CK(Clk), .RN(n106471), .Q(
        n109964) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23196 ), .CK(Clk), .RN(Rst), .Q(n109965)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][17]  ( .D(n104001), 
        .CK(Clk), .RN(n106466), .Q(n109966) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23132 ), .CK(Clk), .RN(n106474), .Q(
        n109967) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23100 ), .CK(Clk), .RN(Rst), .Q(n109968)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23068 ), .CK(Clk), .RN(Rst), .Q(n109969)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23036 ), .CK(Clk), .RN(n106401), .Q(
        n109970) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23004 ), .CK(Clk), .RN(Rst), .Q(n109971)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22972 ), .CK(Clk), .RN(Rst), .Q(n109972)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22940 ), .CK(Clk), .RN(Rst), .Q(n73074) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22908 ), .CK(Clk), .RN(Rst), .Q(n73075) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22876 ), .CK(Clk), .RN(Rst), .Q(n109973)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22844 ), .CK(Clk), .RN(Rst), .Q(n109974)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22812 ), .CK(Clk), .RN(Rst), .Q(n109975)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22780 ), .CK(Clk), .RN(Rst), .Q(n109976)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22748 ), .CK(Clk), .RN(Rst), .Q(n73080) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22716 ), .CK(Clk), .RN(Rst), .Q(n109977)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22684 ), .CK(Clk), .RN(Rst), .Q(n109978)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22652 ), .CK(Clk), .RN(Rst), .Q(n109979)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22620 ), .CK(Clk), .RN(Rst), .Q(n109980)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22588 ), .CK(Clk), .RN(n106430), .Q(
        n109981) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25884 ), .CK(Clk), .RN(Rst), .Q(n73087) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][17]  ( .D(n104279), 
        .CK(Clk), .RN(n106487), .Q(n109983) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25948 ), .CK(Clk), .RN(n106399), .Q(
        n109984) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25980 ), .CK(Clk), .RN(Rst), .Q(n109985), 
        .QN(n103685) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26012 ), .CK(Clk), .RN(n106449), .Q(
        n109986) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26044 ), .CK(Clk), .RN(n106431), .Q(
        n109987) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26076 ), .CK(Clk), .RN(Rst), .Q(n109988)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26108 ), .CK(Clk), .RN(Rst), .Q(n73094) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26140 ), .CK(Clk), .RN(Rst), .Q(n109989), 
        .QN(n101955) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26172 ), .CK(Clk), .RN(n106372), .Q(n73096) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26204 ), .CK(Clk), .RN(Rst), .Q(n73097) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26236 ), .CK(Clk), .RN(n106459), .Q(
        n109990) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26268 ), .CK(Clk), .RN(Rst), .Q(n73099) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26300 ), .CK(Clk), .RN(n106454), .Q(
        n109991) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26332 ), .CK(Clk), .RN(n106453), .Q(
        n109992) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26364 ), .CK(Clk), .RN(n106452), .Q(
        n109993) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26396 ), .CK(Clk), .RN(Rst), .Q(n109994)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26460 ), .CK(Clk), .RN(Rst), .Q(n109996)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26492 ), .CK(Clk), .RN(n106400), .Q(
        n109997), .QN(n103687) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26524 ), .CK(Clk), .RN(n106451), .Q(
        n109998) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26556 ), .CK(Clk), .RN(n106410), .Q(
        n109999) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26588 ), .CK(Clk), .RN(Rst), .Q(n110000)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26620 ), .CK(Clk), .RN(Rst), .Q(n110001)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][17]  ( .D(n106976), 
        .CK(Clk), .RN(Rst), .Q(n110002) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26684 ), .CK(Clk), .RN(Rst), .Q(n110003), 
        .QN(n102528) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26716 ), .CK(Clk), .RN(n106408), .Q(
        n110004), .QN(n103103) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26748 ), .CK(Clk), .RN(Rst), .Q(n73114), 
        .QN(n104542) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][17]  ( .D(n107007), 
        .CK(Clk), .RN(Rst), .Q(n110005), .QN(n101956) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26844 ), .CK(Clk), .RN(Rst), .Q(n110007), 
        .QN(n103104) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[17]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107079), .Q(
        \DLX_Datapath/next_A_IDEX[17] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[17]  ( .D(n106622), .CK(Clk), .RN(n106428), 
        .Q(n110008) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[17]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [17]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [17]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[17]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [17]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [17]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[17]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N130 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [17]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[17]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107045), .Q(
        \DLX_Datapath/next_B_IDEX [17]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[17]  ( .D(n106694), .CK(Clk), .RN(n106405), 
        .Q(n73120), .QN(n104657) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[17]  ( .D(n58894), .CK(Clk), .RN(n106454), 
        .Q(n110010) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[17]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [17]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [17]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[17]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N162 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [17]) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25854 ), .CK(Clk), .RN(n106378), .Q(n73125) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25822 ), .CK(Clk), .RN(n106496), .Q(
        n110013) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25790 ), .CK(Clk), .RN(Rst), .Q(n110014)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25758 ), .CK(Clk), .RN(Rst), .Q(n110015)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25694 ), .CK(Clk), .RN(Rst), .Q(n110016)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25630 ), .CK(Clk), .RN(n106499), .Q(
        n110017) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25598 ), .CK(Clk), .RN(Rst), .Q(n110018)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25566 ), .CK(Clk), .RN(Rst), .Q(n110019)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25534 ), .CK(Clk), .RN(n106374), .Q(
        n110020) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25502 ), .CK(Clk), .RN(n106385), .Q(
        n110021), .QN(n100573) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25470 ), .CK(Clk), .RN(Rst), .Q(n73137) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25438 ), .CK(Clk), .RN(n106448), .Q(
        n110022) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25406 ), .CK(Clk), .RN(n106446), .Q(
        n110023) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25374 ), .CK(Clk), .RN(Rst), .Q(n110024)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][19]  ( .D(n104299), 
        .CK(Clk), .RN(n106447), .Q(n110025) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25310 ), .CK(Clk), .RN(n106377), .Q(
        n110026), .QN(n103138) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25278 ), .CK(Clk), .RN(n106376), .Q(
        n110027), .QN(n102560) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25246 ), .CK(Clk), .RN(n106446), .Q(
        n110028), .QN(n101985) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25214 ), .CK(Clk), .RN(Rst), .Q(n110029)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25182 ), .CK(Clk), .RN(n106375), .Q(n73146) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][19]  ( .D(n104201), 
        .CK(Clk), .RN(Rst), .Q(n110030) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25086 ), .CK(Clk), .RN(n106380), .Q(
        n110031) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25054 ), .CK(Clk), .RN(n106379), .Q(n73150), .QN(n104603) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25022 ), .CK(Clk), .RN(n106378), .Q(
        n110032) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24990 ), .CK(Clk), .RN(Rst), .Q(n110033), 
        .QN(n100605) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24958 ), .CK(Clk), .RN(n106372), .Q(
        n110034) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24926 ), .CK(Clk), .RN(Rst), .Q(n73154) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24894 ), .CK(Clk), .RN(n106391), .Q(
        n110035), .QN(n101160) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24862 ), .CK(Clk), .RN(n106382), .Q(
        n110036) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][19]  ( .D(n104157), 
        .CK(Clk), .RN(Rst), .Q(n110037) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24798 ), .CK(Clk), .RN(n106381), .Q(n73158) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][19]  ( .D(n104163), 
        .CK(Clk), .RN(Rst), .Q(n110038) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24670 ), .CK(Clk), .RN(Rst), .Q(n110039), 
        .QN(n101149) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24638 ), .CK(Clk), .RN(Rst), .Q(n73163) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24606 ), .CK(Clk), .RN(Rst), .Q(n110040)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24542 ), .CK(Clk), .RN(Rst), .Q(n110041)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24510 ), .CK(Clk), .RN(Rst), .Q(n110042), 
        .QN(n102554) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24478 ), .CK(Clk), .RN(n106495), .Q(n73168), .QN(n104624) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][19]  ( .D(n104149), 
        .CK(Clk), .RN(Rst), .Q(n110043) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24414 ), .CK(Clk), .RN(Rst), .Q(n110044)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24382 ), .CK(Clk), .RN(n106492), .Q(
        n110045) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24350 ), .CK(Clk), .RN(n106492), .Q(
        n110046) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24318 ), .CK(Clk), .RN(n106492), .Q(
        n110047) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24286 ), .CK(Clk), .RN(n106492), .Q(
        n110048), .QN(n103133) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24254 ), .CK(Clk), .RN(n106492), .Q(
        n110049) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24222 ), .CK(Clk), .RN(n106492), .Q(
        n110050) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24158 ), .CK(Clk), .RN(n106492), .Q(
        n110051) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24126 ), .CK(Clk), .RN(n106492), .Q(
        n110052) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][19]  ( .D(n104084), 
        .CK(Clk), .RN(n106492), .Q(n110053) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24030 ), .CK(Clk), .RN(n106492), .Q(n73182) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23998 ), .CK(Clk), .RN(Rst), .Q(n110054), 
        .QN(n101062) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23966 ), .CK(Clk), .RN(Rst), .Q(n110055)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][19]  ( .D(n104094), 
        .CK(Clk), .RN(Rst), .Q(n110056), .QN(n103712) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23902 ), .CK(Clk), .RN(Rst), .Q(n110057), 
        .QN(n103131) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23870 ), .CK(Clk), .RN(Rst), .Q(n110058)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][19]  ( .D(n104022), 
        .CK(Clk), .RN(Rst), .Q(n110059) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23774 ), .CK(Clk), .RN(n106499), .Q(
        n110060), .QN(n101033) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23742 ), .CK(Clk), .RN(n106499), .Q(
        n110061) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23710 ), .CK(Clk), .RN(n106499), .Q(n73192) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23678 ), .CK(Clk), .RN(n106499), .Q(
        n110062), .QN(n101002) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23646 ), .CK(Clk), .RN(n106499), .Q(n73194) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23614 ), .CK(Clk), .RN(n106499), .Q(
        n110063) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23582 ), .CK(Clk), .RN(n106499), .Q(
        n110064) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23550 ), .CK(Clk), .RN(n106499), .Q(
        n110065), .QN(n103708) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23518 ), .CK(Clk), .RN(n106499), .Q(
        n110066) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23486 ), .CK(Clk), .RN(n106499), .Q(n73199) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23454 ), .CK(Clk), .RN(Rst), .Q(n73200) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23390 ), .CK(Clk), .RN(n106445), .Q(
        n110067) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23358 ), .CK(Clk), .RN(Rst), .Q(n110068)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23326 ), .CK(Clk), .RN(Rst), .Q(n110069)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23294 ), .CK(Clk), .RN(n106450), .Q(
        n110070) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23262 ), .CK(Clk), .RN(Rst), .Q(n110071), 
        .QN(n103129) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23230 ), .CK(Clk), .RN(n106492), .Q(
        n110072) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23198 ), .CK(Clk), .RN(Rst), .Q(n110073)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23166 ), .CK(Clk), .RN(n106372), .Q(
        n110074) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23134 ), .CK(Clk), .RN(Rst), .Q(n110075)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23102 ), .CK(Clk), .RN(n106485), .Q(
        n110076) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23070 ), .CK(Clk), .RN(Rst), .Q(n110077)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23038 ), .CK(Clk), .RN(n106471), .Q(
        n110078) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23006 ), .CK(Clk), .RN(n106465), .Q(
        n110079) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22974 ), .CK(Clk), .RN(n106470), .Q(
        n110080) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22942 ), .CK(Clk), .RN(n106482), .Q(n73216) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22910 ), .CK(Clk), .RN(n106423), .Q(n73217) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22878 ), .CK(Clk), .RN(n106479), .Q(
        n110081) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22846 ), .CK(Clk), .RN(n106485), .Q(
        n110082) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22814 ), .CK(Clk), .RN(n106460), .Q(
        n110083) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22782 ), .CK(Clk), .RN(n106398), .Q(
        n110084) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22750 ), .CK(Clk), .RN(n106483), .Q(n73222) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22718 ), .CK(Clk), .RN(n106401), .Q(
        n110085) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22686 ), .CK(Clk), .RN(n106466), .Q(
        n110086) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22654 ), .CK(Clk), .RN(Rst), .Q(n110087)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22622 ), .CK(Clk), .RN(Rst), .Q(n110088)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22590 ), .CK(Clk), .RN(Rst), .Q(n110089)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25886 ), .CK(Clk), .RN(Rst), .Q(n73229) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][19]  ( .D(n104272), 
        .CK(Clk), .RN(Rst), .Q(n110091) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25950 ), .CK(Clk), .RN(Rst), .Q(n110092)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25982 ), .CK(Clk), .RN(Rst), .Q(n110093), 
        .QN(n103720) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26014 ), .CK(Clk), .RN(Rst), .Q(n110094)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26046 ), .CK(Clk), .RN(Rst), .Q(n110095)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26078 ), .CK(Clk), .RN(Rst), .Q(n110096)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26110 ), .CK(Clk), .RN(Rst), .Q(n73236) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26142 ), .CK(Clk), .RN(Rst), .Q(n110097), 
        .QN(n101987) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][19]  ( .D(n104247), 
        .CK(Clk), .RN(n106483), .Q(n73238) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26206 ), .CK(Clk), .RN(n106436), .Q(n73239) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26238 ), .CK(Clk), .RN(n106474), .Q(
        n110098) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26270 ), .CK(Clk), .RN(n106472), .Q(n73241) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26302 ), .CK(Clk), .RN(n106471), .Q(
        n110099) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26334 ), .CK(Clk), .RN(n106470), .Q(
        n110100) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26366 ), .CK(Clk), .RN(n106423), .Q(
        n110101) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26398 ), .CK(Clk), .RN(n106489), .Q(
        n110102) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26462 ), .CK(Clk), .RN(n106479), .Q(
        n110104) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26494 ), .CK(Clk), .RN(n106482), .Q(
        n110105), .QN(n103721) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26526 ), .CK(Clk), .RN(n106498), .Q(
        n110106) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26558 ), .CK(Clk), .RN(n106498), .Q(
        n110107) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26590 ), .CK(Clk), .RN(n106498), .Q(
        n110108) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26622 ), .CK(Clk), .RN(n106498), .Q(
        n110109) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][19]  ( .D(n106978), 
        .CK(Clk), .RN(n106498), .Q(n110110) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26686 ), .CK(Clk), .RN(n106498), .Q(
        n110111), .QN(n102562) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26718 ), .CK(Clk), .RN(n106498), .Q(
        n110112), .QN(n103141) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26750 ), .CK(Clk), .RN(n106498), .Q(n73256), .QN(n104544) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][19]  ( .D(n107009), 
        .CK(Clk), .RN(n106498), .Q(n110113), .QN(n101988) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26846 ), .CK(Clk), .RN(n106498), .Q(
        n110115), .QN(n103142) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[19]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107081), .Q(
        \DLX_Datapath/next_A_IDEX[19] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[19]  ( .D(n106623), .CK(Clk), .RN(n106498), 
        .Q(n110116) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[19]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [19]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [19]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[19]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [19]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [19]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[19]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N132 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [19]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[19]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107047), .Q(
        \DLX_Datapath/next_B_IDEX [19]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[19]  ( .D(n106677), .CK(Clk), .RN(n106497), 
        .Q(n73263), .QN(n104659) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[19]  ( .D(n58892), .CK(Clk), .RN(n106497), 
        .Q(n110119) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25853 ), .CK(Clk), .RN(n106497), .Q(n73267) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25821 ), .CK(Clk), .RN(n106497), .Q(
        n110121) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25757 ), .CK(Clk), .RN(n106497), .Q(
        n110122) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25693 ), .CK(Clk), .RN(n106497), .Q(
        n110123) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25629 ), .CK(Clk), .RN(n106497), .Q(
        n110124) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25597 ), .CK(Clk), .RN(n106496), .Q(
        n110125) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25565 ), .CK(Clk), .RN(n106496), .Q(
        n110126) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25533 ), .CK(Clk), .RN(n106496), .Q(
        n110127) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25501 ), .CK(Clk), .RN(n106496), .Q(
        n110128), .QN(n100574) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25469 ), .CK(Clk), .RN(n106496), .Q(n73279) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25437 ), .CK(Clk), .RN(n106496), .Q(
        n110129) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25405 ), .CK(Clk), .RN(n106496), .Q(
        n110130) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25373 ), .CK(Clk), .RN(n106496), .Q(
        n110131) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25341 ), .CK(Clk), .RN(n106496), .Q(
        n110132) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25309 ), .CK(Clk), .RN(n106496), .Q(
        n110133), .QN(n103120) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25277 ), .CK(Clk), .RN(n106496), .Q(
        n110134), .QN(n102543) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25245 ), .CK(Clk), .RN(n106496), .Q(
        n110135), .QN(n101969) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25213 ), .CK(Clk), .RN(Rst), .Q(n110136)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25181 ), .CK(Clk), .RN(Rst), .Q(n73288) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][18]  ( .D(n104202), 
        .CK(Clk), .RN(Rst), .Q(n110137) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25085 ), .CK(Clk), .RN(Rst), .Q(n110138)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25053 ), .CK(Clk), .RN(Rst), .Q(n73292), 
        .QN(n104602) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25021 ), .CK(Clk), .RN(Rst), .Q(n110139)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24989 ), .CK(Clk), .RN(Rst), .Q(n110140), 
        .QN(n100606) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24957 ), .CK(Clk), .RN(Rst), .Q(n110141)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24925 ), .CK(Clk), .RN(Rst), .Q(n73296) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24893 ), .CK(Clk), .RN(Rst), .Q(n110142), 
        .QN(n101161) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24861 ), .CK(Clk), .RN(Rst), .Q(n110143)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24829 ), .CK(Clk), .RN(n106495), .Q(
        n110144) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24797 ), .CK(Clk), .RN(n106495), .Q(n73300) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24701 ), .CK(Clk), .RN(n106495), .Q(
        n110145) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24669 ), .CK(Clk), .RN(n106495), .Q(
        n110146), .QN(n103116) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24637 ), .CK(Clk), .RN(n106495), .Q(n73305) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24605 ), .CK(Clk), .RN(n106495), .Q(
        n110147) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24541 ), .CK(Clk), .RN(n106495), .Q(
        n110148) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24509 ), .CK(Clk), .RN(n106495), .Q(
        n110149), .QN(n102537) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24477 ), .CK(Clk), .RN(n106495), .Q(n73310), .QN(n104623) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24445 ), .CK(Clk), .RN(Rst), .Q(n110150)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24413 ), .CK(Clk), .RN(Rst), .Q(n110151)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24381 ), .CK(Clk), .RN(Rst), .Q(n110152)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24349 ), .CK(Clk), .RN(Rst), .Q(n110153)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24317 ), .CK(Clk), .RN(Rst), .Q(n110154)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24285 ), .CK(Clk), .RN(Rst), .Q(n110155), 
        .QN(n103113) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24253 ), .CK(Clk), .RN(Rst), .Q(n110156)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24221 ), .CK(Clk), .RN(Rst), .Q(n110157)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24157 ), .CK(Clk), .RN(Rst), .Q(n110158)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24125 ), .CK(Clk), .RN(Rst), .Q(n110159)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24061 ), .CK(Clk), .RN(n106494), .Q(
        n110160) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24029 ), .CK(Clk), .RN(n106494), .Q(n73324) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23997 ), .CK(Clk), .RN(n106494), .Q(
        n110161), .QN(n101063) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23965 ), .CK(Clk), .RN(n106494), .Q(
        n110162) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23933 ), .CK(Clk), .RN(n106494), .Q(
        n110163), .QN(n103695) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23901 ), .CK(Clk), .RN(n106494), .Q(
        n110164), .QN(n103111) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23869 ), .CK(Clk), .RN(n106494), .Q(
        n110165) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23805 ), .CK(Clk), .RN(n106494), .Q(
        n110166) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23773 ), .CK(Clk), .RN(n106494), .Q(
        n110167), .QN(n101034) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23741 ), .CK(Clk), .RN(n106494), .Q(
        n110168) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23709 ), .CK(Clk), .RN(n106494), .Q(n73334) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23677 ), .CK(Clk), .RN(Rst), .Q(n110169), 
        .QN(n101003) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23645 ), .CK(Clk), .RN(Rst), .Q(n73336) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23613 ), .CK(Clk), .RN(Rst), .Q(n110170)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23581 ), .CK(Clk), .RN(Rst), .Q(n110171)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23549 ), .CK(Clk), .RN(Rst), .Q(n110172), 
        .QN(n103691) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23517 ), .CK(Clk), .RN(Rst), .Q(n110173)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][18]  ( .D(n104051), 
        .CK(Clk), .RN(Rst), .Q(n73341) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23453 ), .CK(Clk), .RN(Rst), .Q(n73342) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23389 ), .CK(Clk), .RN(Rst), .Q(n110174)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][18]  ( .D(n104067), 
        .CK(Clk), .RN(Rst), .Q(n110175) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23325 ), .CK(Clk), .RN(Rst), .Q(n110176)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23293 ), .CK(Clk), .RN(Rst), .Q(n110177)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23261 ), .CK(Clk), .RN(n106493), .Q(
        n110178), .QN(n103109) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23229 ), .CK(Clk), .RN(n106493), .Q(
        n110179) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23197 ), .CK(Clk), .RN(n106493), .Q(
        n110180) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23165 ), .CK(Clk), .RN(n106493), .Q(
        n110181) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23133 ), .CK(Clk), .RN(n106497), .Q(
        n110182) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23101 ), .CK(Clk), .RN(n106499), .Q(
        n110183) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23069 ), .CK(Clk), .RN(n106459), .Q(
        n110184) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23037 ), .CK(Clk), .RN(Rst), .Q(n110185)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23005 ), .CK(Clk), .RN(Rst), .Q(n110186)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22973 ), .CK(Clk), .RN(Rst), .Q(n110187)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22941 ), .CK(Clk), .RN(Rst), .Q(n73358) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22909 ), .CK(Clk), .RN(n106505), .Q(n73359) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22877 ), .CK(Clk), .RN(Rst), .Q(n110188)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22845 ), .CK(Clk), .RN(Rst), .Q(n110189)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22813 ), .CK(Clk), .RN(Rst), .Q(n110190)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22781 ), .CK(Clk), .RN(Rst), .Q(n110191)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22749 ), .CK(Clk), .RN(Rst), .Q(n73364) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22717 ), .CK(Clk), .RN(Rst), .Q(n110192)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22685 ), .CK(Clk), .RN(Rst), .Q(n110193)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22653 ), .CK(Clk), .RN(Rst), .Q(n110194)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22621 ), .CK(Clk), .RN(Rst), .Q(n110195)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22589 ), .CK(Clk), .RN(Rst), .Q(n110196)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25885 ), .CK(Clk), .RN(Rst), .Q(n73371) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][18]  ( .D(n104278), 
        .CK(Clk), .RN(Rst), .Q(n110198) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25949 ), .CK(Clk), .RN(Rst), .Q(n110199)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25981 ), .CK(Clk), .RN(Rst), .Q(n110200), 
        .QN(n103703) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26013 ), .CK(Clk), .RN(Rst), .Q(n110201)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26045 ), .CK(Clk), .RN(Rst), .Q(n110202)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26077 ), .CK(Clk), .RN(n106469), .Q(
        n110203) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26109 ), .CK(Clk), .RN(n106468), .Q(n73378) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26141 ), .CK(Clk), .RN(n106467), .Q(
        n110204), .QN(n101971) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][18]  ( .D(n104252), 
        .CK(Clk), .RN(n106398), .Q(n73380) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26205 ), .CK(Clk), .RN(n106396), .Q(n73381) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26237 ), .CK(Clk), .RN(n106464), .Q(
        n110205) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26269 ), .CK(Clk), .RN(n106463), .Q(n73383) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26301 ), .CK(Clk), .RN(n106462), .Q(
        n110206) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26333 ), .CK(Clk), .RN(n106372), .Q(
        n110207) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26365 ), .CK(Clk), .RN(Rst), .Q(n110208)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26397 ), .CK(Clk), .RN(Rst), .Q(n110209)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26461 ), .CK(Clk), .RN(n106456), .Q(
        n110211) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26493 ), .CK(Clk), .RN(n106456), .Q(
        n110212), .QN(n103704) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26525 ), .CK(Clk), .RN(n106456), .Q(
        n110213) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26557 ), .CK(Clk), .RN(n106456), .Q(
        n110214) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26589 ), .CK(Clk), .RN(n106456), .Q(
        n110215) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26621 ), .CK(Clk), .RN(n106456), .Q(
        n110216) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][18]  ( .D(n106977), 
        .CK(Clk), .RN(n106456), .Q(n110217) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26685 ), .CK(Clk), .RN(n106456), .Q(
        n110218), .QN(n102545) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26717 ), .CK(Clk), .RN(n106456), .Q(
        n110219), .QN(n103123) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26749 ), .CK(Clk), .RN(n106456), .Q(n73398), .QN(n104543) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][18]  ( .D(n107008), 
        .CK(Clk), .RN(n106456), .Q(n110220), .QN(n101972) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26845 ), .CK(Clk), .RN(Rst), .Q(n110222), 
        .QN(n103124) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[18]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107080), .Q(
        \DLX_Datapath/next_A_IDEX[18] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[18]  ( .D(n106609), .CK(Clk), .RN(Rst), .Q(
        n110223) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[18]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [18]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [18]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[18]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [18]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [18]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[18]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N131 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [18]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[18]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107046), .Q(
        \DLX_Datapath/next_B_IDEX [18]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[18]  ( .D(n106673), .CK(Clk), .RN(Rst), .Q(
        n73405), .QN(n104658) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[18]  ( .D(n58890), .CK(Clk), .RN(Rst), .Q(
        n110226) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[17]  ( .D(n107579), .GN(n60159), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [17]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[18]  ( .D(n107580), .GN(n60159), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [18]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[19]  ( .D(n107581), .GN(n60159), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [19]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[23]  ( .D(n106915), .GN(n106360), 
        .Q(\DLX_Datapath/next_ALUOut_EXMEM [23]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[23]  ( .D(n104355), .CK(Clk), .RN(Rst), .Q(DataAddr[23]), .QN(n58577) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[23]  ( .G(n106369), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [23]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [23]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[23]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N168 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [23]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[22]  ( .D(n106913), .GN(n60158), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [22]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[22]  ( .D(n104356), .CK(Clk), .RN(Rst), .Q(DataAddr[22]), .QN(n58575) );
  DFFR_X2 \DLX_Datapath/PC_reg[22]  ( .D(n60303), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [2]), .QN(n62196) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[22]  ( .D(n106527), .CK(Clk), .RN(Rst), 
        .Q(n110228) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[22]  ( .D(n106650), .CK(Clk), .RN(Rst), 
        .Q(n73411) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[22]  ( .D(n58885), .CK(Clk), .RN(Rst), 
        .Q(n110229), .QN(n59345) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25857 ), .CK(Clk), .RN(n106455), .Q(n73414) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25825 ), .CK(Clk), .RN(n106455), .Q(
        n110231) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25761 ), .CK(Clk), .RN(n106455), .Q(
        n110232) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25697 ), .CK(Clk), .RN(n106455), .Q(
        n110233) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25633 ), .CK(Clk), .RN(n106455), .Q(
        n110234) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25601 ), .CK(Clk), .RN(n106455), .Q(
        n110235) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25569 ), .CK(Clk), .RN(n106455), .Q(
        n110236) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25537 ), .CK(Clk), .RN(n106455), .Q(
        n110237) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25505 ), .CK(Clk), .RN(n106455), .Q(
        n110238), .QN(n100570) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25473 ), .CK(Clk), .RN(n106455), .Q(n73426) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25441 ), .CK(Clk), .RN(Rst), .Q(n110239)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25409 ), .CK(Clk), .RN(Rst), .Q(n110240)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25377 ), .CK(Clk), .RN(n106458), .Q(
        n110241) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][22]  ( .D(n104307), 
        .CK(Clk), .RN(Rst), .Q(n110242) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25313 ), .CK(Clk), .RN(n106457), .Q(
        n110243), .QN(n103196) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25281 ), .CK(Clk), .RN(Rst), .Q(n110244), 
        .QN(n102606) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25249 ), .CK(Clk), .RN(n106393), .Q(
        n110245), .QN(n102036) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25217 ), .CK(Clk), .RN(Rst), .Q(n110246)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25185 ), .CK(Clk), .RN(Rst), .Q(n73435) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25153 ), .CK(Clk), .RN(Rst), .Q(n110247)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25089 ), .CK(Clk), .RN(Rst), .Q(n110248)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25057 ), .CK(Clk), .RN(Rst), .Q(n73439), 
        .QN(n104606) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25025 ), .CK(Clk), .RN(n106480), .Q(
        n110249) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24993 ), .CK(Clk), .RN(Rst), .Q(n110250), 
        .QN(n100602) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24961 ), .CK(Clk), .RN(n106479), .Q(n73442) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24929 ), .CK(Clk), .RN(Rst), .Q(n73443) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24897 ), .CK(Clk), .RN(n106491), .Q(
        n110251), .QN(n101157) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24865 ), .CK(Clk), .RN(Rst), .Q(n110252)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24833 ), .CK(Clk), .RN(Rst), .Q(n110253)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24801 ), .CK(Clk), .RN(Rst), .Q(n73447) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][22]  ( .D(n104165), 
        .CK(Clk), .RN(n106468), .Q(n110254) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24673 ), .CK(Clk), .RN(Rst), .Q(n110255), 
        .QN(n103192) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24641 ), .CK(Clk), .RN(n106436), .Q(n73452) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24609 ), .CK(Clk), .RN(n106401), .Q(
        n110256) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24545 ), .CK(Clk), .RN(n106466), .Q(
        n110257) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24513 ), .CK(Clk), .RN(n106465), .Q(
        n110258), .QN(n102600) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24481 ), .CK(Clk), .RN(Rst), .Q(n73457), 
        .QN(n104627) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][22]  ( .D(n104150), 
        .CK(Clk), .RN(n106469), .Q(n110259) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24417 ), .CK(Clk), .RN(Rst), .Q(n110260)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24385 ), .CK(Clk), .RN(n106397), .Q(
        n110261) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24353 ), .CK(Clk), .RN(n106436), .Q(n73461) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][22]  ( .D(n104102), 
        .CK(Clk), .RN(Rst), .Q(n110262) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24289 ), .CK(Clk), .RN(Rst), .Q(n110263), 
        .QN(n103190) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24257 ), .CK(Clk), .RN(Rst), .Q(n110264)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24225 ), .CK(Clk), .RN(n106429), .Q(
        n110265) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24161 ), .CK(Clk), .RN(n106486), .Q(
        n110266) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24129 ), .CK(Clk), .RN(n106373), .Q(
        n110267) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24065 ), .CK(Clk), .RN(n106496), .Q(
        n110268) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24033 ), .CK(Clk), .RN(Rst), .Q(n73471) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24001 ), .CK(Clk), .RN(n106400), .Q(
        n110269), .QN(n101059) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23969 ), .CK(Clk), .RN(Rst), .Q(n110270)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][22]  ( .D(n104096), 
        .CK(Clk), .RN(Rst), .Q(n110271), .QN(n103763) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23905 ), .CK(Clk), .RN(n106435), .Q(
        n110272), .QN(n103188) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23873 ), .CK(Clk), .RN(Rst), .Q(n73476) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23809 ), .CK(Clk), .RN(n106460), .Q(
        n110273) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23777 ), .CK(Clk), .RN(n106506), .Q(
        n110274), .QN(n101030) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23745 ), .CK(Clk), .RN(Rst), .Q(n110275)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23713 ), .CK(Clk), .RN(n106459), .Q(n73481) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23681 ), .CK(Clk), .RN(n106386), .Q(
        n110276), .QN(n100999) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23649 ), .CK(Clk), .RN(n106391), .Q(n73483) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23617 ), .CK(Clk), .RN(Rst), .Q(n73484) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23585 ), .CK(Clk), .RN(n106447), .Q(
        n110277) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23553 ), .CK(Clk), .RN(n106461), .Q(
        n110278), .QN(n103759) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23521 ), .CK(Clk), .RN(n106496), .Q(
        n110279) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23489 ), .CK(Clk), .RN(Rst), .Q(n73488) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23457 ), .CK(Clk), .RN(Rst), .Q(n73489) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23393 ), .CK(Clk), .RN(Rst), .Q(n110280)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23361 ), .CK(Clk), .RN(n106372), .Q(
        n110281) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23329 ), .CK(Clk), .RN(Rst), .Q(n110282)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23297 ), .CK(Clk), .RN(Rst), .Q(n110283)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23265 ), .CK(Clk), .RN(Rst), .Q(n110284), 
        .QN(n103186) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23233 ), .CK(Clk), .RN(Rst), .Q(n110285)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23201 ), .CK(Clk), .RN(n106372), .Q(
        n110286) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23169 ), .CK(Clk), .RN(Rst), .Q(n110287)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23137 ), .CK(Clk), .RN(n106382), .Q(
        n110288) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][22]  ( .D(n104009), 
        .CK(Clk), .RN(n106456), .Q(n110289) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23073 ), .CK(Clk), .RN(n106381), .Q(
        n110290) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23041 ), .CK(Clk), .RN(Rst), .Q(n110291)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23009 ), .CK(Clk), .RN(n106397), .Q(
        n110292) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22977 ), .CK(Clk), .RN(Rst), .Q(n110293)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22945 ), .CK(Clk), .RN(n106500), .Q(n73505) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22913 ), .CK(Clk), .RN(Rst), .Q(n73506) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22881 ), .CK(Clk), .RN(n106455), .Q(
        n110294) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22849 ), .CK(Clk), .RN(n106434), .Q(
        n110295) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22817 ), .CK(Clk), .RN(n106459), .Q(
        n110296) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22785 ), .CK(Clk), .RN(n106380), .Q(
        n110297) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22753 ), .CK(Clk), .RN(n106402), .Q(n73511) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22721 ), .CK(Clk), .RN(Rst), .Q(n110298)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22689 ), .CK(Clk), .RN(Rst), .Q(n110299)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22657 ), .CK(Clk), .RN(Rst), .Q(n110300)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22625 ), .CK(Clk), .RN(Rst), .Q(n110301)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22593 ), .CK(Clk), .RN(Rst), .Q(n110302)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25889 ), .CK(Clk), .RN(n106506), .Q(n73518) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][22]  ( .D(n104267), 
        .CK(Clk), .RN(n106508), .Q(n110304) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25953 ), .CK(Clk), .RN(n106408), .Q(
        n110305) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25985 ), .CK(Clk), .RN(Rst), .Q(n110306), 
        .QN(n103770) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26017 ), .CK(Clk), .RN(n106459), .Q(
        n110307) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26049 ), .CK(Clk), .RN(n106459), .Q(
        n110308) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26081 ), .CK(Clk), .RN(n106459), .Q(
        n110309) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26113 ), .CK(Clk), .RN(n106459), .Q(n73525) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26145 ), .CK(Clk), .RN(n106459), .Q(
        n110310), .QN(n102040) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][22]  ( .D(n104246), 
        .CK(Clk), .RN(n106459), .Q(n73527) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26209 ), .CK(Clk), .RN(n106459), .Q(n73528) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26241 ), .CK(Clk), .RN(n106459), .Q(
        n110311) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26273 ), .CK(Clk), .RN(n106459), .Q(n73530) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26305 ), .CK(Clk), .RN(n106459), .Q(
        n110312) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26337 ), .CK(Clk), .RN(n106459), .Q(
        n110313) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26369 ), .CK(Clk), .RN(n106459), .Q(
        n110314) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26401 ), .CK(Clk), .RN(n106388), .Q(
        n110315) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26465 ), .CK(Clk), .RN(n106387), .Q(
        n110317) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26497 ), .CK(Clk), .RN(n106386), .Q(
        n110318), .QN(n103771) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26529 ), .CK(Clk), .RN(n106385), .Q(
        n110319) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26561 ), .CK(Clk), .RN(n106425), .Q(
        n110320) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26593 ), .CK(Clk), .RN(n106384), .Q(
        n110321) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26625 ), .CK(Clk), .RN(Rst), .Q(n110322)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][22]  ( .D(n106981), 
        .CK(Clk), .RN(Rst), .Q(n110323) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26689 ), .CK(Clk), .RN(n106383), .Q(
        n110324), .QN(n102608) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26721 ), .CK(Clk), .RN(Rst), .Q(n110325), 
        .QN(n103199) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26753 ), .CK(Clk), .RN(Rst), .Q(n73545), 
        .QN(n104547) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][22]  ( .D(n107012), 
        .CK(Clk), .RN(n106411), .Q(n110326), .QN(n102041) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26849 ), .CK(Clk), .RN(Rst), .Q(n110328), 
        .QN(n103200) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[22]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107084), .Q(
        \DLX_Datapath/next_A_IDEX[22] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[22]  ( .D(n106626), .CK(Clk), .RN(n106405), 
        .Q(n110329) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[22]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [22]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [22]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[22]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [22]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [22]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[22]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N135 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [22]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[22]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107050), .Q(
        \DLX_Datapath/next_B_IDEX [22]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[22]  ( .D(n106680), .CK(Clk), .RN(n106403), 
        .Q(n73552), .QN(n104662) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[22]  ( .D(n58883), .CK(Clk), .RN(n106404), 
        .Q(n110332) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[22]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [22]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [22]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[22]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N167 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [22]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[20]  ( .D(n104364), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [20]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[21]  ( .D(n106911), .GN(n60158), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [21]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[21]  ( .D(n104357), .CK(Clk), .RN(Rst), .Q(DataAddr[21]), .QN(n58570) );
  DFFR_X2 \DLX_Datapath/PC_reg[21]  ( .D(n60304), .CK(Clk), .RN(n106393), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [1]), .QN(n62204) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[20]  ( .D(n106529), .CK(Clk), .RN(n106391), .Q(n110334) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[20]  ( .D(n106638), .CK(Clk), .RN(n106392), .Q(n73558) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[20]  ( .D(n58880), .CK(Clk), .RN(Rst), 
        .Q(n110335), .QN(n59343) );
  DFFR_X2 \DLX_Datapath/NPC_IFID_reg[21]  ( .D(n106528), .CK(Clk), .RN(n106457), .Q(n110336) );
  DFFR_X2 \DLX_Datapath/LPC_IDEX_reg[21]  ( .D(n106649), .CK(Clk), .RN(Rst), 
        .Q(n73560) );
  DFFR_X2 \DLX_Datapath/LPC_EXMEM_reg[21]  ( .D(n58879), .CK(Clk), .RN(n106445), .Q(n110337), .QN(n59344) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25855 ), .CK(Clk), .RN(n106500), .Q(n73563) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25823 ), .CK(Clk), .RN(Rst), .Q(n110339)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25759 ), .CK(Clk), .RN(n106371), .Q(
        n110340) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25695 ), .CK(Clk), .RN(Rst), .Q(n110341)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25631 ), .CK(Clk), .RN(Rst), .Q(n110342)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25599 ), .CK(Clk), .RN(Rst), .Q(n110343)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25567 ), .CK(Clk), .RN(Rst), .Q(n110344)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25535 ), .CK(Clk), .RN(n106375), .Q(
        n110345) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25503 ), .CK(Clk), .RN(n106374), .Q(
        n110346), .QN(n100572) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25471 ), .CK(Clk), .RN(n106386), .Q(n73575) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25439 ), .CK(Clk), .RN(n106383), .Q(
        n110347) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25407 ), .CK(Clk), .RN(n106416), .Q(
        n110348) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25375 ), .CK(Clk), .RN(n106387), .Q(
        n110349) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][20]  ( .D(n104305), 
        .CK(Clk), .RN(Rst), .Q(n110350) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25311 ), .CK(Clk), .RN(Rst), .Q(n110351), 
        .QN(n103158) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25279 ), .CK(Clk), .RN(n106377), .Q(
        n110352), .QN(n102576) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25247 ), .CK(Clk), .RN(n106448), .Q(
        n110353), .QN(n102001) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25215 ), .CK(Clk), .RN(n106376), .Q(
        n110354) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25183 ), .CK(Clk), .RN(n106378), .Q(n73584) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25151 ), .CK(Clk), .RN(Rst), .Q(n110355)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25087 ), .CK(Clk), .RN(n106422), .Q(
        n110356) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25055 ), .CK(Clk), .RN(Rst), .Q(n73588), 
        .QN(n104604) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25023 ), .CK(Clk), .RN(Rst), .Q(n110357)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24991 ), .CK(Clk), .RN(Rst), .Q(n110358), 
        .QN(n100604) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24959 ), .CK(Clk), .RN(n106382), .Q(n73591) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24927 ), .CK(Clk), .RN(n106381), .Q(n73592) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24895 ), .CK(Clk), .RN(n106380), .Q(
        n110359), .QN(n101159) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24863 ), .CK(Clk), .RN(n106379), .Q(
        n110360) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][20]  ( .D(n104158), 
        .CK(Clk), .RN(Rst), .Q(n110361) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24799 ), .CK(Clk), .RN(n106389), .Q(n73596) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][20]  ( .D(n104164), 
        .CK(Clk), .RN(n106476), .Q(n110362) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24671 ), .CK(Clk), .RN(Rst), .Q(n110363), 
        .QN(n103154) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24639 ), .CK(Clk), .RN(n106449), .Q(n73601) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24607 ), .CK(Clk), .RN(n106388), .Q(
        n110364) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24543 ), .CK(Clk), .RN(Rst), .Q(n110365)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24511 ), .CK(Clk), .RN(Rst), .Q(n110366), 
        .QN(n102570) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24479 ), .CK(Clk), .RN(n106435), .Q(n73606), .QN(n104625) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][20]  ( .D(n104141), 
        .CK(Clk), .RN(Rst), .Q(n110367) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24415 ), .CK(Clk), .RN(Rst), .Q(n110368)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24383 ), .CK(Clk), .RN(Rst), .Q(n110369)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24351 ), .CK(Clk), .RN(Rst), .Q(n110370)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][20]  ( .D(n104103), 
        .CK(Clk), .RN(Rst), .Q(n110371) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24287 ), .CK(Clk), .RN(Rst), .Q(n110372), 
        .QN(n103151) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24255 ), .CK(Clk), .RN(n106497), .Q(
        n110373) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24223 ), .CK(Clk), .RN(n106376), .Q(
        n110374) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24159 ), .CK(Clk), .RN(Rst), .Q(n110375)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24127 ), .CK(Clk), .RN(Rst), .Q(n110376)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24063 ), .CK(Clk), .RN(Rst), .Q(n110377)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24031 ), .CK(Clk), .RN(Rst), .Q(n73620) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23999 ), .CK(Clk), .RN(Rst), .Q(n110378), 
        .QN(n101061) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23967 ), .CK(Clk), .RN(n106390), .Q(
        n110379) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][20]  ( .D(n104095), 
        .CK(Clk), .RN(n106397), .Q(n110380), .QN(n103729) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23903 ), .CK(Clk), .RN(Rst), .Q(n110381), 
        .QN(n103149) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23871 ), .CK(Clk), .RN(Rst), .Q(n73625) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23807 ), .CK(Clk), .RN(n106474), .Q(n73627) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23775 ), .CK(Clk), .RN(n106472), .Q(
        n110382), .QN(n101032) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23743 ), .CK(Clk), .RN(n106471), .Q(
        n110383) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23711 ), .CK(Clk), .RN(n106470), .Q(n73630) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23679 ), .CK(Clk), .RN(n106458), .Q(
        n110384), .QN(n101001) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23647 ), .CK(Clk), .RN(n106458), .Q(n73632) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23615 ), .CK(Clk), .RN(n106458), .Q(
        n110385) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23583 ), .CK(Clk), .RN(n106458), .Q(
        n110386) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23551 ), .CK(Clk), .RN(n106458), .Q(
        n110387), .QN(n103726) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23519 ), .CK(Clk), .RN(n106458), .Q(
        n110388) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][20]  ( .D(n104055), 
        .CK(Clk), .RN(n106458), .Q(n73637) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23455 ), .CK(Clk), .RN(n106458), .Q(n73638) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23391 ), .CK(Clk), .RN(n106458), .Q(
        n110389) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][20]  ( .D(n104068), 
        .CK(Clk), .RN(n106458), .Q(n110390) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23327 ), .CK(Clk), .RN(n106458), .Q(
        n110391) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23295 ), .CK(Clk), .RN(n106458), .Q(
        n110392) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23263 ), .CK(Clk), .RN(Rst), .Q(n110393), 
        .QN(n103147) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23231 ), .CK(Clk), .RN(Rst), .Q(n110394)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23199 ), .CK(Clk), .RN(Rst), .Q(n110395)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23167 ), .CK(Clk), .RN(Rst), .Q(n110396)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23135 ), .CK(Clk), .RN(Rst), .Q(n110397)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][20]  ( .D(n104010), 
        .CK(Clk), .RN(Rst), .Q(n110398) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23071 ), .CK(Clk), .RN(Rst), .Q(n110399)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23039 ), .CK(Clk), .RN(Rst), .Q(n110400)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23007 ), .CK(Clk), .RN(Rst), .Q(n110401)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][20]  ( .D(n104016), 
        .CK(Clk), .RN(Rst), .Q(n110402) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22943 ), .CK(Clk), .RN(Rst), .Q(n73654) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22911 ), .CK(Clk), .RN(Rst), .Q(n73655) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22879 ), .CK(Clk), .RN(n106457), .Q(
        n110403) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22847 ), .CK(Clk), .RN(n106457), .Q(
        n110404) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22815 ), .CK(Clk), .RN(n106457), .Q(
        n110405) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22783 ), .CK(Clk), .RN(n106457), .Q(
        n110406) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22751 ), .CK(Clk), .RN(n106457), .Q(n73660) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22719 ), .CK(Clk), .RN(n106457), .Q(
        n110407) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22687 ), .CK(Clk), .RN(n106457), .Q(
        n110408) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22655 ), .CK(Clk), .RN(n106457), .Q(
        n110409) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22623 ), .CK(Clk), .RN(n106457), .Q(
        n110410) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22591 ), .CK(Clk), .RN(n106457), .Q(
        n110411) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25887 ), .CK(Clk), .RN(n106457), .Q(n73667) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25919 ), .CK(Clk), .RN(Rst), .Q(n110413)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25951 ), .CK(Clk), .RN(Rst), .Q(n110414)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25983 ), .CK(Clk), .RN(n106392), .Q(
        n110415), .QN(n103736) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26015 ), .CK(Clk), .RN(n106411), .Q(
        n110416) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26047 ), .CK(Clk), .RN(n106410), .Q(
        n110417) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26079 ), .CK(Clk), .RN(n106409), .Q(
        n110418) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26111 ), .CK(Clk), .RN(n106408), .Q(n73674) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26143 ), .CK(Clk), .RN(n106407), .Q(
        n110419), .QN(n102005) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][20]  ( .D(n104248), 
        .CK(Clk), .RN(n106404), .Q(n73676) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26207 ), .CK(Clk), .RN(n106418), .Q(n73677) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26239 ), .CK(Clk), .RN(Rst), .Q(n110420)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26271 ), .CK(Clk), .RN(n106406), .Q(n73679) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26303 ), .CK(Clk), .RN(Rst), .Q(n110421)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26335 ), .CK(Clk), .RN(n106405), .Q(
        n110422) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26367 ), .CK(Clk), .RN(n106451), .Q(
        n110423) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26399 ), .CK(Clk), .RN(n106451), .Q(
        n110424) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26463 ), .CK(Clk), .RN(n106451), .Q(
        n110426) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26495 ), .CK(Clk), .RN(n106451), .Q(
        n110427), .QN(n103737) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26527 ), .CK(Clk), .RN(n106451), .Q(
        n110428) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26559 ), .CK(Clk), .RN(n106451), .Q(
        n110429) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26591 ), .CK(Clk), .RN(n106451), .Q(
        n110430) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26623 ), .CK(Clk), .RN(n106451), .Q(
        n110431) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][20]  ( .D(n106979), 
        .CK(Clk), .RN(n106451), .Q(n110432) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26687 ), .CK(Clk), .RN(n106451), .Q(
        n110433), .QN(n102578) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26719 ), .CK(Clk), .RN(n106451), .Q(
        n110434), .QN(n103161) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26751 ), .CK(Clk), .RN(n106450), .Q(n73694), .QN(n104545) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][20]  ( .D(n107010), 
        .CK(Clk), .RN(n106450), .Q(n110435), .QN(n102006) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26847 ), .CK(Clk), .RN(n106450), .Q(
        n110437), .QN(n103162) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[20]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107082), .Q(
        \DLX_Datapath/next_A_IDEX[20] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[20]  ( .D(n106624), .CK(Clk), .RN(n106450), 
        .Q(n110438) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[20]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107048), .Q(
        \DLX_Datapath/next_B_IDEX [20]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[20]  ( .D(n106678), .CK(Clk), .RN(n106450), 
        .Q(n73699), .QN(n104660) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[20]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [20]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [20]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[20]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N165 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [20]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Z_reg[20]  ( .D(n103917), .GN(n60158), .Q(
        \DLX_Datapath/next_ALUOut_EXMEM [20]) );
  DFFR_X2 \DLX_Datapath/ALUOut_EXMEM_reg[20]  ( .D(n104358), .CK(Clk), .RN(
        n106450), .Q(DataAddr[20]), .QN(n58565) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[20]  ( .D(n58875), .CK(Clk), .RN(n106450), 
        .Q(n110439) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[20]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [20]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [20]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[20]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [20]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [20]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[20]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N133 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [20]) );
  DFFR_X2 \DLX_Datapath/PC_reg[20]  ( .D(n60305), .CK(Clk), .RN(n106450), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [0]), .QN(n62185) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[20]  ( .D(n60273), .CK(Clk), .RN(n106450), 
        .Q(n110443) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[21]  ( .D(n60272), .CK(Clk), .RN(n106450), 
        .Q(n110444) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[22]  ( .D(n60271), .CK(Clk), .RN(n106450), 
        .Q(n110445) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[23]  ( .D(n60270), .CK(Clk), .RN(n106476), 
        .Q(n110446) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25858 ), .CK(Clk), .RN(n106416), .Q(n73710) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25826 ), .CK(Clk), .RN(Rst), .Q(n110448)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25794 ), .CK(Clk), .RN(n106417), .Q(
        n110449) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25762 ), .CK(Clk), .RN(n106413), .Q(
        n110450) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25698 ), .CK(Clk), .RN(Rst), .Q(n110451)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25634 ), .CK(Clk), .RN(n106414), .Q(
        n110452) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25602 ), .CK(Clk), .RN(n106415), .Q(
        n110453) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25570 ), .CK(Clk), .RN(Rst), .Q(n110454)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25538 ), .CK(Clk), .RN(Rst), .Q(n110455)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25506 ), .CK(Clk), .RN(Rst), .Q(n110456), 
        .QN(n100569) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25474 ), .CK(Clk), .RN(Rst), .Q(n73722) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25442 ), .CK(Clk), .RN(Rst), .Q(n110457)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25410 ), .CK(Clk), .RN(Rst), .Q(n110458)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25378 ), .CK(Clk), .RN(Rst), .Q(n110459)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25346 ), .CK(Clk), .RN(Rst), .Q(n110460)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25314 ), .CK(Clk), .RN(Rst), .Q(n110461), 
        .QN(n103214) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25282 ), .CK(Clk), .RN(Rst), .Q(n110462), 
        .QN(n102620) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25250 ), .CK(Clk), .RN(Rst), .Q(n110463), 
        .QN(n102052) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25218 ), .CK(Clk), .RN(Rst), .Q(n110464)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25186 ), .CK(Clk), .RN(Rst), .Q(n73731) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25154 ), .CK(Clk), .RN(Rst), .Q(n110465)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25090 ), .CK(Clk), .RN(Rst), .Q(n110466)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25058 ), .CK(Clk), .RN(Rst), .Q(n73735), 
        .QN(n104607) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25026 ), .CK(Clk), .RN(Rst), .Q(n110467)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24994 ), .CK(Clk), .RN(Rst), .Q(n110468), 
        .QN(n100601) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24962 ), .CK(Clk), .RN(Rst), .Q(n73738) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24930 ), .CK(Clk), .RN(n106385), .Q(n73739) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24898 ), .CK(Clk), .RN(n106417), .Q(
        n110469), .QN(n101156) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24866 ), .CK(Clk), .RN(n106386), .Q(
        n110470) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24834 ), .CK(Clk), .RN(n106387), .Q(
        n110471) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24802 ), .CK(Clk), .RN(Rst), .Q(n73743) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24706 ), .CK(Clk), .RN(Rst), .Q(n110472)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24674 ), .CK(Clk), .RN(n106448), .Q(
        n110473), .QN(n103211) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24642 ), .CK(Clk), .RN(Rst), .Q(n73748) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24610 ), .CK(Clk), .RN(n106440), .Q(
        n110474) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24546 ), .CK(Clk), .RN(Rst), .Q(n110475)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24514 ), .CK(Clk), .RN(n106424), .Q(
        n110476), .QN(n102614) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24482 ), .CK(Clk), .RN(Rst), .Q(n73753), 
        .QN(n104628) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24450 ), .CK(Clk), .RN(Rst), .Q(n110477)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24418 ), .CK(Clk), .RN(Rst), .Q(n110478)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24386 ), .CK(Clk), .RN(Rst), .Q(n110479)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24354 ), .CK(Clk), .RN(Rst), .Q(n73757) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24322 ), .CK(Clk), .RN(Rst), .Q(n110480)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24290 ), .CK(Clk), .RN(Rst), .Q(n110481), 
        .QN(n103209) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24258 ), .CK(Clk), .RN(Rst), .Q(n110482)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24226 ), .CK(Clk), .RN(Rst), .Q(n110483)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24162 ), .CK(Clk), .RN(Rst), .Q(n110484)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24130 ), .CK(Clk), .RN(Rst), .Q(n110485)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24034 ), .CK(Clk), .RN(n106405), .Q(n73767) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24002 ), .CK(Clk), .RN(n106374), .Q(
        n110486), .QN(n101058) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23970 ), .CK(Clk), .RN(n106375), .Q(
        n110487) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23938 ), .CK(Clk), .RN(Rst), .Q(n110488), 
        .QN(n103780) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23906 ), .CK(Clk), .RN(n106376), .Q(
        n110489), .QN(n103207) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23874 ), .CK(Clk), .RN(n106377), .Q(n73772) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23810 ), .CK(Clk), .RN(n106445), .Q(
        n110490) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23778 ), .CK(Clk), .RN(n106446), .Q(
        n110491), .QN(n101029) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23746 ), .CK(Clk), .RN(n106447), .Q(
        n110492) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23714 ), .CK(Clk), .RN(n106448), .Q(n73777) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23682 ), .CK(Clk), .RN(Rst), .Q(n110493), 
        .QN(n100998) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23650 ), .CK(Clk), .RN(Rst), .Q(n73779) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23618 ), .CK(Clk), .RN(Rst), .Q(n73780) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23586 ), .CK(Clk), .RN(Rst), .Q(n110494)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23522 ), .CK(Clk), .RN(n106421), .Q(
        n110495) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][23]  ( .D(n104057), 
        .CK(Clk), .RN(n106379), .Q(n73784) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23458 ), .CK(Clk), .RN(Rst), .Q(n73785) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23426 ), .CK(Clk), .RN(n106378), .Q(
        n110496) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23394 ), .CK(Clk), .RN(n106388), .Q(
        n110497) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][23]  ( .D(n104062), 
        .CK(Clk), .RN(n106380), .Q(n110498) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23330 ), .CK(Clk), .RN(n106447), .Q(
        n110499) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23298 ), .CK(Clk), .RN(n106452), .Q(
        n110500) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23266 ), .CK(Clk), .RN(Rst), .Q(n110501), 
        .QN(n103205) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23234 ), .CK(Clk), .RN(Rst), .Q(n110502)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23202 ), .CK(Clk), .RN(Rst), .Q(n110503)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23170 ), .CK(Clk), .RN(Rst), .Q(n110504)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23138 ), .CK(Clk), .RN(Rst), .Q(n110505)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23106 ), .CK(Clk), .RN(Rst), .Q(n110506)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23074 ), .CK(Clk), .RN(Rst), .Q(n110507)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23042 ), .CK(Clk), .RN(Rst), .Q(n110508)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23010 ), .CK(Clk), .RN(Rst), .Q(n110509)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22978 ), .CK(Clk), .RN(Rst), .Q(n110510)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22946 ), .CK(Clk), .RN(Rst), .Q(n73801) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22914 ), .CK(Clk), .RN(Rst), .Q(n73802) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22882 ), .CK(Clk), .RN(Rst), .Q(n110511)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22850 ), .CK(Clk), .RN(n106449), .Q(
        n110512) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22818 ), .CK(Clk), .RN(n106449), .Q(n73805) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22786 ), .CK(Clk), .RN(n106449), .Q(
        n110513) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22754 ), .CK(Clk), .RN(n106449), .Q(n73807) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22722 ), .CK(Clk), .RN(n106449), .Q(
        n110514) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22690 ), .CK(Clk), .RN(n106449), .Q(
        n110515) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][23]  ( .D(n103956), 
        .CK(Clk), .RN(n106449), .Q(n110516) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22626 ), .CK(Clk), .RN(n106449), .Q(
        n110517) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22594 ), .CK(Clk), .RN(n106449), .Q(n73812) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25890 ), .CK(Clk), .RN(n106449), .Q(n73814) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25922 ), .CK(Clk), .RN(n106449), .Q(
        n110519) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25954 ), .CK(Clk), .RN(Rst), .Q(n110520)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25986 ), .CK(Clk), .RN(Rst), .Q(n110521), 
        .QN(n103787) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26018 ), .CK(Clk), .RN(Rst), .Q(n110522)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26050 ), .CK(Clk), .RN(n106448), .Q(
        n110523) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26082 ), .CK(Clk), .RN(Rst), .Q(n110524)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26114 ), .CK(Clk), .RN(n106395), .Q(n73821) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26146 ), .CK(Clk), .RN(Rst), .Q(n110525), 
        .QN(n102056) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26178 ), .CK(Clk), .RN(Rst), .Q(n73823) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26210 ), .CK(Clk), .RN(Rst), .Q(n73824) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26242 ), .CK(Clk), .RN(n106449), .Q(
        n110526) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26274 ), .CK(Clk), .RN(n106422), .Q(n73826) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26306 ), .CK(Clk), .RN(n106421), .Q(
        n110527) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26338 ), .CK(Clk), .RN(Rst), .Q(n110528)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26370 ), .CK(Clk), .RN(Rst), .Q(n110529)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26402 ), .CK(Clk), .RN(Rst), .Q(n110530)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26466 ), .CK(Clk), .RN(Rst), .Q(n110532)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26498 ), .CK(Clk), .RN(Rst), .Q(n110533), 
        .QN(n103788) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26530 ), .CK(Clk), .RN(Rst), .Q(n110534)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26562 ), .CK(Clk), .RN(Rst), .Q(n110535)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26594 ), .CK(Clk), .RN(Rst), .Q(n110536)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26626 ), .CK(Clk), .RN(Rst), .Q(n110537)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][23]  ( .D(n106982), 
        .CK(Clk), .RN(n106437), .Q(n110538) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26690 ), .CK(Clk), .RN(n106432), .Q(
        n110539), .QN(n102622) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26722 ), .CK(Clk), .RN(n106398), .Q(
        n110540), .QN(n103217) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26754 ), .CK(Clk), .RN(Rst), .Q(n73841), 
        .QN(n104548) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][23]  ( .D(n107013), 
        .CK(Clk), .RN(Rst), .Q(n110541), .QN(n102057) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26850 ), .CK(Clk), .RN(n106439), .Q(
        n110543), .QN(n103218) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[23]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107085), .Q(
        \DLX_Datapath/next_A_IDEX[23] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[23]  ( .D(n106610), .CK(Clk), .RN(Rst), .Q(
        n110544) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[23]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [23]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [23]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[23]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [23]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [23]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[23]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N136 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [23]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[23]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107051), .Q(
        \DLX_Datapath/next_B_IDEX [23]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[23]  ( .D(n106681), .CK(Clk), .RN(n106433), 
        .Q(n73847), .QN(n104663) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[23]  ( .D(n58873), .CK(Clk), .RN(Rst), .Q(
        n110546) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25856 ), .CK(Clk), .RN(n106438), .Q(n73851) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25824 ), .CK(Clk), .RN(n106489), .Q(
        n110548) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25760 ), .CK(Clk), .RN(n106400), .Q(
        n110549) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25696 ), .CK(Clk), .RN(n106451), .Q(
        n110550) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25632 ), .CK(Clk), .RN(n106450), .Q(
        n110551) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25600 ), .CK(Clk), .RN(n106439), .Q(
        n110552) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25568 ), .CK(Clk), .RN(Rst), .Q(n110553)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25536 ), .CK(Clk), .RN(Rst), .Q(n110554)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25504 ), .CK(Clk), .RN(n106401), .Q(
        n110555), .QN(n100571) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25472 ), .CK(Clk), .RN(Rst), .Q(n73863) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25440 ), .CK(Clk), .RN(Rst), .Q(n110556)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25408 ), .CK(Clk), .RN(Rst), .Q(n110557)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25376 ), .CK(Clk), .RN(Rst), .Q(n110558)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25344 ), .CK(Clk), .RN(Rst), .Q(n110559)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25312 ), .CK(Clk), .RN(n106371), .Q(
        n110560), .QN(n103177) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25280 ), .CK(Clk), .RN(Rst), .Q(n110561), 
        .QN(n102591) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25248 ), .CK(Clk), .RN(n106454), .Q(
        n110562), .QN(n102019) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25216 ), .CK(Clk), .RN(n106494), .Q(
        n110563) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25184 ), .CK(Clk), .RN(Rst), .Q(n73872) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25152 ), .CK(Clk), .RN(n106371), .Q(
        n110564) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25088 ), .CK(Clk), .RN(n106386), .Q(
        n110565) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25056 ), .CK(Clk), .RN(n106493), .Q(n73876), .QN(n104605) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25024 ), .CK(Clk), .RN(Rst), .Q(n110566)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24992 ), .CK(Clk), .RN(n106386), .Q(
        n110567), .QN(n100603) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24960 ), .CK(Clk), .RN(Rst), .Q(n73879) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24928 ), .CK(Clk), .RN(n106493), .Q(n73880) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24896 ), .CK(Clk), .RN(n106409), .Q(
        n110568), .QN(n101158) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24864 ), .CK(Clk), .RN(Rst), .Q(n110569)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24832 ), .CK(Clk), .RN(Rst), .Q(n110570)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24800 ), .CK(Clk), .RN(n106385), .Q(n73884) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24704 ), .CK(Clk), .RN(n106506), .Q(
        n110571) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24672 ), .CK(Clk), .RN(Rst), .Q(n110572), 
        .QN(n103173) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24640 ), .CK(Clk), .RN(Rst), .Q(n73889) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24608 ), .CK(Clk), .RN(n106372), .Q(
        n110573) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24544 ), .CK(Clk), .RN(Rst), .Q(n110574)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24512 ), .CK(Clk), .RN(n106414), .Q(
        n110575), .QN(n102585) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24480 ), .CK(Clk), .RN(n106384), .Q(n73894), .QN(n104626) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24448 ), .CK(Clk), .RN(n106504), .Q(
        n110576) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24416 ), .CK(Clk), .RN(Rst), .Q(n110577)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24384 ), .CK(Clk), .RN(Rst), .Q(n110578)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24352 ), .CK(Clk), .RN(n106372), .Q(
        n110579) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24320 ), .CK(Clk), .RN(n106371), .Q(
        n110580) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24288 ), .CK(Clk), .RN(Rst), .Q(n110581), 
        .QN(n103171) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24256 ), .CK(Clk), .RN(n106454), .Q(
        n110582) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24224 ), .CK(Clk), .RN(n106454), .Q(
        n110583) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24160 ), .CK(Clk), .RN(n106454), .Q(
        n110584) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24128 ), .CK(Clk), .RN(n106454), .Q(
        n110585) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24064 ), .CK(Clk), .RN(n106454), .Q(
        n110586) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24032 ), .CK(Clk), .RN(n106454), .Q(n73908) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24000 ), .CK(Clk), .RN(n106454), .Q(
        n110587), .QN(n101060) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23968 ), .CK(Clk), .RN(n106454), .Q(
        n110588) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23936 ), .CK(Clk), .RN(n106454), .Q(
        n110589), .QN(n103746) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23904 ), .CK(Clk), .RN(n106453), .Q(
        n110590), .QN(n103169) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23872 ), .CK(Clk), .RN(n106453), .Q(n73913) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23808 ), .CK(Clk), .RN(n106453), .Q(
        n110591) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23776 ), .CK(Clk), .RN(n106453), .Q(
        n110592), .QN(n101031) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23744 ), .CK(Clk), .RN(n106453), .Q(
        n110593) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23712 ), .CK(Clk), .RN(n106453), .Q(n73918) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23680 ), .CK(Clk), .RN(n106453), .Q(
        n110594), .QN(n101000) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23648 ), .CK(Clk), .RN(n106453), .Q(n73920) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][21]  ( .D(n104043), 
        .CK(Clk), .RN(n106453), .Q(n110595) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23584 ), .CK(Clk), .RN(n106453), .Q(
        n110596) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23552 ), .CK(Clk), .RN(n106453), .Q(
        n110597), .QN(n103742) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23520 ), .CK(Clk), .RN(n106452), .Q(
        n110598) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][21]  ( .D(n104056), 
        .CK(Clk), .RN(n106452), .Q(n73925) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23456 ), .CK(Clk), .RN(n106452), .Q(n73926) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23424 ), .CK(Clk), .RN(n106452), .Q(
        n110599) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23392 ), .CK(Clk), .RN(n106452), .Q(
        n110600) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][21]  ( .D(n104070), 
        .CK(Clk), .RN(n106452), .Q(n110601) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23328 ), .CK(Clk), .RN(n106452), .Q(
        n110602) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23296 ), .CK(Clk), .RN(n106452), .Q(
        n110603) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23264 ), .CK(Clk), .RN(n106452), .Q(
        n110604), .QN(n103167) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23232 ), .CK(Clk), .RN(n106452), .Q(
        n110605) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23200 ), .CK(Clk), .RN(n106452), .Q(
        n110606) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23168 ), .CK(Clk), .RN(n106452), .Q(
        n110607) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23136 ), .CK(Clk), .RN(Rst), .Q(n110608)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23104 ), .CK(Clk), .RN(Rst), .Q(n110609)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23072 ), .CK(Clk), .RN(Rst), .Q(n110610)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23040 ), .CK(Clk), .RN(Rst), .Q(n110611)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23008 ), .CK(Clk), .RN(Rst), .Q(n110612)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22976 ), .CK(Clk), .RN(Rst), .Q(n110613)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22944 ), .CK(Clk), .RN(Rst), .Q(n73942) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22912 ), .CK(Clk), .RN(Rst), .Q(n73943) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22880 ), .CK(Clk), .RN(Rst), .Q(n110614)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22848 ), .CK(Clk), .RN(Rst), .Q(n110615)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22816 ), .CK(Clk), .RN(Rst), .Q(n110616)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22784 ), .CK(Clk), .RN(Rst), .Q(n110617)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22752 ), .CK(Clk), .RN(Rst), .Q(n110618)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22720 ), .CK(Clk), .RN(Rst), .Q(n110619)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22688 ), .CK(Clk), .RN(Rst), .Q(n110620)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22656 ), .CK(Clk), .RN(Rst), .Q(n110621)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22624 ), .CK(Clk), .RN(Rst), .Q(n110622)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22592 ), .CK(Clk), .RN(Rst), .Q(n73953) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25888 ), .CK(Clk), .RN(Rst), .Q(n73955) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25920 ), .CK(Clk), .RN(Rst), .Q(n110624)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25952 ), .CK(Clk), .RN(Rst), .Q(n110625)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25984 ), .CK(Clk), .RN(Rst), .Q(n110626), 
        .QN(n103753) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26016 ), .CK(Clk), .RN(Rst), .Q(n110627)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26048 ), .CK(Clk), .RN(Rst), .Q(n110628)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26080 ), .CK(Clk), .RN(Rst), .Q(n110629)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26112 ), .CK(Clk), .RN(Rst), .Q(n73962) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26144 ), .CK(Clk), .RN(Rst), .Q(n110630), 
        .QN(n102023) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26176 ), .CK(Clk), .RN(Rst), .Q(n73964) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26208 ), .CK(Clk), .RN(n106416), .Q(n73965) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26240 ), .CK(Clk), .RN(Rst), .Q(n110631)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26272 ), .CK(Clk), .RN(Rst), .Q(n73967) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26304 ), .CK(Clk), .RN(Rst), .Q(n110632)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26336 ), .CK(Clk), .RN(Rst), .Q(n110633)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26368 ), .CK(Clk), .RN(n106415), .Q(
        n110634) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26400 ), .CK(Clk), .RN(Rst), .Q(n110635)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26464 ), .CK(Clk), .RN(Rst), .Q(n110637)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26496 ), .CK(Clk), .RN(Rst), .Q(n110638), 
        .QN(n103754) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26528 ), .CK(Clk), .RN(Rst), .Q(n110639)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26560 ), .CK(Clk), .RN(Rst), .Q(n110640)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26592 ), .CK(Clk), .RN(Rst), .Q(n110641)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26624 ), .CK(Clk), .RN(Rst), .Q(n110642)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][21]  ( .D(n106980), 
        .CK(Clk), .RN(Rst), .Q(n110643) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26688 ), .CK(Clk), .RN(Rst), .Q(n110644), 
        .QN(n102593) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26720 ), .CK(Clk), .RN(Rst), .Q(n110645), 
        .QN(n103180) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26752 ), .CK(Clk), .RN(Rst), .Q(n73982), 
        .QN(n104546) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][21]  ( .D(n107011), 
        .CK(Clk), .RN(Rst), .Q(n110646), .QN(n102024) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26848 ), .CK(Clk), .RN(n106454), .Q(
        n110648), .QN(n103181) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[21]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107083), .Q(
        \DLX_Datapath/next_A_IDEX[21] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[21]  ( .D(n106625), .CK(Clk), .RN(Rst), .Q(
        n110649) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[21]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [21]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [21]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[21]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [21]), .GN(n106949), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [21]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[21]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N134 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [21]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[21]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107049), .Q(
        \DLX_Datapath/next_B_IDEX [21]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[21]  ( .D(n106679), .CK(Clk), .RN(Rst), .Q(
        n73988), .QN(n104661) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[21]  ( .D(n58871), .CK(Clk), .RN(Rst), .Q(
        n110652) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[21]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [21]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [21]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[21]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N166 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [21]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[21]  ( .D(n107583), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [21]) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25862 ), .CK(Clk), .RN(n106494), .Q(n73993) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25830 ), .CK(Clk), .RN(n106408), .Q(
        n110655) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25798 ), .CK(Clk), .RN(Rst), .Q(n110656)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25766 ), .CK(Clk), .RN(Rst), .Q(n110657)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25702 ), .CK(Clk), .RN(n106423), .Q(
        n110658) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25638 ), .CK(Clk), .RN(Rst), .Q(n110659)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25606 ), .CK(Clk), .RN(n106412), .Q(
        n110660) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25574 ), .CK(Clk), .RN(n106505), .Q(
        n110661) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25542 ), .CK(Clk), .RN(Rst), .Q(n110662)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25510 ), .CK(Clk), .RN(Rst), .Q(n110663), 
        .QN(n100565) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25478 ), .CK(Clk), .RN(Rst), .Q(n74005) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25446 ), .CK(Clk), .RN(Rst), .Q(n110664)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25414 ), .CK(Clk), .RN(n106411), .Q(
        n110665) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25382 ), .CK(Clk), .RN(Rst), .Q(n110666)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][27]  ( .D(n104311), 
        .CK(Clk), .RN(Rst), .Q(n110667) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25318 ), .CK(Clk), .RN(Rst), .Q(n110668), 
        .QN(n103290) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25286 ), .CK(Clk), .RN(Rst), .Q(n110669), 
        .QN(n102686) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25254 ), .CK(Clk), .RN(Rst), .Q(n110670), 
        .QN(n102115) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25222 ), .CK(Clk), .RN(Rst), .Q(n110671)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25190 ), .CK(Clk), .RN(Rst), .Q(n74014) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25158 ), .CK(Clk), .RN(Rst), .Q(n110672)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25094 ), .CK(Clk), .RN(Rst), .Q(n110673)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25062 ), .CK(Clk), .RN(Rst), .Q(n74018), 
        .QN(n104611) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25030 ), .CK(Clk), .RN(Rst), .Q(n110674)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24998 ), .CK(Clk), .RN(Rst), .Q(n110675), 
        .QN(n100597) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24966 ), .CK(Clk), .RN(Rst), .Q(n74021) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24934 ), .CK(Clk), .RN(n106476), .Q(n74022) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24902 ), .CK(Clk), .RN(n106476), .Q(
        n110676), .QN(n101153) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24870 ), .CK(Clk), .RN(n106476), .Q(
        n110677) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24838 ), .CK(Clk), .RN(n106476), .Q(
        n110678) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24806 ), .CK(Clk), .RN(n106476), .Q(n74026) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24774 ), .CK(Clk), .RN(n106476), .Q(
        n110679) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][27]  ( .D(n104169), 
        .CK(Clk), .RN(n106476), .Q(n110680) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24678 ), .CK(Clk), .RN(n106476), .Q(
        n110681), .QN(n103286) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24646 ), .CK(Clk), .RN(n106476), .Q(n74031) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24614 ), .CK(Clk), .RN(n106476), .Q(n74032) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24550 ), .CK(Clk), .RN(n106476), .Q(
        n110682) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24518 ), .CK(Clk), .RN(n106432), .Q(
        n110683), .QN(n102679) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24486 ), .CK(Clk), .RN(n106401), .Q(n74036), .QN(n104632) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][27]  ( .D(n104151), 
        .CK(Clk), .RN(Rst), .Q(n110684) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24422 ), .CK(Clk), .RN(Rst), .Q(n110685)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24390 ), .CK(Clk), .RN(n106508), .Q(
        n110686) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24358 ), .CK(Clk), .RN(Rst), .Q(n110687)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24326 ), .CK(Clk), .RN(Rst), .Q(n110688)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24294 ), .CK(Clk), .RN(Rst), .Q(n110689), 
        .QN(n103284) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24262 ), .CK(Clk), .RN(Rst), .Q(n110690)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24166 ), .CK(Clk), .RN(n106433), .Q(
        n110691) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24134 ), .CK(Clk), .RN(Rst), .Q(n110692)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][27]  ( .D(n104078), 
        .CK(Clk), .RN(Rst), .Q(n110693) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24038 ), .CK(Clk), .RN(Rst), .Q(n74050) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24006 ), .CK(Clk), .RN(Rst), .Q(n110694), 
        .QN(n101055) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23974 ), .CK(Clk), .RN(Rst), .Q(n74052) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][27]  ( .D(n104089), 
        .CK(Clk), .RN(Rst), .Q(n110695), .QN(n103843) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23910 ), .CK(Clk), .RN(Rst), .Q(n110696), 
        .QN(n103282) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23878 ), .CK(Clk), .RN(Rst), .Q(n74055) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23814 ), .CK(Clk), .RN(Rst), .Q(n74057) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23782 ), .CK(Clk), .RN(Rst), .Q(n110697), 
        .QN(n101025) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23750 ), .CK(Clk), .RN(n106475), .Q(
        n110698) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23718 ), .CK(Clk), .RN(n106475), .Q(n74060) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23686 ), .CK(Clk), .RN(n106475), .Q(n74061), .QN(n104651) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23654 ), .CK(Clk), .RN(n106475), .Q(n74062) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23622 ), .CK(Clk), .RN(n106475), .Q(
        n110699) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23590 ), .CK(Clk), .RN(n106475), .Q(
        n110700) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23558 ), .CK(Clk), .RN(n106475), .Q(n74065) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23526 ), .CK(Clk), .RN(n106475), .Q(
        n110701) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23494 ), .CK(Clk), .RN(n106475), .Q(n74067) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23462 ), .CK(Clk), .RN(n106475), .Q(n74068) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23430 ), .CK(Clk), .RN(n106475), .Q(n74069) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23398 ), .CK(Clk), .RN(n106474), .Q(
        n110702) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][27]  ( .D(n104063), 
        .CK(Clk), .RN(n106474), .Q(n74071) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23334 ), .CK(Clk), .RN(n106474), .Q(
        n110703) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][27]  ( .D(n104007), 
        .CK(Clk), .RN(n106474), .Q(n110704) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23270 ), .CK(Clk), .RN(n106474), .Q(
        n110705), .QN(n103280) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23238 ), .CK(Clk), .RN(n106474), .Q(
        n110706) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23206 ), .CK(Clk), .RN(n106474), .Q(
        n110707) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23142 ), .CK(Clk), .RN(n106474), .Q(
        n110708) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23110 ), .CK(Clk), .RN(n106474), .Q(
        n110709) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23078 ), .CK(Clk), .RN(n106474), .Q(
        n110710) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23046 ), .CK(Clk), .RN(n106474), .Q(
        n110711) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23014 ), .CK(Clk), .RN(Rst), .Q(n110712)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22982 ), .CK(Clk), .RN(Rst), .Q(n110713)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22950 ), .CK(Clk), .RN(Rst), .Q(n74084) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22918 ), .CK(Clk), .RN(Rst), .Q(n74085) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22886 ), .CK(Clk), .RN(Rst), .Q(n110714)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22854 ), .CK(Clk), .RN(Rst), .Q(n110715)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22822 ), .CK(Clk), .RN(Rst), .Q(n74088) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22790 ), .CK(Clk), .RN(Rst), .Q(n110716)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22758 ), .CK(Clk), .RN(Rst), .Q(n74090) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22726 ), .CK(Clk), .RN(Rst), .Q(n110717)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22694 ), .CK(Clk), .RN(Rst), .Q(n110718)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22662 ), .CK(Clk), .RN(Rst), .Q(n110719)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22630 ), .CK(Clk), .RN(Rst), .Q(n110720)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22598 ), .CK(Clk), .RN(Rst), .Q(n74095) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25894 ), .CK(Clk), .RN(Rst), .Q(n74097) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25926 ), .CK(Clk), .RN(Rst), .Q(n110722)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25958 ), .CK(Clk), .RN(Rst), .Q(n110723)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25990 ), .CK(Clk), .RN(Rst), .Q(n110724), 
        .QN(n103850) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26022 ), .CK(Clk), .RN(Rst), .Q(n110725)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26054 ), .CK(Clk), .RN(Rst), .Q(n110726)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26086 ), .CK(Clk), .RN(Rst), .Q(n110727)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26150 ), .CK(Clk), .RN(Rst), .Q(n110728), 
        .QN(n102119) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][27]  ( .D(n104249), 
        .CK(Clk), .RN(Rst), .Q(n74106) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26214 ), .CK(Clk), .RN(Rst), .Q(n74107) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26246 ), .CK(Clk), .RN(Rst), .Q(n110729)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26278 ), .CK(Clk), .RN(Rst), .Q(n74109) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26310 ), .CK(Clk), .RN(Rst), .Q(n110730)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26342 ), .CK(Clk), .RN(Rst), .Q(n110731)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26374 ), .CK(Clk), .RN(Rst), .Q(n110732)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26406 ), .CK(Clk), .RN(Rst), .Q(n110733)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26438 ), .CK(Clk), .RN(Rst), .Q(n110734)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26470 ), .CK(Clk), .RN(Rst), .Q(n110735)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26502 ), .CK(Clk), .RN(Rst), .Q(n110736), 
        .QN(n103851) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26534 ), .CK(Clk), .RN(Rst), .Q(n110737)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26598 ), .CK(Clk), .RN(n106473), .Q(
        n110739) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26630 ), .CK(Clk), .RN(n106473), .Q(
        n110740) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][27]  ( .D(n106986), 
        .CK(Clk), .RN(n106473), .Q(n110741) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26694 ), .CK(Clk), .RN(n106473), .Q(
        n110742), .QN(n102688) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26726 ), .CK(Clk), .RN(n106473), .Q(
        n110743), .QN(n103293) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26758 ), .CK(Clk), .RN(n106473), .Q(n74124), .QN(n104552) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][27]  ( .D(n107017), 
        .CK(Clk), .RN(n106473), .Q(n110744), .QN(n102120) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26854 ), .CK(Clk), .RN(n106473), .Q(
        n110746), .QN(n103294) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[27]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107089), .Q(
        \DLX_Datapath/next_A_IDEX[27] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[27]  ( .D(n106612), .CK(Clk), .RN(n106473), 
        .Q(n110747) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_log_reg[27]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInA [27]), .Q(
        \DLX_Datapath/ArithLogUnit/A_log [27]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/A_shf_reg[27]  ( .D(
        \DLX_Datapath/MUX_HDU_ALUInA [27]), .GN(n105198), .Q(
        \DLX_Datapath/ArithLogUnit/A_shf [27]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[27]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N140 ), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [27]) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[27]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107055), .Q(
        \DLX_Datapath/next_B_IDEX [27]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[27]  ( .D(n106685), .CK(Clk), .RN(n106473), 
        .Q(n74130), .QN(n104667) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[27]  ( .D(n58869), .CK(Clk), .RN(Rst), .Q(
        n110750) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25860 ), .CK(Clk), .RN(Rst), .Q(n74134) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25828 ), .CK(Clk), .RN(Rst), .Q(n110752)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25796 ), .CK(Clk), .RN(Rst), .Q(n110753)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25764 ), .CK(Clk), .RN(Rst), .Q(n110754)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25700 ), .CK(Clk), .RN(Rst), .Q(n110755)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25636 ), .CK(Clk), .RN(Rst), .Q(n110756)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25604 ), .CK(Clk), .RN(Rst), .Q(n110757)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25572 ), .CK(Clk), .RN(Rst), .Q(n110758)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25540 ), .CK(Clk), .RN(Rst), .Q(n110759)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25508 ), .CK(Clk), .RN(Rst), .Q(n110760), 
        .QN(n100567) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25476 ), .CK(Clk), .RN(n106475), .Q(n74146) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25444 ), .CK(Clk), .RN(Rst), .Q(n110761)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25412 ), .CK(Clk), .RN(n106436), .Q(
        n110762) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25380 ), .CK(Clk), .RN(Rst), .Q(n110763)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25348 ), .CK(Clk), .RN(n106446), .Q(
        n110764) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25316 ), .CK(Clk), .RN(Rst), .Q(n110765), 
        .QN(n103252) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25284 ), .CK(Clk), .RN(n106438), .Q(
        n110766), .QN(n102653) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25252 ), .CK(Clk), .RN(n106395), .Q(
        n110767), .QN(n102087) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25220 ), .CK(Clk), .RN(n106428), .Q(
        n110768) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25188 ), .CK(Clk), .RN(n106420), .Q(n74155) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25156 ), .CK(Clk), .RN(Rst), .Q(n110769)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25092 ), .CK(Clk), .RN(Rst), .Q(n110770)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25060 ), .CK(Clk), .RN(Rst), .Q(n74159), 
        .QN(n104609) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25028 ), .CK(Clk), .RN(Rst), .Q(n110771)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24996 ), .CK(Clk), .RN(Rst), .Q(n110772), 
        .QN(n100599) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][25]  ( .D(n104295), 
        .CK(Clk), .RN(Rst), .Q(n74162) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24932 ), .CK(Clk), .RN(n106475), .Q(n74163) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24900 ), .CK(Clk), .RN(n106373), .Q(
        n110773), .QN(n101155) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24868 ), .CK(Clk), .RN(n106473), .Q(
        n110774) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24836 ), .CK(Clk), .RN(Rst), .Q(n110775)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24804 ), .CK(Clk), .RN(Rst), .Q(n74167) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24772 ), .CK(Clk), .RN(n106439), .Q(
        n110776) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][25]  ( .D(n104168), 
        .CK(Clk), .RN(n106447), .Q(n110777) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24676 ), .CK(Clk), .RN(n106479), .Q(
        n110778), .QN(n103248) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24644 ), .CK(Clk), .RN(n106405), .Q(n74172) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24612 ), .CK(Clk), .RN(n106403), .Q(
        n110779) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24548 ), .CK(Clk), .RN(n106387), .Q(
        n110780) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24516 ), .CK(Clk), .RN(n106384), .Q(
        n110781), .QN(n102646) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24484 ), .CK(Clk), .RN(n106382), .Q(n74177), .QN(n104630) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][25]  ( .D(n104145), 
        .CK(Clk), .RN(n106389), .Q(n110782) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24420 ), .CK(Clk), .RN(Rst), .Q(n110783)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24388 ), .CK(Clk), .RN(n106383), .Q(
        n110784) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24356 ), .CK(Clk), .RN(Rst), .Q(n110785)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24324 ), .CK(Clk), .RN(Rst), .Q(n110786)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24292 ), .CK(Clk), .RN(Rst), .Q(n110787), 
        .QN(n103246) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24260 ), .CK(Clk), .RN(Rst), .Q(n110788)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24228 ), .CK(Clk), .RN(Rst), .Q(n110789)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24164 ), .CK(Clk), .RN(n106502), .Q(
        n110790) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24132 ), .CK(Clk), .RN(Rst), .Q(n110791)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][25]  ( .D(n104077), 
        .CK(Clk), .RN(Rst), .Q(n110792) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24036 ), .CK(Clk), .RN(Rst), .Q(n74191) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24004 ), .CK(Clk), .RN(Rst), .Q(n110793), 
        .QN(n101056) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23972 ), .CK(Clk), .RN(Rst), .Q(n110794)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][25]  ( .D(n104088), 
        .CK(Clk), .RN(Rst), .Q(n110795), .QN(n103812) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23908 ), .CK(Clk), .RN(Rst), .Q(n110796), 
        .QN(n103244) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23876 ), .CK(Clk), .RN(Rst), .Q(n74196) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23812 ), .CK(Clk), .RN(Rst), .Q(n110797)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23780 ), .CK(Clk), .RN(Rst), .Q(n110798), 
        .QN(n101027) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23748 ), .CK(Clk), .RN(Rst), .Q(n110799)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23716 ), .CK(Clk), .RN(Rst), .Q(n74201) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23684 ), .CK(Clk), .RN(Rst), .Q(n110800), 
        .QN(n100997) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23652 ), .CK(Clk), .RN(Rst), .Q(n74203) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23620 ), .CK(Clk), .RN(Rst), .Q(n110801)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23588 ), .CK(Clk), .RN(Rst), .Q(n110802)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23556 ), .CK(Clk), .RN(Rst), .Q(n74206) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23524 ), .CK(Clk), .RN(Rst), .Q(n110803)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23492 ), .CK(Clk), .RN(Rst), .Q(n74208) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23460 ), .CK(Clk), .RN(Rst), .Q(n74209) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23428 ), .CK(Clk), .RN(Rst), .Q(n74210) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23396 ), .CK(Clk), .RN(Rst), .Q(n110804)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23364 ), .CK(Clk), .RN(Rst), .Q(n74212) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23332 ), .CK(Clk), .RN(Rst), .Q(n110805)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][25]  ( .D(n104006), 
        .CK(Clk), .RN(Rst), .Q(n110806) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23268 ), .CK(Clk), .RN(Rst), .Q(n110807), 
        .QN(n103242) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23236 ), .CK(Clk), .RN(Rst), .Q(n110808)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23204 ), .CK(Clk), .RN(Rst), .Q(n110809)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23140 ), .CK(Clk), .RN(Rst), .Q(n110810)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23108 ), .CK(Clk), .RN(Rst), .Q(n110811)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23076 ), .CK(Clk), .RN(Rst), .Q(n110812)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][25]  ( .D(n103992), 
        .CK(Clk), .RN(Rst), .Q(n110813) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23012 ), .CK(Clk), .RN(Rst), .Q(n110814)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22980 ), .CK(Clk), .RN(Rst), .Q(n110815)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22948 ), .CK(Clk), .RN(Rst), .Q(n74225) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22916 ), .CK(Clk), .RN(Rst), .Q(n74226) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22884 ), .CK(Clk), .RN(Rst), .Q(n110816)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22852 ), .CK(Clk), .RN(Rst), .Q(n110817)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22820 ), .CK(Clk), .RN(Rst), .Q(n74229) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22788 ), .CK(Clk), .RN(Rst), .Q(n110818)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22756 ), .CK(Clk), .RN(Rst), .Q(n74231) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22724 ), .CK(Clk), .RN(Rst), .Q(n110819)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22692 ), .CK(Clk), .RN(Rst), .Q(n110820)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22660 ), .CK(Clk), .RN(Rst), .Q(n110821)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22628 ), .CK(Clk), .RN(Rst), .Q(n110822)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22596 ), .CK(Clk), .RN(Rst), .Q(n110823)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25892 ), .CK(Clk), .RN(Rst), .Q(n74238) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25924 ), .CK(Clk), .RN(Rst), .Q(n110825)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25956 ), .CK(Clk), .RN(Rst), .Q(n110826)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25988 ), .CK(Clk), .RN(Rst), .Q(n110827), 
        .QN(n103820) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26020 ), .CK(Clk), .RN(Rst), .Q(n110828)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26052 ), .CK(Clk), .RN(Rst), .Q(n110829)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26084 ), .CK(Clk), .RN(Rst), .Q(n110830)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26148 ), .CK(Clk), .RN(Rst), .Q(n110831), 
        .QN(n102091) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][25]  ( .D(n104250), 
        .CK(Clk), .RN(Rst), .Q(n74247) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26212 ), .CK(Clk), .RN(Rst), .Q(n74248) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26244 ), .CK(Clk), .RN(Rst), .Q(n110832)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26276 ), .CK(Clk), .RN(n106478), .Q(n74250) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26308 ), .CK(Clk), .RN(n106478), .Q(
        n110833) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26340 ), .CK(Clk), .RN(n106478), .Q(
        n110834) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26372 ), .CK(Clk), .RN(n106478), .Q(
        n110835) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26404 ), .CK(Clk), .RN(n106478), .Q(
        n110836) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26436 ), .CK(Clk), .RN(n106478), .Q(
        n110837) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26468 ), .CK(Clk), .RN(n106478), .Q(
        n110838) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26500 ), .CK(Clk), .RN(n106478), .Q(
        n110839), .QN(n103821) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26532 ), .CK(Clk), .RN(n106478), .Q(
        n110840) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26596 ), .CK(Clk), .RN(n106478), .Q(
        n110842) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26628 ), .CK(Clk), .RN(n106478), .Q(
        n110843) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][25]  ( .D(n106984), 
        .CK(Clk), .RN(n106477), .Q(n110844) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26692 ), .CK(Clk), .RN(n106477), .Q(
        n110845), .QN(n102655) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26724 ), .CK(Clk), .RN(n106477), .Q(
        n110846), .QN(n103255) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26756 ), .CK(Clk), .RN(n106477), .Q(n74265), .QN(n104550) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][25]  ( .D(n107015), 
        .CK(Clk), .RN(n106477), .Q(n110847), .QN(n102092) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26852 ), .CK(Clk), .RN(n106477), .Q(
        n110849), .QN(n103256) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[25]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107087), .Q(
        \DLX_Datapath/next_A_IDEX[25] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[25]  ( .D(n106627), .CK(Clk), .RN(n106477), 
        .Q(n110850) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[25]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107053), .Q(
        \DLX_Datapath/next_B_IDEX [25]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[25]  ( .D(n106683), .CK(Clk), .RN(n106477), 
        .Q(n74270), .QN(n104665) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[25]  ( .D(n58867), .CK(Clk), .RN(n106477), 
        .Q(n110851) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[32][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25859 ), .CK(Clk), .RN(Rst), .Q(n74274) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[33][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25827 ), .CK(Clk), .RN(Rst), .Q(n110853)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25795 ), .CK(Clk), .RN(Rst), .Q(n110854)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[35][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25763 ), .CK(Clk), .RN(Rst), .Q(n110855)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[37][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25699 ), .CK(Clk), .RN(Rst), .Q(n110856)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[39][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25635 ), .CK(Clk), .RN(Rst), .Q(n110857)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[40][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25603 ), .CK(Clk), .RN(Rst), .Q(n110858)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[41][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25571 ), .CK(Clk), .RN(Rst), .Q(n110859)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[42][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25539 ), .CK(Clk), .RN(Rst), .Q(n110860)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[43][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25507 ), .CK(Clk), .RN(Rst), .Q(n110861), 
        .QN(n100568) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[44][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25475 ), .CK(Clk), .RN(n106381), .Q(n74286) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[45][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25443 ), .CK(Clk), .RN(n106502), .Q(
        n110862) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[46][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25411 ), .CK(Clk), .RN(Rst), .Q(n110863)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[47][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25379 ), .CK(Clk), .RN(Rst), .Q(n110864)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[48][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25347 ), .CK(Clk), .RN(Rst), .Q(n110865)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25315 ), .CK(Clk), .RN(Rst), .Q(n110866), 
        .QN(n103233) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[50][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25283 ), .CK(Clk), .RN(Rst), .Q(n110867), 
        .QN(n102637) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[51][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25251 ), .CK(Clk), .RN(Rst), .Q(n110868), 
        .QN(n102070) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[52][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25219 ), .CK(Clk), .RN(n106371), .Q(
        n110869) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[53][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25187 ), .CK(Clk), .RN(Rst), .Q(n74295) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[54][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25155 ), .CK(Clk), .RN(n106497), .Q(
        n110870) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[56][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25091 ), .CK(Clk), .RN(n106497), .Q(
        n110871) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[57][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25059 ), .CK(Clk), .RN(n106407), .Q(n74299), .QN(n104608) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[58][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25027 ), .CK(Clk), .RN(Rst), .Q(n110872)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[59][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24995 ), .CK(Clk), .RN(n106429), .Q(
        n110873), .QN(n100600) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[60][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24963 ), .CK(Clk), .RN(Rst), .Q(n74302) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[61][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24931 ), .CK(Clk), .RN(Rst), .Q(n74303) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[62][24]  ( .D(n104204), 
        .CK(Clk), .RN(n106373), .Q(n110874), .QN(n100771) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[63][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24867 ), .CK(Clk), .RN(Rst), .Q(n110875)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[64][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24835 ), .CK(Clk), .RN(n106473), .Q(
        n110876) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[65][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24803 ), .CK(Clk), .RN(Rst), .Q(n74307) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24771 ), .CK(Clk), .RN(Rst), .Q(n110877)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[68][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24707 ), .CK(Clk), .RN(Rst), .Q(n110878)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[69][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24675 ), .CK(Clk), .RN(n106431), .Q(
        n110879), .QN(n103229) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[70][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24643 ), .CK(Clk), .RN(Rst), .Q(n74312) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[71][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24611 ), .CK(Clk), .RN(Rst), .Q(n110880)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24547 ), .CK(Clk), .RN(Rst), .Q(n110881)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[74][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24515 ), .CK(Clk), .RN(Rst), .Q(n110882), 
        .QN(n102630) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[75][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24483 ), .CK(Clk), .RN(Rst), .Q(n74317), 
        .QN(n104629) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[76][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24451 ), .CK(Clk), .RN(Rst), .Q(n110883)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[77][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24419 ), .CK(Clk), .RN(Rst), .Q(n74319) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[78][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24387 ), .CK(Clk), .RN(Rst), .Q(n110884)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[79][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24355 ), .CK(Clk), .RN(Rst), .Q(n110885)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[80][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24323 ), .CK(Clk), .RN(Rst), .Q(n110886)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[81][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24291 ), .CK(Clk), .RN(Rst), .Q(n110887), 
        .QN(n103227) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[82][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24259 ), .CK(Clk), .RN(Rst), .Q(n110888)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24227 ), .CK(Clk), .RN(n106500), .Q(
        n110889) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[85][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24163 ), .CK(Clk), .RN(Rst), .Q(n110890)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[86][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24131 ), .CK(Clk), .RN(Rst), .Q(n110891)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[89][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24035 ), .CK(Clk), .RN(Rst), .Q(n74331) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[90][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24003 ), .CK(Clk), .RN(Rst), .Q(n110892), 
        .QN(n101057) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[91][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23971 ), .CK(Clk), .RN(Rst), .Q(n110893)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[92][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23939 ), .CK(Clk), .RN(n106415), .Q(
        n110894), .QN(n103796) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[93][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23907 ), .CK(Clk), .RN(Rst), .Q(n110895), 
        .QN(n103225) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[94][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23875 ), .CK(Clk), .RN(Rst), .Q(n74336) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[96][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23811 ), .CK(Clk), .RN(n106467), .Q(n74338) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[97][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23779 ), .CK(Clk), .RN(Rst), .Q(n110896), 
        .QN(n101028) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[98][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23747 ), .CK(Clk), .RN(Rst), .Q(n110897)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[99][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23715 ), .CK(Clk), .RN(Rst), .Q(n74341) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[100][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23683 ), .CK(Clk), .RN(Rst), .Q(n74342), 
        .QN(n104650) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[101][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23651 ), .CK(Clk), .RN(Rst), .Q(n74343) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[102][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23619 ), .CK(Clk), .RN(Rst), .Q(n110898)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[103][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23587 ), .CK(Clk), .RN(n106468), .Q(
        n110899) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[105][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23523 ), .CK(Clk), .RN(Rst), .Q(n110900)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[106][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23491 ), .CK(Clk), .RN(n106492), .Q(n74348) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[107][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23459 ), .CK(Clk), .RN(n106394), .Q(n74349) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23427 ), .CK(Clk), .RN(n106372), .Q(
        n110901) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[109][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23395 ), .CK(Clk), .RN(Rst), .Q(n110902)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[110][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23363 ), .CK(Clk), .RN(n106508), .Q(
        n110903) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[111][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23331 ), .CK(Clk), .RN(Rst), .Q(n110904)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23299 ), .CK(Clk), .RN(n106372), .Q(
        n110905) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23267 ), .CK(Clk), .RN(n106488), .Q(
        n110906), .QN(n103223) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[114][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23235 ), .CK(Clk), .RN(n106489), .Q(
        n110907) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[115][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23203 ), .CK(Clk), .RN(n106490), .Q(
        n110908) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23171 ), .CK(Clk), .RN(n106372), .Q(
        n110909) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23139 ), .CK(Clk), .RN(Rst), .Q(n110910)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[118][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23107 ), .CK(Clk), .RN(n106372), .Q(
        n110911) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[119][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23075 ), .CK(Clk), .RN(n106508), .Q(
        n110912) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[120][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23043 ), .CK(Clk), .RN(n106461), .Q(
        n110913) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[121][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23011 ), .CK(Clk), .RN(n106461), .Q(
        n110914) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[122][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22979 ), .CK(Clk), .RN(n106461), .Q(
        n110915) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[123][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22947 ), .CK(Clk), .RN(n106461), .Q(n74365) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[124][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22915 ), .CK(Clk), .RN(n106461), .Q(n74366) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[125][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22883 ), .CK(Clk), .RN(n106461), .Q(
        n110916) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[126][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22851 ), .CK(Clk), .RN(n106461), .Q(
        n110917) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[127][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22819 ), .CK(Clk), .RN(n106461), .Q(
        n110918) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[128][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22787 ), .CK(Clk), .RN(n106461), .Q(
        n110919) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[129][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22755 ), .CK(Clk), .RN(n106461), .Q(n74371) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22723 ), .CK(Clk), .RN(n106461), .Q(
        n110920) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[131][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22691 ), .CK(Clk), .RN(n106461), .Q(
        n110921) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[132][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22659 ), .CK(Clk), .RN(Rst), .Q(n110922)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[133][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22627 ), .CK(Clk), .RN(n106498), .Q(
        n110923) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[134][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22595 ), .CK(Clk), .RN(Rst), .Q(n110924)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25891 ), .CK(Clk), .RN(n106503), .Q(n74378) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[30][24]  ( .D(n104266), 
        .CK(Clk), .RN(n106472), .Q(n110926) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[29][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25955 ), .CK(Clk), .RN(n106502), .Q(
        n110927) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[28][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25987 ), .CK(Clk), .RN(n106501), .Q(
        n110928), .QN(n103804) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[27][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26019 ), .CK(Clk), .RN(n106500), .Q(
        n110929) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[26][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26051 ), .CK(Clk), .RN(n106499), .Q(
        n110930) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[25][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26083 ), .CK(Clk), .RN(Rst), .Q(n110931)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[23][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26147 ), .CK(Clk), .RN(Rst), .Q(n110932), 
        .QN(n102074) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[22][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26179 ), .CK(Clk), .RN(n106422), .Q(n74387) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[21][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26211 ), .CK(Clk), .RN(n106421), .Q(n74388) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[20][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26243 ), .CK(Clk), .RN(n106420), .Q(
        n110933) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[19][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26275 ), .CK(Clk), .RN(n106484), .Q(n74390) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[18][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26307 ), .CK(Clk), .RN(n106419), .Q(
        n110934) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[17][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26339 ), .CK(Clk), .RN(n106418), .Q(
        n110935) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[16][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26371 ), .CK(Clk), .RN(n106394), .Q(
        n110936) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[15][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26403 ), .CK(Clk), .RN(n106478), .Q(
        n110937) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26435 ), .CK(Clk), .RN(n106477), .Q(
        n110938) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[13][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26467 ), .CK(Clk), .RN(n106477), .Q(
        n110939) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[12][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26499 ), .CK(Clk), .RN(Rst), .Q(n110940), 
        .QN(n103805) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[11][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26531 ), .CK(Clk), .RN(Rst), .Q(n110941)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[9][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26595 ), .CK(Clk), .RN(n106428), .Q(
        n110943) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[8][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26627 ), .CK(Clk), .RN(n106427), .Q(
        n110944) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[7][24]  ( .D(n106983), 
        .CK(Clk), .RN(Rst), .Q(n110945) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[6][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26691 ), .CK(Clk), .RN(n106426), .Q(
        n110946), .QN(n102639) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[5][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26723 ), .CK(Clk), .RN(n106425), .Q(
        n110947), .QN(n103236) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[4][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26755 ), .CK(Clk), .RN(n106472), .Q(n74405), .QN(n104549) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[3][24]  ( .D(n107014), 
        .CK(Clk), .RN(Rst), .Q(n110948), .QN(n102075) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[1][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26851 ), .CK(Clk), .RN(n106424), .Q(
        n110950), .QN(n103237) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out1_reg[24]  ( .G(
        \DLX_Datapath/RegisterFile/N46898 ), .D(n107086), .Q(
        \DLX_Datapath/next_A_IDEX[24] ) );
  DFFR_X2 \DLX_Datapath/A_IDEX_reg[24]  ( .D(n106611), .CK(Clk), .RN(Rst), .Q(
        n110951) );
  DLH_X2 \DLX_Datapath/RegisterFile/Out2_reg[24]  ( .G(
        \DLX_Datapath/RegisterFile/N46899 ), .D(n107052), .Q(
        \DLX_Datapath/next_B_IDEX [24]) );
  DFFR_X2 \DLX_Datapath/B_IDEX_reg[24]  ( .D(n106682), .CK(Clk), .RN(Rst), .Q(
        n74410), .QN(n104664) );
  DFFR_X2 \DLX_Datapath/B_EXMEM_reg[24]  ( .D(n58865), .CK(Clk), .RN(Rst), .Q(
        n110952) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[22]  ( .D(n107584), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [22]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[23]  ( .D(n107585), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [23]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[24]  ( .D(n104365), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [24]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[24]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N137 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [24]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[24]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [24]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [24]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[24]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N169 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [24]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[25]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N138 ), .Q(\DLX_Datapath/ArithLogUnit/A_add [25]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[25]  ( .G(n106370), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [25]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [25]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[25]  ( .G(n106368), .D(
        \DLX_Datapath/ArithLogUnit/N170 ), .Q(
        \DLX_Datapath/ArithLogUnit/B_add [25]) );
  DFFR_X2 \DLX_Datapath/PC_reg[25]  ( .D(n60300), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [1]), .QN(n57428) );
  DFFR_X2 \DLX_Datapath/PC_reg[24]  ( .D(n60301), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [0]), .QN(n59477) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[25]  ( .D(n107593), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [25]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[26]  ( .D(n107594), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [26]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[27]  ( .D(n107595), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [27]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[28]  ( .D(n104366), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [28]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[29]  ( .D(n107588), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [29]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/A_add_reg[30]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(n106877), .Q(
        \DLX_Datapath/ArithLogUnit/A_add [30]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_log_reg[30]  ( .G(
        \DLX_Datapath/ArithLogUnit/N178 ), .D(
        \DLX_Datapath/MUX_HDU_ALUInB [30]), .Q(
        \DLX_Datapath/ArithLogUnit/B_log [30]) );
  DLH_X2 \DLX_Datapath/ArithLogUnit/B_add_reg[30]  ( .G(
        \DLX_Datapath/ArithLogUnit/N112 ), .D(\DLX_Datapath/ArithLogUnit/N175 ), .Q(\DLX_Datapath/ArithLogUnit/B_add [30]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[30]  ( .D(n107589), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [30]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/useBorrow_cmp_reg  ( .D(
        \DLX_Datapath/ArithLogUnit/N187 ), .GN(n106359), .Q(
        \DLX_Datapath/ArithLogUnit/useBorrow_cmp ) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Sum_cmp_reg[31]  ( .D(n107590), .GN(
        n106359), .Q(\DLX_Datapath/ArithLogUnit/Sum_cmp [31]) );
  DLL_X2 \DLX_Datapath/ArithLogUnit/Cout_cmp_reg  ( .D(n69975), .GN(n106359), 
        .Q(\DLX_Datapath/ArithLogUnit/Cout_cmp ) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[19]  ( .D(n103940), .CK(Clk), .RN(Rst), 
        .Q(n110958) );
  DFFR_X2 \DLX_Datapath/PC_IFID_reg[2]  ( .D(n60227), .CK(Clk), .RN(Rst), .Q(
        n110959), .QN(n61666) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[1][1]  ( .D(n60163), .CK(
        Clk), .RN(Rst), .Q(n110960) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[9][1]  ( .D(n60179), .CK(
        Clk), .RN(Rst), .Q(n110961) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[17][1]  ( .D(n60195), 
        .CK(Clk), .RN(Rst), .Q(n110962) );
  DFFR_X2 \DLX_Datapath/PC_reg[29]  ( .D(n60296), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0 [1]), .QN(n57429) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[28]  ( .D(n105053), .CK(Clk), .RN(Rst), 
        .Q(n110964) );
  DFFR_X2 \DLX_Datapath/PC_reg[28]  ( .D(n60297), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0 [0]), .QN(n57426) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[29]  ( .D(n103954), .CK(Clk), .RN(Rst), 
        .Q(net2411318) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[30]  ( .D(n103942), .CK(Clk), .RN(Rst), 
        .Q(n110965) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[31]  ( .D(n103947), .CK(Clk), .RN(Rst), 
        .Q(n110966) );
  DFFR_X2 \DLX_Datapath/PC_IFID_reg[1]  ( .D(n60228), .CK(Clk), .RN(Rst), .Q(
        n110967), .QN(n59421) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[5][1]  ( .D(n60171), .CK(
        Clk), .RN(Rst), .Q(n110968) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[13][0]  ( .D(n60188), 
        .CK(Clk), .RN(Rst), .Q(n110969) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[13][1]  ( .D(n60187), 
        .CK(Clk), .RN(Rst), .Q(n110970) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[21][0]  ( .D(n60204), 
        .CK(Clk), .RN(Rst), .Q(n110971) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[21][1]  ( .D(n60203), 
        .CK(Clk), .RN(Rst), .Q(n110972) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[29][1]  ( .D(n60219), 
        .CK(Clk), .RN(Rst), .Q(n110973) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[4][0]  ( .D(n60170), .CK(
        Clk), .RN(Rst), .Q(n110974) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[4][1]  ( .D(n60169), .CK(
        Clk), .RN(Rst), .Q(n110975) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[12][0]  ( .D(n60186), 
        .CK(Clk), .RN(Rst), .Q(n110976) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[12][1]  ( .D(n60185), 
        .CK(Clk), .RN(Rst), .Q(n110977) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[20][0]  ( .D(n60202), 
        .CK(Clk), .RN(Rst), .Q(n110978) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[20][1]  ( .D(n60201), 
        .CK(Clk), .RN(Rst), .Q(n110979) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[28][1]  ( .D(n60217), 
        .CK(Clk), .RN(Rst), .Q(n110980) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[0][0]  ( .D(n60162), .CK(
        Clk), .RN(Rst), .Q(n110981) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[0][1]  ( .D(n60161), .CK(
        Clk), .RN(Rst), .Q(n110982) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[8][0]  ( .D(n60178), .CK(
        Clk), .RN(Rst), .Q(n110983) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[8][1]  ( .D(n60177), .CK(
        Clk), .RN(n106460), .Q(n110984) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[16][0]  ( .D(n60194), 
        .CK(Clk), .RN(n106460), .Q(n110985) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[16][1]  ( .D(n60193), 
        .CK(Clk), .RN(n106460), .Q(n110986) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[24][0]  ( .D(n60210), 
        .CK(Clk), .RN(n106460), .Q(n110987) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[24][1]  ( .D(n60209), 
        .CK(Clk), .RN(n106460), .Q(n110988) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[7][0]  ( .D(n60176), .CK(
        Clk), .RN(n106460), .Q(n110989) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[7][1]  ( .D(n60175), .CK(
        Clk), .RN(n106460), .Q(n110990) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[15][0]  ( .D(n60192), 
        .CK(Clk), .RN(n106460), .Q(n110991) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[15][1]  ( .D(n60191), 
        .CK(Clk), .RN(n106460), .Q(n110992) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[23][0]  ( .D(n60208), 
        .CK(Clk), .RN(n106460), .Q(n110993) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[23][1]  ( .D(n60207), 
        .CK(Clk), .RN(n106460), .Q(n110994) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[31][1]  ( .D(n60223), 
        .CK(Clk), .RN(n106460), .Q(n110995) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[6][1]  ( .D(n60173), .CK(
        Clk), .RN(n106407), .Q(n110996) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[14][0]  ( .D(n60190), 
        .CK(Clk), .RN(n106390), .Q(n110997) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[14][1]  ( .D(n60189), 
        .CK(Clk), .RN(n106497), .Q(n110998) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[22][0]  ( .D(n60206), 
        .CK(Clk), .RN(Rst), .Q(n110999) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[22][1]  ( .D(n60205), 
        .CK(Clk), .RN(Rst), .Q(n111000) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[30][1]  ( .D(n60221), 
        .CK(Clk), .RN(Rst), .Q(n111001) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[3][1]  ( .D(n60167), .CK(
        Clk), .RN(Rst), .Q(n111002) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[11][0]  ( .D(n60184), 
        .CK(Clk), .RN(Rst), .Q(n111003) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[11][1]  ( .D(n60183), 
        .CK(Clk), .RN(Rst), .Q(n111004) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[19][0]  ( .D(n60200), 
        .CK(Clk), .RN(Rst), .Q(n111005) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[19][1]  ( .D(n60199), 
        .CK(Clk), .RN(Rst), .Q(n111006) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[27][0]  ( .D(n60216), 
        .CK(Clk), .RN(n106472), .Q(n111007) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[27][1]  ( .D(n60215), 
        .CK(Clk), .RN(n106472), .Q(n111008) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[2][1]  ( .D(n60165), .CK(
        Clk), .RN(n106472), .Q(n111009) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[10][0]  ( .D(n60182), 
        .CK(Clk), .RN(n106472), .Q(n111010) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[10][1]  ( .D(n60181), 
        .CK(Clk), .RN(n106472), .Q(n111011) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[18][0]  ( .D(n60198), 
        .CK(Clk), .RN(n106472), .Q(n111012) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[18][1]  ( .D(n60197), 
        .CK(Clk), .RN(n106472), .Q(n111013) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[26][0]  ( .D(n60214), 
        .CK(Clk), .RN(n106472), .Q(n111014) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[26][1]  ( .D(n60213), 
        .CK(Clk), .RN(n106472), .Q(n111015) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[127]  ( .A(n58864), .EN(
        n106365), .Z(stackBus_Out[127]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[126]  ( .A(n58863), .EN(
        n58746), .Z(stackBus_Out[126]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[125]  ( .A(n58862), .EN(
        n106367), .Z(stackBus_Out[125]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[124]  ( .A(n58861), .EN(
        n106361), .Z(stackBus_Out[124]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[123]  ( .A(n58860), .EN(
        n106364), .Z(stackBus_Out[123]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[122]  ( .A(n58859), .EN(
        n106366), .Z(stackBus_Out[122]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[121]  ( .A(n58858), .EN(
        n106365), .Z(stackBus_Out[121]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[120]  ( .A(n58857), .EN(
        n106362), .Z(stackBus_Out[120]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[119]  ( .A(n58856), .EN(
        n58746), .Z(stackBus_Out[119]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[118]  ( .A(n58855), .EN(
        n106364), .Z(stackBus_Out[118]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[117]  ( .A(n58854), .EN(
        n106362), .Z(stackBus_Out[117]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[116]  ( .A(n58853), .EN(
        n106365), .Z(stackBus_Out[116]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[115]  ( .A(n58852), .EN(
        n58746), .Z(stackBus_Out[115]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[114]  ( .A(n58851), .EN(
        n106367), .Z(stackBus_Out[114]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[113]  ( .A(n58850), .EN(
        n106364), .Z(stackBus_Out[113]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[112]  ( .A(n58849), .EN(
        n106364), .Z(stackBus_Out[112]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[111]  ( .A(n58848), .EN(
        n106365), .Z(stackBus_Out[111]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[110]  ( .A(n58847), .EN(
        n106365), .Z(stackBus_Out[110]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[109]  ( .A(n58846), .EN(
        n106367), .Z(stackBus_Out[109]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[108]  ( .A(n58845), .EN(
        n106364), .Z(stackBus_Out[108]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[107]  ( .A(n58844), .EN(
        n106367), .Z(stackBus_Out[107]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[106]  ( .A(n58843), .EN(
        n106365), .Z(stackBus_Out[106]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[105]  ( .A(n58842), .EN(
        n106366), .Z(stackBus_Out[105]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[104]  ( .A(n58841), .EN(
        n106367), .Z(stackBus_Out[104]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[103]  ( .A(n58840), .EN(
        n106364), .Z(stackBus_Out[103]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[102]  ( .A(n58839), .EN(
        n106364), .Z(stackBus_Out[102]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[101]  ( .A(n58838), .EN(
        n106363), .Z(stackBus_Out[101]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[100]  ( .A(n58837), .EN(
        n106366), .Z(stackBus_Out[100]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[99]  ( .A(n58836), .EN(
        n106361), .Z(stackBus_Out[99]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[98]  ( .A(n58835), .EN(
        n58746), .Z(stackBus_Out[98]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[97]  ( .A(n58834), .EN(
        n106362), .Z(stackBus_Out[97]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[96]  ( .A(n58833), .EN(
        n106361), .Z(stackBus_Out[96]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[95]  ( .A(n106732), .EN(
        n106363), .Z(stackBus_Out[95]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[94]  ( .A(n106731), .EN(
        n106362), .Z(stackBus_Out[94]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[93]  ( .A(n106730), .EN(
        n106364), .Z(stackBus_Out[93]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[92]  ( .A(n106729), .EN(
        n106361), .Z(stackBus_Out[92]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[91]  ( .A(n106728), .EN(
        n106366), .Z(stackBus_Out[91]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[90]  ( .A(n106727), .EN(
        n58746), .Z(stackBus_Out[90]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[89]  ( .A(n106726), .EN(
        n106361), .Z(stackBus_Out[89]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[88]  ( .A(n106725), .EN(
        n106364), .Z(stackBus_Out[88]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[87]  ( .A(n106724), .EN(
        n106362), .Z(stackBus_Out[87]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[86]  ( .A(n106723), .EN(
        n106366), .Z(stackBus_Out[86]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[85]  ( .A(n106722), .EN(
        n106361), .Z(stackBus_Out[85]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[84]  ( .A(n106721), .EN(
        n106362), .Z(stackBus_Out[84]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[83]  ( .A(n106720), .EN(
        n106362), .Z(stackBus_Out[83]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[82]  ( .A(n106719), .EN(
        n106365), .Z(stackBus_Out[82]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[81]  ( .A(n106718), .EN(
        n106365), .Z(stackBus_Out[81]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[80]  ( .A(n106717), .EN(
        n106366), .Z(stackBus_Out[80]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[79]  ( .A(n106716), .EN(
        n58746), .Z(stackBus_Out[79]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[78]  ( .A(n106715), .EN(
        n106361), .Z(stackBus_Out[78]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[77]  ( .A(n106714), .EN(
        n106362), .Z(stackBus_Out[77]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[76]  ( .A(n106713), .EN(
        n106367), .Z(stackBus_Out[76]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[75]  ( .A(n106712), .EN(
        n106363), .Z(stackBus_Out[75]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[74]  ( .A(n106711), .EN(
        n106365), .Z(stackBus_Out[74]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[73]  ( .A(n106710), .EN(
        n106361), .Z(stackBus_Out[73]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[72]  ( .A(n106709), .EN(
        n106364), .Z(stackBus_Out[72]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[71]  ( .A(n106708), .EN(
        n106367), .Z(stackBus_Out[71]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[70]  ( .A(n106707), .EN(
        n106366), .Z(stackBus_Out[70]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[69]  ( .A(n106706), .EN(
        n106363), .Z(stackBus_Out[69]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[68]  ( .A(n106705), .EN(
        n106365), .Z(stackBus_Out[68]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[67]  ( .A(n106704), .EN(
        n106364), .Z(stackBus_Out[67]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[66]  ( .A(n106703), .EN(
        n106366), .Z(stackBus_Out[66]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[65]  ( .A(n106702), .EN(
        n106361), .Z(stackBus_Out[65]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[64]  ( .A(n106701), .EN(
        n106361), .Z(stackBus_Out[64]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[63]  ( .A(n58800), .EN(
        n106361), .Z(stackBus_Out[63]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[62]  ( .A(n58799), .EN(
        n106365), .Z(stackBus_Out[62]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[61]  ( .A(n58798), .EN(
        n106362), .Z(stackBus_Out[61]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[60]  ( .A(n58797), .EN(
        n106362), .Z(stackBus_Out[60]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[59]  ( .A(n58796), .EN(
        n106362), .Z(stackBus_Out[59]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[58]  ( .A(n58795), .EN(
        n106367), .Z(stackBus_Out[58]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[57]  ( .A(n58794), .EN(
        n106363), .Z(stackBus_Out[57]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[56]  ( .A(n58793), .EN(
        n106365), .Z(stackBus_Out[56]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[55]  ( .A(n58792), .EN(
        n106365), .Z(stackBus_Out[55]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[54]  ( .A(n58791), .EN(
        n106364), .Z(stackBus_Out[54]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[53]  ( .A(n58790), .EN(
        n106366), .Z(stackBus_Out[53]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[52]  ( .A(n58789), .EN(
        n106367), .Z(stackBus_Out[52]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[51]  ( .A(n58788), .EN(
        n106367), .Z(stackBus_Out[51]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[50]  ( .A(n58787), .EN(
        n106366), .Z(stackBus_Out[50]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[49]  ( .A(n58786), .EN(
        n106363), .Z(stackBus_Out[49]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[48]  ( .A(n58785), .EN(
        n106362), .Z(stackBus_Out[48]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[47]  ( .A(n58784), .EN(
        n106367), .Z(stackBus_Out[47]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[46]  ( .A(n58783), .EN(
        n106366), .Z(stackBus_Out[46]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[45]  ( .A(n58782), .EN(
        n106361), .Z(stackBus_Out[45]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[44]  ( .A(n58781), .EN(
        n106363), .Z(stackBus_Out[44]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[43]  ( .A(n58780), .EN(
        n106363), .Z(stackBus_Out[43]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[42]  ( .A(n58779), .EN(
        n106365), .Z(stackBus_Out[42]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[41]  ( .A(n58778), .EN(
        n106363), .Z(stackBus_Out[41]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[40]  ( .A(n58777), .EN(
        n106365), .Z(stackBus_Out[40]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[39]  ( .A(n58776), .EN(
        n106366), .Z(stackBus_Out[39]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[38]  ( .A(n58775), .EN(
        n106363), .Z(stackBus_Out[38]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[37]  ( .A(n58774), .EN(
        n106362), .Z(stackBus_Out[37]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[36]  ( .A(n58773), .EN(
        n106363), .Z(stackBus_Out[36]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[35]  ( .A(n58772), .EN(
        n106366), .Z(stackBus_Out[35]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[34]  ( .A(n58771), .EN(
        n106363), .Z(stackBus_Out[34]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[33]  ( .A(n58770), .EN(
        n106366), .Z(stackBus_Out[33]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[32]  ( .A(n58769), .EN(
        n106363), .Z(stackBus_Out[32]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[31]  ( .A(n103969), .EN(
        n58746), .Z(stackBus_Out[31]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[30]  ( .A(n103970), .EN(
        n106363), .Z(stackBus_Out[30]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[29]  ( .A(n103971), .EN(
        n106363), .Z(stackBus_Out[29]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[28]  ( .A(n103972), .EN(
        n106365), .Z(stackBus_Out[28]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[27]  ( .A(n103973), .EN(
        n106363), .Z(stackBus_Out[27]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[26]  ( .A(n103974), .EN(
        n106362), .Z(stackBus_Out[26]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[25]  ( .A(n103975), .EN(
        n106363), .Z(stackBus_Out[25]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[24]  ( .A(n103976), .EN(
        n106363), .Z(stackBus_Out[24]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[23]  ( .A(n103977), .EN(
        n106364), .Z(stackBus_Out[23]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[22]  ( .A(n103978), .EN(
        n106365), .Z(stackBus_Out[22]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[21]  ( .A(n103979), .EN(
        n106364), .Z(stackBus_Out[21]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[20]  ( .A(n103980), .EN(
        n106366), .Z(stackBus_Out[20]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[19]  ( .A(n103981), .EN(
        n106361), .Z(stackBus_Out[19]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[18]  ( .A(n103982), .EN(
        n106367), .Z(stackBus_Out[18]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[17]  ( .A(n103983), .EN(
        n106362), .Z(stackBus_Out[17]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[16]  ( .A(n103984), .EN(
        n106361), .Z(stackBus_Out[16]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[15]  ( .A(n103985), .EN(
        n106364), .Z(stackBus_Out[15]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[14]  ( .A(n103986), .EN(
        n106364), .Z(stackBus_Out[14]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[13]  ( .A(n103987), .EN(
        n106367), .Z(stackBus_Out[13]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[12]  ( .A(n103988), .EN(
        n106367), .Z(stackBus_Out[12]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[11]  ( .A(n103957), .EN(
        n106367), .Z(stackBus_Out[11]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[10]  ( .A(n103958), .EN(
        n106367), .Z(stackBus_Out[10]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[9]  ( .A(n103959), .EN(
        n106364), .Z(stackBus_Out[9]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[8]  ( .A(n103960), .EN(
        n106362), .Z(stackBus_Out[8]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[7]  ( .A(n103961), .EN(
        n106366), .Z(stackBus_Out[7]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[6]  ( .A(n103962), .EN(
        n106366), .Z(stackBus_Out[6]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[5]  ( .A(n103963), .EN(
        n106361), .Z(stackBus_Out[5]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[4]  ( .A(n103964), .EN(
        n106362), .Z(stackBus_Out[4]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[3]  ( .A(n103965), .EN(
        n106364), .Z(stackBus_Out[3]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[2]  ( .A(n103966), .EN(
        n58746), .Z(stackBus_Out[2]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[1]  ( .A(n103967), .EN(
        n106366), .Z(stackBus_Out[1]) );
  TBUF_X4 \DLX_Datapath/RegisterFile/memBus_out_tri[0]  ( .A(n103968), .EN(
        n106367), .Z(stackBus_Out[0]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [29]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [29]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [30]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [30]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [31]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [31]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_0/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [29]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [29]), .CI(n104369), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_0/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [30]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [30]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_0/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [31]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [31]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [25]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [25]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [26]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [26]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [27]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [27]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_0/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [25]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [25]), .CI(n104376), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_0/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [26]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [26]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_0/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [27]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [27]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [21]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [21]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [22]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [22]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [23]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [23]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_0/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [21]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [21]), .CI(n104375), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_0/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [22]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [22]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_0/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [23]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [23]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [17]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [17]), .CI(n109894), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [18]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [18]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [19]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [19]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [17]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [17]), .CI(n104374), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [18]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [18]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [19]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [19]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [13]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [13]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [14]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [14]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [15]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [15]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [13]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [13]), .CI(n104373), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [14]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [14]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [15]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [15]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [9]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [9]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [10]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [10]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [11]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [11]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [9]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [9]), .CI(n104372), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [10]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [10]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [11]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [11]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [5]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [5]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [6]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [6]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [7]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [7]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [5]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [5]), .CI(n104370), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [6]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [6]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [7]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [7]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [1]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [1]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [2]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [2]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [3]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [3]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/U1_1  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [1]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [1]), .CI(n104367), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/U1_2  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [2]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [2]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/U1_3  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_add [3]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [3]), .CI(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/U1_1  ( 
        .A(n111131), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [1]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/S_1[1] ) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/U1_1  ( 
        .A(n111131), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [1]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/S_0[1] ) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/U1_1  ( 
        .A(IR_in[13]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [1]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/U1_2  ( 
        .A(IR_in[14]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [2]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/U1_3  ( 
        .A(IR_in[15]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [3]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/U1_1  ( 
        .A(IR_in[13]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [1]), 
        .CI(n104368), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/U1_2  ( 
        .A(IR_in[14]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [2]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/U1_3  ( 
        .A(IR_in[15]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [3]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/U1_1  ( 
        .A(IR_in[9]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [1]), 
        .CI(net68723), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/U1_2  ( 
        .A(IR_in[10]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [2]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/U1_3  ( 
        .A(IR_in[11]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [3]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/U1_1  ( 
        .A(IR_in[9]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [1]), 
        .CI(net68722), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/U1_2  ( 
        .A(IR_in[10]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [2]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/U1_3  ( 
        .A(IR_in[11]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [3]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/U1_1  ( 
        .A(IR_in[5]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [1]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[1] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[2] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_1 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/U1_2  ( 
        .A(IR_in[6]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [2]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_1 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/U1_3  ( 
        .A(IR_in[7]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [3]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_1 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/U1_1  ( 
        .A(IR_in[5]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [1]), 
        .CI(n104371), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/U1_2  ( 
        .A(IR_in[6]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [2]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/U1_3  ( 
        .A(IR_in[7]), .B(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [3]), 
        .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_0 [3]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/U1_1  ( 
        .A(IR_in[1]), .B(PC_out[1]), .CI(n104326), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[2] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 [1]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/U1_2  ( 
        .A(IR_in[2]), .B(n74605), .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[2] ), .CO(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 [2]) );
  FA_X1 \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/U1_3  ( 
        .A(IR_in[3]), .B(PC_out[3]), .CI(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/RCA_0/add_38_2/carry[3] ), .S(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 [3]) );
  FA_X1 \add_0_root_r2411/U1_5  ( .A(\DLX_Datapath/RegisterFile/old_CWP2[1] ), 
        .B(n104757), .CI(n105034), .CO(\add_0_root_r2411/carry[6] ), .S(
        \DLX_Datapath/RegisterFile/N46177 ) );
  FA_X1 \add_0_root_r2411/U1_6  ( .A(\DLX_Datapath/RegisterFile/old_CWP2[2] ), 
        .B(n104757), .CI(\add_0_root_r2411/carry[6] ), .CO(
        \add_0_root_r2411/carry[7] ), .S(\DLX_Datapath/RegisterFile/N46178 )
         );
  FA_X1 \add_0_root_sub_0_root_DLX_Datapath/RegisterFile/add_172/U1_5  ( .A(
        \DLX_Datapath/RegisterFile/old_CWP2[1] ), .B(n104757), .CI(n62664), 
        .CO(\add_0_root_sub_0_root_DLX_Datapath/RegisterFile/add_172/carry[6] ), .S(\DLX_Datapath/RegisterFile/N9337 ) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[14]  ( .D(n64127), .CK(Clk), .RN(n106472), 
        .Q(\DLX_Datapath/HazardDetUnit/N112 ), .QN(n62574) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[15]  ( .D(n64126), .CK(Clk), .RN(n106472), 
        .Q(\DLX_Datapath/IR_IDEX[15] ), .QN(n62573) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24067 ), .CK(Clk), .RN(n106472), .Q(
        n111016) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[88][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24066 ), .CK(Clk), .RN(n106471), .Q(
        n111017) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25792 ), .CK(Clk), .RN(n106471), .Q(
        n111018) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25791 ), .CK(Clk), .RN(n106471), .Q(
        n111019) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25793 ), .CK(Clk), .RN(n106471), .Q(
        n111020) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[34][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25789 ), .CK(Clk), .RN(n106471), .Q(
        n111021) );
  DFFS_X2 \DLX_Datapath/IR_EXMEM_reg[30]  ( .D(n69315), .CK(Clk), .SN(Rst), 
        .Q(n111022), .QN(n57379) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[13]  ( .D(
        \DLX_Datapath/HazardDetUnit/N111 ), .CK(Clk), .RN(n106470), .Q(
        \DLX_Datapath/HazardDetUnit/N139 ), .QN(n100419) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[12]  ( .D(
        \DLX_Datapath/HazardDetUnit/N110 ), .CK(Clk), .RN(n106470), .Q(
        \DLX_Datapath/HazardDetUnit/N138 ), .QN(n100420) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[11]  ( .D(
        \DLX_Datapath/HazardDetUnit/N109 ), .CK(Clk), .RN(n106470), .Q(
        \DLX_Datapath/HazardDetUnit/N137 ), .QN(n100418) );
  DFFR_X2 \DLX_Datapath/RegisterFile/old_CWP2_reg[0]  ( .D(
        \DLX_Datapath/RegisterFile/old_CWP1 [0]), .CK(Clk), .RN(n106470), .QN(
        n100801) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[16]  ( .D(
        \DLX_Datapath/HazardDetUnit/N95 ), .CK(Clk), .RN(n106470), .Q(
        \DLX_Datapath/HazardDetUnit/N123 ), .QN(n100796) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[18]  ( .D(
        \DLX_Datapath/HazardDetUnit/N97 ), .CK(Clk), .RN(n106470), .Q(
        \DLX_Datapath/HazardDetUnit/N125 ), .QN(n100422) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[17]  ( .D(
        \DLX_Datapath/HazardDetUnit/N96 ), .CK(Clk), .RN(n106470), .Q(
        \DLX_Datapath/HazardDetUnit/N124 ), .QN(n100423) );
  DFFR_X2 \DLX_Datapath/RegisterFile/to_transfer_reg[0]  ( .D(
        \DLX_Datapath/RegisterFile/next_to_transfer [0]), .CK(Clk), .RN(
        n106469), .Q(n104582), .QN(n62190) );
  DFFR_X2 \DLX_Datapath/RegisterFile/to_transfer_reg[1]  ( .D(
        \DLX_Datapath/RegisterFile/next_to_transfer [1]), .CK(Clk), .RN(
        n106469), .Q(n111027), .QN(n62212) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[25]  ( .D(\DLX_Datapath/N352 ), .CK(Clk), 
        .RN(n106469), .Q(n111028), .QN(n61799) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[24]  ( .D(\DLX_Datapath/N351 ), .CK(Clk), 
        .RN(n106469), .Q(n104441), .QN(n100893) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[23]  ( .D(\DLX_Datapath/N350 ), .CK(Clk), 
        .RN(n106469), .QN(n100429) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[22]  ( .D(\DLX_Datapath/N349 ), .CK(Clk), 
        .RN(n106469), .QN(n100430) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[21]  ( .D(\DLX_Datapath/N348 ), .CK(Clk), 
        .RN(n106469), .QN(n100428) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[17]  ( .D(\DLX_Datapath/N344 ), .CK(Clk), 
        .RN(n106469), .Q(\DLX_Datapath/HazardDetUnit/N96 ), .QN(n100719) );
  DFFR_X2 \DLX_Datapath/IR_IDEX_reg[18]  ( .D(\DLX_Datapath/N345 ), .CK(Clk), 
        .RN(n106468), .Q(\DLX_Datapath/HazardDetUnit/N97 ), .QN(n100427) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[0]  ( .D(n106556), .CK(Clk), .RN(n106468), 
        .Q(\DLX_ControlUnit/cw2 [0]) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[15]  ( .D(n106557), .CK(Clk), .RN(n106467), 
        .Q(\DLX_ControlUnit/cw2 [15]) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[13]  ( .D(n106582), .CK(Clk), .RN(n106467), 
        .Q(\DLX_ControlUnit/cw2 [13]) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[8]  ( .D(n103927), .CK(Clk), .RN(n106467), 
        .QN(n100779) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[10]  ( .D(n106560), .CK(Clk), .RN(n106467), 
        .Q(\DLX_ControlUnit/cw2 [10]) );
  DFFR_X2 \DLX_ControlUnit/ALUop2_reg[1]  ( .D(n60328), .CK(Clk), .RN(n106467), 
        .Q(n111033), .QN(n100784) );
  DFFR_X2 \DLX_ControlUnit/ALUop2_reg[0]  ( .D(n60329), .CK(Clk), .RN(n106467), 
        .Q(n111034), .QN(n100795) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23421 ), .CK(Clk), .RN(n106467), .Q(
        n111035) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23554 ), .CK(Clk), .RN(n106467), .Q(
        n111036), .QN(n103776) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[104][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23555 ), .CK(Clk), .RN(n106466), .Q(
        n111037), .QN(n103793) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23423 ), .CK(Clk), .RN(n106466), .Q(
        n111038) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23425 ), .CK(Clk), .RN(n106466), .Q(
        n111039) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[108][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23422 ), .CK(Clk), .RN(n106466), .Q(
        n111040) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[6][0]  ( .D(n60174), .CK(
        Clk), .RN(n106466), .Q(n111041) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[5][0]  ( .D(n60172), .CK(
        Clk), .RN(n106466), .Q(n111042) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[3][0]  ( .D(n60168), .CK(
        Clk), .RN(n106466), .Q(n111043) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[2][0]  ( .D(n60166), .CK(
        Clk), .RN(n106466), .Q(n111044) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[31][0]  ( .D(n60224), 
        .CK(Clk), .RN(n106466), .Q(n111045) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[30][0]  ( .D(n60222), 
        .CK(Clk), .RN(n106466), .Q(n111046) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[29][0]  ( .D(n60220), 
        .CK(Clk), .RN(n106466), .Q(n111047) );
  DFFR_X2 \DLX_Datapath/BrancJump_logic/pred_mem_reg[28][0]  ( .D(n60218), 
        .CK(Clk), .RN(n106466), .Q(n111048) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[22]  ( .D(n58886), .CK(Clk), .RN(Rst), 
        .Q(n111066), .QN(n100667) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[21]  ( .D(n58881), .CK(Clk), .RN(Rst), 
        .Q(n111067), .QN(n100669) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[20]  ( .D(n58876), .CK(Clk), .RN(Rst), 
        .Q(n111068), .QN(n100671) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[31]  ( .D(n58996), .CK(Clk), .RN(Rst), 
        .Q(n111069), .QN(n100649) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[29]  ( .D(n59054), .CK(Clk), .RN(Rst), 
        .Q(n111070), .QN(n100653) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[23]  ( .D(n58888), .CK(Clk), .RN(Rst), 
        .Q(n111071), .QN(n100665) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[19]  ( .D(n58907), .CK(Clk), .RN(Rst), 
        .Q(n111072), .QN(n100673) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[18]  ( .D(n58905), .CK(Clk), .RN(Rst), 
        .Q(n111073), .QN(n100675) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[16]  ( .D(n58899), .CK(Clk), .RN(Rst), 
        .Q(n111074), .QN(n100679) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[9]  ( .D(n58920), .CK(Clk), .RN(Rst), 
        .Q(n111075), .QN(n100693) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[8]  ( .D(n58915), .CK(Clk), .RN(Rst), 
        .Q(n111076), .QN(n100695) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[5]  ( .D(n58925), .CK(Clk), .RN(Rst), 
        .Q(n111077), .QN(n100701) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[17]  ( .D(n58903), .CK(Clk), .RN(
        n106464), .Q(n111078), .QN(n100677) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[14]  ( .D(n58972), .CK(Clk), .RN(
        n106464), .Q(n111079), .QN(n100683) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[13]  ( .D(n58964), .CK(Clk), .RN(
        n106464), .Q(n111080), .QN(n100685) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[11]  ( .D(n58961), .CK(Clk), .RN(
        n106464), .Q(n111081), .QN(n100689) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[10]  ( .D(n58959), .CK(Clk), .RN(
        n106464), .Q(n111082), .QN(n100691) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[6]  ( .D(n58935), .CK(Clk), .RN(
        n106464), .Q(n111083), .QN(n100699) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[3]  ( .D(n58955), .CK(Clk), .RN(
        n106464), .Q(n111084), .QN(n100705) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[2]  ( .D(n58943), .CK(Clk), .RN(
        n106464), .Q(n111085), .QN(n100707) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[1]  ( .D(n58946), .CK(Clk), .RN(
        n106464), .Q(n111086), .QN(n100709) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[0]  ( .D(n59053), .CK(Clk), .RN(
        n106464), .Q(n111087), .QN(n100711) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[7]  ( .D(n58940), .CK(Clk), .RN(
        n106464), .Q(n111088), .QN(n100697) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[4]  ( .D(n58929), .CK(Clk), .RN(
        n106464), .Q(n111089), .QN(n100703) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[30]  ( .D(n58993), .CK(Clk), .RN(
        n106463), .Q(n111090), .QN(n100651) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[28]  ( .D(n58999), .CK(Clk), .RN(
        n106463), .Q(n111091), .QN(n100655) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[27]  ( .D(n58990), .CK(Clk), .RN(
        n106463), .Q(n111092), .QN(n100657) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[26]  ( .D(n58988), .CK(Clk), .RN(
        n106463), .Q(n111093), .QN(n100659) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[25]  ( .D(n58981), .CK(Clk), .RN(
        n106463), .Q(n111094), .QN(n100661) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[24]  ( .D(n58979), .CK(Clk), .RN(
        n106463), .Q(n111095), .QN(n100663) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[15]  ( .D(n58977), .CK(Clk), .RN(
        n106463), .Q(n111096), .QN(n100681) );
  DFFR_X2 \DLX_Datapath/ALUOut_MEMWB_reg[12]  ( .D(n59006), .CK(Clk), .RN(
        n106463), .Q(n111097), .QN(n100687) );
  DFFR_X2 \DLX_Datapath/IR_EXMEM_reg[31]  ( .D(\DLX_Datapath/IR_IDEX[31] ), 
        .CK(Clk), .RN(Rst), .Q(\DLX_Datapath/IR_EXMEM[31] ), .QN(n59326) );
  OAI21_X1 U64741 ( .B1(n62189), .B2(n58698), .A(n79652), .ZN(n104329) );
  NAND2_X1 U64742 ( .A1(n62189), .A2(\DLX_Datapath/next_ALUOut_EXMEM [12]), 
        .ZN(n79652) );
  OAI21_X1 U64743 ( .B1(n62189), .B2(n58691), .A(n79653), .ZN(n104330) );
  NAND2_X1 U64744 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [28]), .A2(n62189), 
        .ZN(n79653) );
  OAI21_X1 U64745 ( .B1(n62189), .B2(n58688), .A(n79654), .ZN(n104331) );
  NAND2_X1 U64746 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [31]), .A2(n62189), 
        .ZN(n79654) );
  OAI21_X1 U64747 ( .B1(n62189), .B2(n58685), .A(n79655), .ZN(n104332) );
  NAND2_X1 U64748 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [30]), .A2(n62189), 
        .ZN(n79655) );
  OAI21_X1 U64749 ( .B1(n62189), .B2(n58682), .A(n79656), .ZN(n104333) );
  NAND2_X1 U64750 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [27]), .A2(n62189), 
        .ZN(n79656) );
  OAI21_X1 U64751 ( .B1(n62189), .B2(n58680), .A(n79657), .ZN(n104334) );
  NAND2_X1 U64752 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [26]), .A2(n62189), 
        .ZN(n79657) );
  OAI21_X1 U64753 ( .B1(n62189), .B2(n58673), .A(n79658), .ZN(n104335) );
  NAND2_X1 U64754 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [25]), .A2(n62189), 
        .ZN(n79658) );
  OAI21_X1 U64755 ( .B1(n62189), .B2(n58671), .A(n79659), .ZN(n104336) );
  NAND2_X1 U64756 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [24]), .A2(n106358), 
        .ZN(n79659) );
  OAI21_X1 U64757 ( .B1(n62189), .B2(n58669), .A(n79660), .ZN(n104337) );
  NAND2_X1 U64758 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [15]), .A2(n62189), 
        .ZN(n79660) );
  OAI21_X1 U64759 ( .B1(n62189), .B2(n58664), .A(n79661), .ZN(n104338) );
  NAND2_X1 U64760 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [14]), .A2(n106358), 
        .ZN(n79661) );
  OAI21_X1 U64761 ( .B1(n62189), .B2(n58656), .A(n79662), .ZN(n104339) );
  NAND2_X1 U64762 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [13]), .A2(n106358), 
        .ZN(n79662) );
  OAI21_X1 U64763 ( .B1(n62189), .B2(n58653), .A(n79663), .ZN(n104340) );
  NAND2_X1 U64764 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [11]), .A2(n106358), 
        .ZN(n79663) );
  OAI21_X1 U64765 ( .B1(n62189), .B2(n58651), .A(n79664), .ZN(n104341) );
  NAND2_X1 U64766 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [10]), .A2(n106358), 
        .ZN(n79664) );
  OAI21_X1 U64767 ( .B1(n62189), .B2(n58647), .A(n79665), .ZN(n104342) );
  NAND2_X1 U64768 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [3]), .A2(n106358), 
        .ZN(n79665) );
  OAI21_X1 U64769 ( .B1(n62189), .B2(n58635), .A(n79666), .ZN(n104343) );
  NAND2_X1 U64770 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [1]), .A2(n106358), 
        .ZN(n79666) );
  OAI21_X1 U64771 ( .B1(n62189), .B2(n58632), .A(n79667), .ZN(n104344) );
  NAND2_X1 U64772 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [2]), .A2(n106358), 
        .ZN(n79667) );
  OAI21_X1 U64773 ( .B1(n62189), .B2(n58629), .A(n79668), .ZN(n104345) );
  NAND2_X1 U64774 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [7]), .A2(n106358), 
        .ZN(n79668) );
  OAI21_X1 U64775 ( .B1(n62189), .B2(n58624), .A(n79669), .ZN(n104346) );
  NAND2_X1 U64776 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [6]), .A2(n106358), 
        .ZN(n79669) );
  OAI21_X1 U64777 ( .B1(n62189), .B2(n58618), .A(n79670), .ZN(n104347) );
  NAND2_X1 U64778 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [4]), .A2(n106358), 
        .ZN(n79670) );
  OAI21_X1 U64779 ( .B1(n62189), .B2(n58614), .A(n79671), .ZN(n104348) );
  NAND2_X1 U64780 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [5]), .A2(n62189), 
        .ZN(n79671) );
  OAI21_X1 U64781 ( .B1(n62189), .B2(n58609), .A(n79672), .ZN(n104349) );
  NAND2_X1 U64782 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [9]), .A2(n62189), 
        .ZN(n79672) );
  OAI21_X1 U64783 ( .B1(n62189), .B2(n58604), .A(n79673), .ZN(n104350) );
  NAND2_X1 U64784 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [8]), .A2(n62189), 
        .ZN(n79673) );
  OAI21_X1 U64785 ( .B1(n62189), .B2(n58596), .A(n79674), .ZN(n104351) );
  NAND2_X1 U64786 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [19]), .A2(n62189), 
        .ZN(n79674) );
  OAI21_X1 U64787 ( .B1(n62189), .B2(n58594), .A(n79675), .ZN(n104352) );
  NAND2_X1 U64788 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [18]), .A2(n62189), 
        .ZN(n79675) );
  OAI21_X1 U64789 ( .B1(n62189), .B2(n58592), .A(n79676), .ZN(n104353) );
  NAND2_X1 U64790 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [17]), .A2(n62189), 
        .ZN(n79676) );
  OAI21_X1 U64791 ( .B1(n62189), .B2(n58588), .A(n79677), .ZN(n104354) );
  NAND2_X1 U64792 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [16]), .A2(n62189), 
        .ZN(n79677) );
  OAI21_X1 U64793 ( .B1(n62189), .B2(n58577), .A(n79678), .ZN(n104355) );
  NAND2_X1 U64794 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [23]), .A2(n62189), 
        .ZN(n79678) );
  OAI21_X1 U64795 ( .B1(n106358), .B2(n58575), .A(n79679), .ZN(n104356) );
  NAND2_X1 U64796 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [22]), .A2(n106358), 
        .ZN(n79679) );
  OAI21_X1 U64797 ( .B1(n62189), .B2(n58570), .A(n79680), .ZN(n104357) );
  NAND2_X1 U64798 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [21]), .A2(n62189), 
        .ZN(n79680) );
  OAI21_X1 U64799 ( .B1(n106358), .B2(n58565), .A(n79681), .ZN(n104358) );
  NAND2_X1 U64800 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [20]), .A2(n106358), 
        .ZN(n79681) );
  NOR4_X1 U64801 ( .A1(n79707), .A2(n79708), .A3(n79709), .A4(n79710), .ZN(
        n79706) );
  NOR2_X1 U64802 ( .A1(n79711), .A2(n107950), .ZN(n79710) );
  AOI22_X1 U64803 ( .A1(n79712), .A2(n107949), .B1(n79713), .B2(
        \DLX_Datapath/ArithLogUnit/A_log [31]), .ZN(n79711) );
  NOR3_X1 U64804 ( .A1(n107949), .A2(\DLX_Datapath/ArithLogUnit/B_log [31]), 
        .A3(n106357), .ZN(n79709) );
  OAI21_X1 U64805 ( .B1(n106926), .B2(n106954), .A(n79715), .ZN(n79708) );
  NAND2_X1 U64806 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N39 ), .A2(
        n106356), .ZN(n79715) );
  OAI21_X1 U64807 ( .B1(n106948), .B2(n79703), .A(n79717), .ZN(n79707) );
  AOI22_X1 U64808 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N71 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N103 ), .B2(n79719), .ZN(n79717) );
  AOI22_X1 U64809 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_1 [3]), .A2(
        n107591), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_0 [3]), .B2(
        n79720), .ZN(n79703) );
  NOR4_X1 U64810 ( .A1(n79722), .A2(n79723), .A3(n79724), .A4(n79725), .ZN(
        n79721) );
  NOR2_X1 U64811 ( .A1(n79726), .A2(n110956), .ZN(n79725) );
  AOI22_X1 U64812 ( .A1(n79712), .A2(n108045), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [30]), .B2(n79713), .ZN(n79726) );
  NOR3_X1 U64813 ( .A1(n108045), .A2(\DLX_Datapath/ArithLogUnit/B_log [30]), 
        .A3(n106357), .ZN(n79724) );
  OAI21_X1 U64814 ( .B1(n106924), .B2(n106954), .A(n79727), .ZN(n79723) );
  NAND2_X1 U64815 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N38 ), .A2(
        n106356), .ZN(n79727) );
  OAI21_X1 U64816 ( .B1(n106948), .B2(n79704), .A(n79728), .ZN(n79722) );
  AOI22_X1 U64817 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N70 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N102 ), .B2(n79719), .ZN(n79728) );
  AOI22_X1 U64818 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_1 [2]), .A2(
        n107591), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_0 [2]), .B2(
        n79720), .ZN(n79704) );
  NOR4_X1 U64819 ( .A1(n79730), .A2(n79731), .A3(n79732), .A4(n79733), .ZN(
        n79729) );
  NOR2_X1 U64820 ( .A1(n79734), .A2(n107574), .ZN(n79733) );
  AOI22_X1 U64821 ( .A1(n79712), .A2(n107572), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [29]), .B2(n79713), .ZN(n79734) );
  NOR3_X1 U64822 ( .A1(n107572), .A2(\DLX_Datapath/ArithLogUnit/B_log [29]), 
        .A3(n106357), .ZN(n79732) );
  OAI21_X1 U64823 ( .B1(n106840), .B2(n106954), .A(n79735), .ZN(n79731) );
  NAND2_X1 U64824 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N37 ), .A2(
        n106356), .ZN(n79735) );
  OAI21_X1 U64825 ( .B1(n106948), .B2(n79705), .A(n79736), .ZN(n79730) );
  AOI22_X1 U64826 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N69 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N101 ), .B2(n79719), .ZN(n79736) );
  AOI22_X1 U64827 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_1 [1]), .A2(
        n107591), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/S_0 [1]), .B2(
        n79720), .ZN(n79705) );
  NAND4_X2 U64828 ( .A1(n79737), .A2(n79738), .A3(n79739), .A4(n79740), .ZN(
        n103915) );
  AOI22_X1 U64831 ( .A1(n79712), .A2(n107854), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [28]), .B2(n79713), .ZN(n79743) );
  NOR2_X1 U64832 ( .A1(\DLX_Datapath/ArithLogUnit/B_log [28]), .A2(n106357), 
        .ZN(n79741) );
  AOI22_X1 U64833 ( .A1(n104366), .A2(n79744), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N36 ), .B2(n79716), .ZN(n79739)
         );
  XOR2_X1 U64834 ( .A(n79745), .B(n79720), .Z(n104366) );
  XNOR2_X1 U64835 ( .A(\DLX_Datapath/ArithLogUnit/A_add [28]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [28]), .ZN(n79745) );
  NAND2_X1 U64836 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N100 ), .A2(
        n79719), .ZN(n79738) );
  AOI22_X1 U64837 ( .A1(n105123), .A2(\DLX_Datapath/MUX_HDU_ALUInB [28]), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N68 ), .B2(n79718), .ZN(n79737)
         );
  NOR4_X1 U64838 ( .A1(n79748), .A2(n79749), .A3(n79750), .A4(n79751), .ZN(
        n79747) );
  NOR2_X1 U64839 ( .A1(n79752), .A2(n108046), .ZN(n79751) );
  AOI22_X1 U64840 ( .A1(n79712), .A2(n110748), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [27]), .B2(n79713), .ZN(n79752) );
  NOR3_X1 U64841 ( .A1(n110748), .A2(\DLX_Datapath/ArithLogUnit/B_log [27]), 
        .A3(n106357), .ZN(n79750) );
  OAI21_X1 U64842 ( .B1(n106922), .B2(n106954), .A(n79753), .ZN(n79749) );
  NAND2_X1 U64843 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N35 ), .A2(
        n106356), .ZN(n79753) );
  OAI21_X1 U64844 ( .B1(n106948), .B2(n79700), .A(n79754), .ZN(n79748) );
  AOI22_X1 U64845 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N67 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N99 ), .B2(n79719), .ZN(n79754) );
  AOI22_X1 U64846 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_1 [3]), .A2(
        n107596), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_0 [3]), .B2(
        n79755), .ZN(n79700) );
  NOR4_X1 U64847 ( .A1(n79757), .A2(n79758), .A3(n79759), .A4(n79760), .ZN(
        n79756) );
  NOR2_X1 U64848 ( .A1(n79761), .A2(n108155), .ZN(n79760) );
  AOI22_X1 U64849 ( .A1(n79712), .A2(n108153), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [26]), .B2(n79713), .ZN(n79761) );
  NOR3_X1 U64850 ( .A1(n108153), .A2(\DLX_Datapath/ArithLogUnit/B_log [26]), 
        .A3(n106357), .ZN(n79759) );
  OAI21_X1 U64851 ( .B1(n106920), .B2(n106954), .A(n79762), .ZN(n79758) );
  NAND2_X1 U64852 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N34 ), .A2(
        n106356), .ZN(n79762) );
  OAI21_X1 U64853 ( .B1(n106948), .B2(n79701), .A(n79763), .ZN(n79757) );
  AOI22_X1 U64854 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N66 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N98 ), .B2(n79719), .ZN(n79763) );
  AOI22_X1 U64855 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_1 [2]), .A2(
        n107596), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_0 [2]), .B2(
        n79755), .ZN(n79701) );
  NOR4_X1 U64856 ( .A1(n79765), .A2(n79766), .A3(n79767), .A4(n79768), .ZN(
        n79764) );
  NOR2_X1 U64857 ( .A1(n79769), .A2(n110954), .ZN(n79768) );
  AOI22_X1 U64858 ( .A1(n79712), .A2(n108156), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [25]), .B2(n79713), .ZN(n79769) );
  NOR3_X1 U64859 ( .A1(n108156), .A2(\DLX_Datapath/ArithLogUnit/B_log [25]), 
        .A3(n106357), .ZN(n79767) );
  OAI21_X1 U64860 ( .B1(n106918), .B2(n106954), .A(n79770), .ZN(n79766) );
  NAND2_X1 U64861 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N33 ), .A2(
        n106356), .ZN(n79770) );
  OAI21_X1 U64862 ( .B1(n106948), .B2(n79702), .A(n79771), .ZN(n79765) );
  AOI22_X1 U64863 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N65 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N97 ), .B2(n79719), .ZN(n79771) );
  AOI22_X1 U64864 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_1 [1]), .A2(
        n107596), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/S_0 [1]), .B2(
        n79755), .ZN(n79702) );
  NAND4_X2 U64865 ( .A1(n79772), .A2(n79773), .A3(n79774), .A4(n79775), .ZN(
        n103916) );
  AOI22_X1 U64868 ( .A1(n79712), .A2(n108157), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [24]), .B2(n79713), .ZN(n79778) );
  NOR2_X1 U64869 ( .A1(\DLX_Datapath/ArithLogUnit/B_log [24]), .A2(n106357), 
        .ZN(n79776) );
  AOI22_X1 U64870 ( .A1(n104365), .A2(n79744), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N32 ), .B2(n79716), .ZN(n79774)
         );
  XOR2_X1 U64871 ( .A(n107596), .B(n79779), .Z(n104365) );
  XOR2_X1 U64872 ( .A(\DLX_Datapath/ArithLogUnit/B_add [24]), .B(
        \DLX_Datapath/ArithLogUnit/A_add [24]), .Z(n79779) );
  NAND2_X1 U64873 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N96 ), .A2(n79719), .ZN(n79773) );
  AOI22_X1 U64874 ( .A1(n105123), .A2(\DLX_Datapath/MUX_HDU_ALUInB [24]), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N64 ), .B2(n79718), .ZN(n79772)
         );
  NOR4_X1 U64875 ( .A1(n79781), .A2(n79782), .A3(n79783), .A4(n79784), .ZN(
        n79780) );
  NOR2_X1 U64876 ( .A1(n79785), .A2(n110227), .ZN(n79784) );
  AOI22_X1 U64877 ( .A1(n79712), .A2(n110545), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [23]), .B2(n79713), .ZN(n79785) );
  NOR3_X1 U64878 ( .A1(n110545), .A2(\DLX_Datapath/ArithLogUnit/B_log [23]), 
        .A3(n79714), .ZN(n79783) );
  OAI21_X1 U64879 ( .B1(n106916), .B2(n106954), .A(n79786), .ZN(n79782) );
  NAND2_X1 U64880 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N31 ), .A2(
        n106356), .ZN(n79786) );
  OAI21_X1 U64881 ( .B1(n106948), .B2(n79697), .A(n79787), .ZN(n79781) );
  AOI22_X1 U64882 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N63 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N95 ), .B2(n79719), .ZN(n79787) );
  AOI22_X1 U64883 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_0 [3]), .A2(
        n107586), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_1 [3]), .B2(
        n79788), .ZN(n79697) );
  NOR4_X1 U64884 ( .A1(n79790), .A2(n79791), .A3(n79792), .A4(n79793), .ZN(
        n79789) );
  NOR2_X1 U64885 ( .A1(n79794), .A2(n110333), .ZN(n79793) );
  AOI22_X1 U64886 ( .A1(n79712), .A2(n110330), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [22]), .B2(n79713), .ZN(n79794) );
  NOR3_X1 U64887 ( .A1(n110330), .A2(\DLX_Datapath/ArithLogUnit/B_log [22]), 
        .A3(n106357), .ZN(n79792) );
  OAI21_X1 U64888 ( .B1(n106914), .B2(n106954), .A(n79795), .ZN(n79791) );
  NAND2_X1 U64889 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N30 ), .A2(
        n106356), .ZN(n79795) );
  OAI21_X1 U64890 ( .B1(n106948), .B2(n79698), .A(n79796), .ZN(n79790) );
  AOI22_X1 U64891 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N62 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N94 ), .B2(n79719), .ZN(n79796) );
  AOI22_X1 U64892 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_0 [2]), .A2(
        n107586), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_1 [2]), .B2(
        n79788), .ZN(n79698) );
  NOR4_X1 U64893 ( .A1(n79798), .A2(n79799), .A3(n79800), .A4(n79801), .ZN(
        n79797) );
  NOR2_X1 U64894 ( .A1(n79802), .A2(n110653), .ZN(n79801) );
  AOI22_X1 U64895 ( .A1(n79712), .A2(n110650), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [21]), .B2(n79713), .ZN(n79802) );
  NOR3_X1 U64896 ( .A1(n110650), .A2(\DLX_Datapath/ArithLogUnit/B_log [21]), 
        .A3(n79714), .ZN(n79800) );
  OAI21_X1 U64897 ( .B1(n106912), .B2(n106954), .A(n79803), .ZN(n79799) );
  NAND2_X1 U64898 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N29 ), .A2(
        n106356), .ZN(n79803) );
  OAI21_X1 U64899 ( .B1(n106948), .B2(n79699), .A(n79804), .ZN(n79798) );
  AOI22_X1 U64900 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N61 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N93 ), .B2(n79719), .ZN(n79804) );
  AOI22_X1 U64901 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_0 [1]), .A2(
        n107586), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/S_1 [1]), .B2(
        n79788), .ZN(n79699) );
  NAND4_X2 U64902 ( .A1(n79805), .A2(n79806), .A3(n79807), .A4(n79808), .ZN(
        n103917) );
  AOI22_X1 U64905 ( .A1(n79712), .A2(n110440), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [20]), .B2(n79713), .ZN(n79811) );
  NOR2_X1 U64906 ( .A1(\DLX_Datapath/ArithLogUnit/B_log [20]), .A2(n106357), 
        .ZN(n79809) );
  AOI22_X1 U64907 ( .A1(n104364), .A2(n79744), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N28 ), .B2(n79716), .ZN(n79807)
         );
  XOR2_X1 U64908 ( .A(n79788), .B(n79812), .Z(n104364) );
  XOR2_X1 U64909 ( .A(\DLX_Datapath/ArithLogUnit/B_add [20]), .B(
        \DLX_Datapath/ArithLogUnit/A_add [20]), .Z(n79812) );
  NAND2_X1 U64910 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N92 ), .A2(n79719), .ZN(n79806) );
  AOI22_X1 U64911 ( .A1(n105123), .A2(\DLX_Datapath/MUX_HDU_ALUInB [20]), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N60 ), .B2(n79718), .ZN(n79805)
         );
  NOR4_X1 U64912 ( .A1(n79814), .A2(n79815), .A3(n79816), .A4(n79817), .ZN(
        n79813) );
  NOR2_X1 U64913 ( .A1(n79818), .A2(n109778), .ZN(n79817) );
  AOI22_X1 U64914 ( .A1(n79712), .A2(n110117), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [19]), .B2(n79713), .ZN(n79818) );
  NOR3_X1 U64915 ( .A1(n110117), .A2(\DLX_Datapath/ArithLogUnit/B_log [19]), 
        .A3(n79714), .ZN(n79816) );
  OAI21_X1 U64916 ( .B1(n106910), .B2(n106954), .A(n79819), .ZN(n79815) );
  NAND2_X1 U64917 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N27 ), .A2(
        n106356), .ZN(n79819) );
  OAI21_X1 U64918 ( .B1(n106948), .B2(n79694), .A(n79820), .ZN(n79814) );
  AOI22_X1 U64919 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N59 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N91 ), .B2(n79719), .ZN(n79820) );
  AOI22_X1 U64920 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_1 [3]), .A2(
        n107582), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_0 [3]), .B2(
        n79821), .ZN(n79694) );
  NOR4_X1 U64921 ( .A1(n79823), .A2(n79824), .A3(n79825), .A4(n79826), .ZN(
        n79822) );
  NOR2_X1 U64922 ( .A1(n79827), .A2(n109780), .ZN(n79826) );
  AOI22_X1 U64923 ( .A1(n79712), .A2(n110224), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [18]), .B2(n79713), .ZN(n79827) );
  NOR3_X1 U64924 ( .A1(n110224), .A2(\DLX_Datapath/ArithLogUnit/B_log [18]), 
        .A3(n106357), .ZN(n79825) );
  OAI21_X1 U64925 ( .B1(n106908), .B2(n106954), .A(n79828), .ZN(n79824) );
  NAND2_X1 U64926 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N26 ), .A2(
        n106356), .ZN(n79828) );
  OAI21_X1 U64927 ( .B1(n106948), .B2(n79695), .A(n79829), .ZN(n79823) );
  AOI22_X1 U64928 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N58 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N90 ), .B2(n79719), .ZN(n79829) );
  AOI22_X1 U64929 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_1 [2]), .A2(
        n107582), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_0 [2]), .B2(
        n79821), .ZN(n79695) );
  NOR4_X1 U64930 ( .A1(n79831), .A2(n79832), .A3(n79833), .A4(n79834), .ZN(
        n79830) );
  NOR2_X1 U64931 ( .A1(n79835), .A2(n110011), .ZN(n79834) );
  AOI22_X1 U64932 ( .A1(n79712), .A2(n110009), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [17]), .B2(n79713), .ZN(n79835) );
  NOR3_X1 U64933 ( .A1(n110009), .A2(\DLX_Datapath/ArithLogUnit/B_log [17]), 
        .A3(n79714), .ZN(n79833) );
  OAI21_X1 U64934 ( .B1(n106906), .B2(n106954), .A(n79836), .ZN(n79832) );
  NAND2_X1 U64935 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N25 ), .A2(
        n106356), .ZN(n79836) );
  OAI21_X1 U64936 ( .B1(n106948), .B2(n79696), .A(n79837), .ZN(n79831) );
  AOI22_X1 U64937 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N57 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N89 ), .B2(n79719), .ZN(n79837) );
  AOI22_X1 U64938 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_1 [1]), .A2(
        n107582), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_4/S_0 [1]), .B2(
        n79821), .ZN(n79696) );
  NAND4_X2 U64939 ( .A1(n79838), .A2(n79839), .A3(n79840), .A4(n79841), .ZN(
        n103918) );
  AOI22_X1 U64942 ( .A1(n79712), .A2(n109896), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [16]), .B2(n79713), .ZN(n79844) );
  NOR2_X1 U64943 ( .A1(\DLX_Datapath/ArithLogUnit/B_log [16]), .A2(n106357), 
        .ZN(n79842) );
  AOI22_X1 U64944 ( .A1(n104363), .A2(n79744), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N24 ), .B2(n79716), .ZN(n79840)
         );
  XOR2_X1 U64945 ( .A(n79845), .B(n79821), .Z(n104363) );
  XNOR2_X1 U64946 ( .A(\DLX_Datapath/ArithLogUnit/A_add [16]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [16]), .ZN(n79845) );
  NAND2_X1 U64947 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N88 ), .A2(n79719), .ZN(n79839) );
  AOI22_X1 U64948 ( .A1(n105123), .A2(\DLX_Datapath/MUX_HDU_ALUInB [16]), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N56 ), .B2(n79718), .ZN(n79838)
         );
  NOR4_X1 U64949 ( .A1(n79847), .A2(n79848), .A3(n79849), .A4(n79850), .ZN(
        n79846) );
  NOR2_X1 U64950 ( .A1(n79851), .A2(n108274), .ZN(n79850) );
  AOI22_X1 U64951 ( .A1(n79712), .A2(n108269), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [15]), .B2(n79713), .ZN(n79851) );
  NOR3_X1 U64952 ( .A1(n108269), .A2(\DLX_Datapath/ArithLogUnit/B_log [15]), 
        .A3(n106357), .ZN(n79849) );
  OAI21_X1 U64953 ( .B1(n106904), .B2(n106954), .A(n79852), .ZN(n79848) );
  NAND2_X1 U64954 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N23 ), .A2(
        n106356), .ZN(n79852) );
  OAI21_X1 U64955 ( .B1(n106948), .B2(n79691), .A(n79853), .ZN(n79847) );
  AOI22_X1 U64956 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N55 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N87 ), .B2(n79719), .ZN(n79853) );
  AOI22_X1 U64957 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_1 [3]), .A2(
        n107604), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_0 [3]), .B2(
        n79854), .ZN(n79691) );
  NOR4_X1 U64958 ( .A1(n79856), .A2(n79857), .A3(n79858), .A4(n79859), .ZN(
        n79855) );
  NOR2_X1 U64959 ( .A1(n79860), .A2(n108393), .ZN(n79859) );
  AOI22_X1 U64960 ( .A1(n79712), .A2(n108390), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [14]), .B2(n79713), .ZN(n79860) );
  NOR3_X1 U64961 ( .A1(n108390), .A2(\DLX_Datapath/ArithLogUnit/B_log [14]), 
        .A3(n79714), .ZN(n79858) );
  OAI21_X1 U64962 ( .B1(n106902), .B2(n106954), .A(n79861), .ZN(n79857) );
  NAND2_X1 U64963 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N22 ), .A2(
        n106356), .ZN(n79861) );
  OAI21_X1 U64964 ( .B1(n106948), .B2(n79692), .A(n79862), .ZN(n79856) );
  AOI22_X1 U64965 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N54 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N86 ), .B2(n79719), .ZN(n79862) );
  AOI22_X1 U64966 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_1 [2]), .A2(
        n107604), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_0 [2]), .B2(
        n79854), .ZN(n79692) );
  NOR4_X1 U64967 ( .A1(n79864), .A2(n79865), .A3(n79866), .A4(n79867), .ZN(
        n79863) );
  NOR2_X1 U64968 ( .A1(n79868), .A2(n109773), .ZN(n79867) );
  AOI22_X1 U64969 ( .A1(n79712), .A2(n109768), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [13]), .B2(n79713), .ZN(n79868) );
  NOR3_X1 U64970 ( .A1(n109768), .A2(\DLX_Datapath/ArithLogUnit/B_log [13]), 
        .A3(n79714), .ZN(n79866) );
  OAI21_X1 U64971 ( .B1(n106900), .B2(n106954), .A(n79869), .ZN(n79865) );
  NAND2_X1 U64972 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N21 ), .A2(
        n106356), .ZN(n79869) );
  OAI21_X1 U64973 ( .B1(n106948), .B2(n79693), .A(n79870), .ZN(n79864) );
  AOI22_X1 U64974 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N53 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N85 ), .B2(n79719), .ZN(n79870) );
  AOI22_X1 U64975 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_1 [1]), .A2(
        n107604), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/S_0 [1]), .B2(
        n79854), .ZN(n79693) );
  NAND4_X2 U64976 ( .A1(n79871), .A2(n79872), .A3(n79873), .A4(n79874), .ZN(
        n103919) );
  AOI22_X1 U64979 ( .A1(n79712), .A2(n107743), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [12]), .B2(n79713), .ZN(n79877) );
  NOR2_X1 U64980 ( .A1(\DLX_Datapath/ArithLogUnit/B_log [12]), .A2(n106357), 
        .ZN(n79875) );
  AOI22_X1 U64981 ( .A1(n104362), .A2(n79744), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N20 ), .B2(n79716), .ZN(n79873)
         );
  XOR2_X1 U64982 ( .A(n79878), .B(n79854), .Z(n104362) );
  XNOR2_X1 U64983 ( .A(\DLX_Datapath/ArithLogUnit/A_add [12]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [12]), .ZN(n79878) );
  NAND2_X1 U64984 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N84 ), .A2(n79719), .ZN(n79872) );
  AOI22_X1 U64985 ( .A1(n105123), .A2(\DLX_Datapath/MUX_HDU_ALUInB [12]), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N52 ), .B2(n79718), .ZN(n79871)
         );
  NOR4_X1 U64986 ( .A1(n79880), .A2(n79881), .A3(n79882), .A4(n79883), .ZN(
        n79879) );
  NOR2_X1 U64987 ( .A1(n79884), .A2(n108506), .ZN(n79883) );
  AOI22_X1 U64988 ( .A1(n79712), .A2(n109653), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [11]), .B2(n79713), .ZN(n79884) );
  NOR3_X1 U64989 ( .A1(n109653), .A2(\DLX_Datapath/ArithLogUnit/B_log [11]), 
        .A3(n79714), .ZN(n79882) );
  OAI21_X1 U64990 ( .B1(n106898), .B2(n106954), .A(n79885), .ZN(n79881) );
  NAND2_X1 U64991 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N19 ), .A2(
        n106356), .ZN(n79885) );
  OAI21_X1 U64992 ( .B1(n106948), .B2(n79688), .A(n79886), .ZN(n79880) );
  AOI22_X1 U64993 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N51 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N83 ), .B2(n79719), .ZN(n79886) );
  AOI22_X1 U64994 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_1 [3]), .A2(
        n107609), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_0 [3]), .B2(
        n79887), .ZN(n79688) );
  NOR4_X1 U64995 ( .A1(n79889), .A2(n79890), .A3(n79891), .A4(n79892), .ZN(
        n79888) );
  NOR2_X1 U64996 ( .A1(n79893), .A2(n109767), .ZN(n79892) );
  AOI22_X1 U64997 ( .A1(n79712), .A2(n109765), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [10]), .B2(n79713), .ZN(n79893) );
  NOR3_X1 U64998 ( .A1(n109765), .A2(\DLX_Datapath/ArithLogUnit/B_log [10]), 
        .A3(n79714), .ZN(n79891) );
  OAI21_X1 U64999 ( .B1(n106896), .B2(n106954), .A(n79894), .ZN(n79890) );
  NAND2_X1 U65000 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N18 ), .A2(
        n106356), .ZN(n79894) );
  OAI21_X1 U65001 ( .B1(n106948), .B2(n79689), .A(n79895), .ZN(n79889) );
  AOI22_X1 U65002 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N50 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N82 ), .B2(n79719), .ZN(n79895) );
  AOI22_X1 U65003 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_1 [2]), .A2(
        n107609), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_0 [2]), .B2(
        n79887), .ZN(n79689) );
  NOR4_X1 U65004 ( .A1(n79897), .A2(n79898), .A3(n79899), .A4(n79900), .ZN(
        n79896) );
  NOR2_X1 U65005 ( .A1(n79901), .A2(n109763), .ZN(n79900) );
  AOI22_X1 U65006 ( .A1(n79712), .A2(n109760), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [9]), .B2(n79713), .ZN(n79901) );
  NOR3_X1 U65007 ( .A1(n109760), .A2(\DLX_Datapath/ArithLogUnit/B_log [9]), 
        .A3(n79714), .ZN(n79899) );
  OAI21_X1 U65008 ( .B1(n106894), .B2(n106954), .A(n79902), .ZN(n79898) );
  NAND2_X1 U65009 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N17 ), .A2(
        n106356), .ZN(n79902) );
  OAI21_X1 U65010 ( .B1(n106948), .B2(n79690), .A(n79903), .ZN(n79897) );
  AOI22_X1 U65011 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N49 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N81 ), .B2(n79719), .ZN(n79903) );
  AOI22_X1 U65012 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_1 [1]), .A2(
        n107609), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/S_0 [1]), .B2(
        n79887), .ZN(n79690) );
  NAND4_X2 U65013 ( .A1(n79904), .A2(n79905), .A3(n79906), .A4(n79907), .ZN(
        n103920) );
  AOI22_X1 U65016 ( .A1(n79712), .A2(n109546), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [8]), .B2(n79713), .ZN(n79910) );
  NOR2_X1 U65017 ( .A1(\DLX_Datapath/ArithLogUnit/B_log [8]), .A2(n106357), 
        .ZN(n79908) );
  AOI22_X1 U65018 ( .A1(n104361), .A2(n79744), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N16 ), .B2(n79716), .ZN(n79906)
         );
  XOR2_X1 U65019 ( .A(n79911), .B(n79887), .Z(n104361) );
  XNOR2_X1 U65020 ( .A(\DLX_Datapath/ArithLogUnit/A_add [8]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [8]), .ZN(n79911) );
  NAND2_X1 U65021 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N80 ), .A2(n79719), .ZN(n79905) );
  AOI22_X1 U65022 ( .A1(n105123), .A2(\DLX_Datapath/MUX_HDU_ALUInB [8]), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N48 ), .B2(n79718), .ZN(n79904)
         );
  NOR4_X1 U65023 ( .A1(n79913), .A2(n79914), .A3(n79915), .A4(n79916), .ZN(
        n79912) );
  NOR2_X1 U65024 ( .A1(n79917), .A2(n109091), .ZN(n79916) );
  AOI22_X1 U65025 ( .A1(n79712), .A2(n109083), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [7]), .B2(n79713), .ZN(n79917) );
  NOR3_X1 U65026 ( .A1(n109083), .A2(\DLX_Datapath/ArithLogUnit/B_log [7]), 
        .A3(n79714), .ZN(n79915) );
  OAI21_X1 U65027 ( .B1(n106892), .B2(n106954), .A(n79918), .ZN(n79914) );
  NAND2_X1 U65028 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N15 ), .A2(
        n106356), .ZN(n79918) );
  OAI21_X1 U65029 ( .B1(n106948), .B2(n79685), .A(n79919), .ZN(n79913) );
  AOI22_X1 U65030 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N47 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N79 ), .B2(n79719), .ZN(n79919) );
  AOI22_X1 U65031 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_1 [3]), .A2(
        n107615), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_0 [3]), .B2(
        n79920), .ZN(n79685) );
  NOR4_X1 U65032 ( .A1(n79922), .A2(n79923), .A3(n79924), .A4(n79925), .ZN(
        n79921) );
  NOR2_X1 U65033 ( .A1(n79926), .A2(n109434), .ZN(n79925) );
  AOI22_X1 U65034 ( .A1(n79712), .A2(n109430), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [6]), .B2(n79713), .ZN(n79926) );
  NOR3_X1 U65035 ( .A1(n109430), .A2(\DLX_Datapath/ArithLogUnit/B_log [6]), 
        .A3(n79714), .ZN(n79924) );
  OAI21_X1 U65036 ( .B1(n106890), .B2(n106954), .A(n79927), .ZN(n79923) );
  NAND2_X1 U65037 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N14 ), .A2(n79716), .ZN(n79927) );
  OAI21_X1 U65038 ( .B1(n106948), .B2(n79686), .A(n79928), .ZN(n79922) );
  AOI22_X1 U65039 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N46 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N78 ), .B2(n79719), .ZN(n79928) );
  AOI22_X1 U65040 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_1 [2]), .A2(
        n107615), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_0 [2]), .B2(
        n79920), .ZN(n79686) );
  NOR4_X1 U65041 ( .A1(n79930), .A2(n79931), .A3(n79932), .A4(n79933), .ZN(
        n79929) );
  NOR2_X1 U65042 ( .A1(n79934), .A2(n109311), .ZN(n79933) );
  AOI22_X1 U65043 ( .A1(n79712), .A2(n109314), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [5]), .B2(n79713), .ZN(n79934) );
  NOR3_X1 U65044 ( .A1(n109314), .A2(\DLX_Datapath/ArithLogUnit/B_log [5]), 
        .A3(n79714), .ZN(n79932) );
  OAI21_X1 U65045 ( .B1(n106888), .B2(n106954), .A(n79935), .ZN(n79931) );
  NAND2_X1 U65046 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N13 ), .A2(n79716), .ZN(n79935) );
  OAI21_X1 U65047 ( .B1(n106948), .B2(n79687), .A(n79936), .ZN(n79930) );
  AOI22_X1 U65048 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N45 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N77 ), .B2(n79719), .ZN(n79936) );
  AOI22_X1 U65049 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_1 [1]), .A2(
        n107615), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/S_0 [1]), .B2(
        n79920), .ZN(n79687) );
  NAND4_X2 U65050 ( .A1(n79937), .A2(n79938), .A3(n79939), .A4(n79940), .ZN(
        n103921) );
  AOI22_X1 U65053 ( .A1(n79712), .A2(n109205), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [4]), .B2(n79713), .ZN(n79943) );
  NOR2_X1 U65054 ( .A1(\DLX_Datapath/ArithLogUnit/B_log [4]), .A2(n106357), 
        .ZN(n79941) );
  AOI22_X1 U65055 ( .A1(n104360), .A2(n79744), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N12 ), .B2(n79716), .ZN(n79939)
         );
  XOR2_X1 U65056 ( .A(n79944), .B(n79920), .Z(n104360) );
  XNOR2_X1 U65057 ( .A(\DLX_Datapath/ArithLogUnit/A_add [4]), .B(
        \DLX_Datapath/ArithLogUnit/B_add [4]), .ZN(n79944) );
  NAND2_X1 U65058 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N76 ), .A2(n79719), .ZN(n79938) );
  AOI22_X1 U65059 ( .A1(n105123), .A2(\DLX_Datapath/MUX_HDU_ALUInB [4]), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_shift/N44 ), .B2(n79718), .ZN(n79937)
         );
  NOR4_X1 U65060 ( .A1(n79946), .A2(n79947), .A3(n79948), .A4(n79949), .ZN(
        n79945) );
  NOR2_X1 U65061 ( .A1(n79950), .A2(n108746), .ZN(n79949) );
  AOI22_X1 U65062 ( .A1(n79712), .A2(n108738), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [3]), .B2(n79713), .ZN(n79950) );
  NOR3_X1 U65063 ( .A1(n108738), .A2(\DLX_Datapath/ArithLogUnit/B_log [3]), 
        .A3(n79714), .ZN(n79948) );
  OAI21_X1 U65064 ( .B1(n106886), .B2(n106954), .A(n79951), .ZN(n79947) );
  NAND2_X1 U65065 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N11 ), .A2(n79716), .ZN(n79951) );
  OAI21_X1 U65066 ( .B1(n106948), .B2(n79684), .A(n79952), .ZN(n79946) );
  AOI22_X1 U65067 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N43 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N75 ), .B2(n79719), .ZN(n79952) );
  AOI22_X1 U65068 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_0 [3]), .A2(
        n107578), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_1 [3]), .B2(
        \DLX_Datapath/ArithLogUnit/Cin_add ), .ZN(n79684) );
  NOR4_X1 U65069 ( .A1(n79954), .A2(n79955), .A3(n79956), .A4(n79957), .ZN(
        n79953) );
  NOR2_X1 U65070 ( .A1(n79958), .A2(n108970), .ZN(n79957) );
  AOI22_X1 U65071 ( .A1(n79712), .A2(n108967), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [2]), .B2(n79713), .ZN(n79958) );
  NOR3_X1 U65072 ( .A1(n108967), .A2(\DLX_Datapath/ArithLogUnit/B_log [2]), 
        .A3(n79714), .ZN(n79956) );
  OAI21_X1 U65073 ( .B1(n106884), .B2(n106954), .A(n79959), .ZN(n79955) );
  NAND2_X1 U65074 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N10 ), .A2(n79716), .ZN(n79959) );
  OAI21_X1 U65075 ( .B1(n106948), .B2(n79683), .A(n79960), .ZN(n79954) );
  AOI22_X1 U65076 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N42 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N74 ), .B2(n79719), .ZN(n79960) );
  AOI22_X1 U65077 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_0 [2]), .A2(
        n107578), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_1 [2]), .B2(
        \DLX_Datapath/ArithLogUnit/Cin_add ), .ZN(n79683) );
  NOR4_X1 U65078 ( .A1(n79962), .A2(n79963), .A3(n79964), .A4(n79965), .ZN(
        n79961) );
  NOR2_X1 U65079 ( .A1(n79966), .A2(n108859), .ZN(n79965) );
  AOI22_X1 U65080 ( .A1(n79712), .A2(n108856), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [1]), .B2(n79713), .ZN(n79966) );
  NOR3_X1 U65081 ( .A1(n108856), .A2(\DLX_Datapath/ArithLogUnit/B_log [1]), 
        .A3(n79714), .ZN(n79964) );
  OAI21_X1 U65082 ( .B1(n106882), .B2(n106954), .A(n79967), .ZN(n79963) );
  NAND2_X1 U65083 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N9 ), .A2(n106356), .ZN(n79967) );
  OAI21_X1 U65084 ( .B1(n106948), .B2(n79682), .A(n79968), .ZN(n79962) );
  AOI22_X1 U65085 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N41 ), .A2(n79718), .B1(\DLX_Datapath/ArithLogUnit/ALU_shift/N73 ), .B2(n79719), .ZN(n79968) );
  AOI22_X1 U65086 ( .A1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_0 [1]), .A2(
        n107578), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/S_1 [1]), .B2(
        \DLX_Datapath/ArithLogUnit/Cin_add ), .ZN(n79682) );
  AOI22_X1 U65087 ( .A1(\DLX_Datapath/next_B_IDEX [17]), .A2(n106355), .B1(
        n106353), .B2(n73120), .ZN(n79969) );
  AOI22_X1 U65088 ( .A1(\DLX_Datapath/next_B_IDEX [15]), .A2(n106354), .B1(
        n106353), .B2(n70872), .ZN(n79972) );
  AOI22_X1 U65089 ( .A1(\DLX_Datapath/next_B_IDEX [13]), .A2(n106355), .B1(
        n106353), .B2(n71169), .ZN(n79973) );
  AOI22_X1 U65090 ( .A1(\DLX_Datapath/next_B_IDEX [11]), .A2(n106355), .B1(
        n106353), .B2(n72661), .ZN(n79974) );
  AOI22_X1 U65091 ( .A1(\DLX_Datapath/next_B_IDEX [9]), .A2(n106354), .B1(
        n106353), .B2(n72803), .ZN(n79975) );
  AOI22_X1 U65092 ( .A1(\DLX_Datapath/next_B_IDEX [7]), .A2(n106354), .B1(
        n106353), .B2(n71913), .ZN(n79976) );
  AOI22_X1 U65093 ( .A1(\DLX_Datapath/next_B_IDEX [31]), .A2(n106355), .B1(
        n106353), .B2(n70427), .ZN(n79977) );
  AOI22_X1 U65094 ( .A1(n106351), .A2(n106825), .B1(n69413), .B2(n106349), 
        .ZN(n79978) );
  AOI22_X1 U65095 ( .A1(n106350), .A2(n106826), .B1(n69414), .B2(n106349), 
        .ZN(n79981) );
  AOI22_X1 U65096 ( .A1(n106350), .A2(n108049), .B1(n70576), .B2(n106349), 
        .ZN(n79982) );
  AOI22_X1 U65097 ( .A1(net2410613), .A2(n106350), .B1(n70575), .B2(n106349), 
        .ZN(n79983) );
  AOI22_X1 U65098 ( .A1(n106350), .A2(n106822), .B1(n69417), .B2(n106349), 
        .ZN(n79984) );
  AOI22_X1 U65099 ( .A1(n106350), .A2(n108158), .B1(n70726), .B2(n106349), 
        .ZN(n79985) );
  AOI22_X1 U65100 ( .A1(n106350), .A2(n108278), .B1(n70882), .B2(n106349), 
        .ZN(n79986) );
  AOI22_X1 U65101 ( .A1(n106350), .A2(n109437), .B1(n72372), .B2(n106349), 
        .ZN(n79987) );
  AOI22_X1 U65102 ( .A1(n106350), .A2(n109092), .B1(n71922), .B2(n106349), 
        .ZN(n79988) );
  AOI22_X1 U65103 ( .A1(n106350), .A2(n108621), .B1(n71327), .B2(n106348), 
        .ZN(n79989) );
  AOI22_X1 U65104 ( .A1(n106350), .A2(n106827), .B1(n69415), .B2(n106348), 
        .ZN(n79990) );
  AOI22_X1 U65105 ( .A1(n106350), .A2(n107747), .B1(n70142), .B2(n106348), 
        .ZN(n79991) );
  AOI22_X1 U65106 ( .A1(n106351), .A2(n110228), .B1(n73411), .B2(n106348), 
        .ZN(n79992) );
  AOI22_X1 U65107 ( .A1(n106351), .A2(n110336), .B1(n73560), .B2(n106348), 
        .ZN(n79993) );
  AOI22_X1 U65108 ( .A1(n106351), .A2(n109783), .B1(n72830), .B2(n106348), 
        .ZN(n79994) );
  AOI22_X1 U65109 ( .A1(n106351), .A2(n109899), .B1(n72978), .B2(n106348), 
        .ZN(n79995) );
  AOI22_X1 U65110 ( .A1(n106351), .A2(n108276), .B1(n70880), .B2(n106348), 
        .ZN(n79996) );
  AOI22_X1 U65111 ( .A1(n106351), .A2(n108508), .B1(n71179), .B2(n106348), 
        .ZN(n79997) );
  AOI22_X1 U65112 ( .A1(n106351), .A2(n108972), .B1(n71772), .B2(n106348), 
        .ZN(n79998) );
  AOI22_X1 U65113 ( .A1(n106351), .A2(n109094), .B1(n71924), .B2(n106348), 
        .ZN(n79999) );
  AOI22_X1 U65114 ( .A1(n106351), .A2(n108619), .B1(n71325), .B2(n106348), 
        .ZN(n80000) );
  NOR2_X1 U65115 ( .A1(n100795), .A2(net113156), .ZN(n103922) );
  NOR2_X1 U65116 ( .A1(n100779), .A2(net113155), .ZN(n103923) );
  NOR2_X1 U65117 ( .A1(n100770), .A2(net113159), .ZN(n103924) );
  NOR2_X1 U65118 ( .A1(n62247), .A2(net113159), .ZN(n103925) );
  NOR2_X1 U65119 ( .A1(n100784), .A2(net113157), .ZN(n103926) );
  AOI22_X1 U65120 ( .A1(\DLX_Datapath/next_B_IDEX [29]), .A2(n106354), .B1(
        n106353), .B2(n69307), .ZN(n80002) );
  AOI22_X1 U65121 ( .A1(\DLX_Datapath/next_B_IDEX [28]), .A2(n106355), .B1(
        n106353), .B2(n70283), .ZN(n80003) );
  AOI22_X1 U65122 ( .A1(\DLX_Datapath/next_B_IDEX [27]), .A2(n106354), .B1(
        n106352), .B2(n74130), .ZN(n80004) );
  AOI22_X1 U65123 ( .A1(\DLX_Datapath/next_B_IDEX [26]), .A2(n79970), .B1(
        n106352), .B2(n70717), .ZN(n80005) );
  AOI22_X1 U65124 ( .A1(\DLX_Datapath/next_B_IDEX [25]), .A2(n106355), .B1(
        n106352), .B2(n74270), .ZN(n80006) );
  AOI22_X1 U65125 ( .A1(\DLX_Datapath/next_B_IDEX [24]), .A2(n106355), .B1(
        n106352), .B2(n74410), .ZN(n80007) );
  AOI22_X1 U65126 ( .A1(\DLX_Datapath/next_B_IDEX [23]), .A2(n106354), .B1(
        n106352), .B2(n73847), .ZN(n80008) );
  AOI22_X1 U65127 ( .A1(\DLX_Datapath/next_B_IDEX [22]), .A2(n79970), .B1(
        n106352), .B2(n73552), .ZN(n80009) );
  AOI22_X1 U65128 ( .A1(\DLX_Datapath/next_B_IDEX [21]), .A2(n106355), .B1(
        n106352), .B2(n73988), .ZN(n80010) );
  AOI22_X1 U65129 ( .A1(\DLX_Datapath/next_B_IDEX [20]), .A2(n106354), .B1(
        n106352), .B2(n73699), .ZN(n80011) );
  AOI22_X1 U65130 ( .A1(\DLX_Datapath/next_B_IDEX [19]), .A2(n79970), .B1(
        n106352), .B2(n73263), .ZN(n80012) );
  AOI22_X1 U65131 ( .A1(\DLX_Datapath/next_B_IDEX [5]), .A2(n106355), .B1(
        n106352), .B2(n72209), .ZN(n80013) );
  AOI22_X1 U65132 ( .A1(\DLX_Datapath/next_B_IDEX [1]), .A2(n106354), .B1(
        n106352), .B2(n71618), .ZN(n80014) );
  AOI22_X1 U65133 ( .A1(\DLX_Datapath/next_B_IDEX [30]), .A2(n106355), .B1(
        n106352), .B2(n70569), .ZN(n80015) );
  AOI22_X1 U65134 ( .A1(\DLX_Datapath/next_B_IDEX [18]), .A2(n106354), .B1(
        n106353), .B2(n73405), .ZN(n80016) );
  AOI22_X1 U65135 ( .A1(\DLX_Datapath/next_B_IDEX [16]), .A2(n79970), .B1(
        n79971), .B2(n72969), .ZN(n80017) );
  AOI22_X1 U65136 ( .A1(\DLX_Datapath/next_B_IDEX [14]), .A2(n106355), .B1(
        n106353), .B2(n71026), .ZN(n80018) );
  AOI22_X1 U65137 ( .A1(\DLX_Datapath/next_B_IDEX [12]), .A2(n106354), .B1(
        n106353), .B2(n70130), .ZN(n80019) );
  AOI22_X1 U65138 ( .A1(\DLX_Datapath/next_B_IDEX [10]), .A2(n79970), .B1(
        n79971), .B2(n72808), .ZN(n80020) );
  AOI22_X1 U65139 ( .A1(\DLX_Datapath/next_B_IDEX [8]), .A2(n106355), .B1(
        n79971), .B2(n72511), .ZN(n80021) );
  AOI22_X1 U65140 ( .A1(\DLX_Datapath/next_B_IDEX [6]), .A2(n106354), .B1(
        n79971), .B2(n72362), .ZN(n80022) );
  AOI22_X1 U65141 ( .A1(\DLX_Datapath/next_B_IDEX [4]), .A2(n79970), .B1(
        n79971), .B2(n72065), .ZN(n80023) );
  AOI22_X1 U65142 ( .A1(\DLX_Datapath/next_B_IDEX [3]), .A2(n106355), .B1(
        n79971), .B2(n71469), .ZN(n80024) );
  AOI22_X1 U65143 ( .A1(\DLX_Datapath/next_B_IDEX [2]), .A2(n106354), .B1(
        n79971), .B2(n71762), .ZN(n80025) );
  AOI22_X1 U65144 ( .A1(\DLX_Datapath/next_B_IDEX [0]), .A2(n106354), .B1(
        n69292), .B2(n106353), .ZN(n80026) );
  NOR2_X1 U65145 ( .A1(net113155), .A2(n79971), .ZN(n79970) );
  NOR2_X1 U65146 ( .A1(n107417), .A2(net113154), .ZN(n79971) );
  AOI22_X1 U65147 ( .A1(n106351), .A2(n106828), .B1(n69303), .B2(n106349), 
        .ZN(n80027) );
  AOI22_X1 U65148 ( .A1(n106351), .A2(n108051), .B1(n70577), .B2(n106349), 
        .ZN(n80028) );
  AOI22_X1 U65149 ( .A1(n106351), .A2(n106824), .B1(n69416), .B2(n106349), 
        .ZN(n80029) );
  AOI22_X1 U65150 ( .A1(n106351), .A2(n110334), .B1(n73558), .B2(n106349), 
        .ZN(n80030) );
  AOI22_X1 U65151 ( .A1(n79979), .A2(n109901), .B1(n72980), .B2(n79980), .ZN(
        n80031) );
  AOI22_X1 U65152 ( .A1(n79979), .A2(n108280), .B1(n70884), .B2(n79980), .ZN(
        n80032) );
  AOI22_X1 U65153 ( .A1(n79979), .A2(n107621), .B1(n69991), .B2(n79980), .ZN(
        n80033) );
  AOI22_X1 U65154 ( .A1(n79979), .A2(n109435), .B1(n72370), .B2(n79980), .ZN(
        n80034) );
  AOI22_X1 U65155 ( .A1(n106351), .A2(n109096), .B1(n71926), .B2(n79980), .ZN(
        n80035) );
  AOI22_X1 U65156 ( .A1(n106350), .A2(n108631), .B1(n71329), .B2(n79980), .ZN(
        n80036) );
  AOI22_X1 U65157 ( .A1(n106350), .A2(n106765), .B1(n69289), .B2(n79980), .ZN(
        n80037) );
  NOR2_X1 U65158 ( .A1(net113159), .A2(n79980), .ZN(n79979) );
  NOR2_X1 U65159 ( .A1(net113154), .A2(n100718), .ZN(n79980) );
  OAI21_X1 U65160 ( .B1(n100779), .B2(net113091), .A(n106598), .ZN(n103927) );
  NOR3_X1 U65161 ( .A1(n80039), .A2(n80040), .A3(n105152), .ZN(n80038) );
  AOI22_X1 U65162 ( .A1(IR_in[28]), .A2(n80042), .B1(n111145), .B2(n111143), 
        .ZN(n80040) );
  AOI22_X1 U65163 ( .A1(IR_in[1]), .A2(n105163), .B1(n69350), .B2(net113156), 
        .ZN(n80043) );
  AOI22_X1 U65164 ( .A1(IR_in[2]), .A2(n105165), .B1(n69351), .B2(net113156), 
        .ZN(n80044) );
  AOI22_X1 U65165 ( .A1(IR_in[3]), .A2(n105163), .B1(n69352), .B2(net113156), 
        .ZN(n80045) );
  AOI22_X1 U65166 ( .A1(IR_in[11]), .A2(n105164), .B1(net113156), .B2(
        \DLX_Datapath/IR_IFID[11] ), .ZN(n80046) );
  AOI22_X1 U65167 ( .A1(IR_in[14]), .A2(n105162), .B1(n69362), .B2(net113159), 
        .ZN(n80047) );
  AOI22_X1 U65168 ( .A1(IR_in[15]), .A2(n105165), .B1(n69369), .B2(net113157), 
        .ZN(n80048) );
  AOI22_X1 U65169 ( .A1(IR_in[16]), .A2(n105163), .B1(net113157), .B2(n107132), 
        .ZN(n80049) );
  AOI22_X1 U65170 ( .A1(IR_in[17]), .A2(n105164), .B1(net113155), .B2(n107134), 
        .ZN(n80050) );
  AOI22_X1 U65171 ( .A1(IR_in[19]), .A2(n105162), .B1(net113157), .B2(n107139), 
        .ZN(n80051) );
  AOI22_X1 U65172 ( .A1(IR_in[24]), .A2(n105165), .B1(net113155), .B2(n104707), 
        .ZN(n80052) );
  AOI22_X1 U65173 ( .A1(IR_in[27]), .A2(n105163), .B1(n69377), .B2(net113155), 
        .ZN(n80053) );
  AOI22_X1 U65174 ( .A1(IR_in[29]), .A2(n105164), .B1(n69379), .B2(net113156), 
        .ZN(n80054) );
  AOI22_X1 U65175 ( .A1(n80056), .A2(n105162), .B1(net113155), .B2(
        \DLX_ControlUnit/cw2 [13]), .ZN(n80055) );
  AOI22_X1 U65176 ( .A1(n105164), .A2(n111119), .B1(net113156), .B2(
        \DLX_ControlUnit/cw2 [6]), .ZN(n80057) );
  AOI22_X1 U65177 ( .A1(n105162), .A2(n111118), .B1(net113155), .B2(
        \DLX_ControlUnit/cw2 [2]), .ZN(n80058) );
  AOI22_X1 U65178 ( .A1(IR_in[6]), .A2(n105165), .B1(n69355), .B2(net113155), 
        .ZN(n80059) );
  AOI22_X1 U65179 ( .A1(IR_in[7]), .A2(n105163), .B1(n69356), .B2(net113159), 
        .ZN(n80060) );
  AOI22_X1 U65180 ( .A1(IR_in[10]), .A2(n105164), .B1(n69359), .B2(net113155), 
        .ZN(n80061) );
  AOI22_X1 U65181 ( .A1(n105162), .A2(IR_in[12]), .B1(net113159), .B2(
        \DLX_Datapath/IR_IFID[12] ), .ZN(n80062) );
  AOI22_X1 U65182 ( .A1(IR_in[25]), .A2(n105162), .B1(net113155), .B2(n104495), 
        .ZN(n80063) );
  OAI21_X1 U65183 ( .B1(n80064), .B2(n80065), .A(n80066), .ZN(n103928) );
  NAND2_X1 U65184 ( .A1(n69283), .A2(net113155), .ZN(n80066) );
  OR2_X1 U65185 ( .A1(n80067), .A2(n105152), .ZN(n80065) );
  AOI22_X1 U65186 ( .A1(n105163), .A2(n80069), .B1(n69765), .B2(net113159), 
        .ZN(n80068) );
  AOI22_X1 U65187 ( .A1(n80071), .A2(n105165), .B1(net113155), .B2(
        \DLX_ControlUnit/cw2 [7]), .ZN(n80070) );
  AOI22_X1 U65188 ( .A1(n105165), .A2(n80073), .B1(net113155), .B2(n104506), 
        .ZN(n80072) );
  AOI22_X1 U65189 ( .A1(IR_in[0]), .A2(n105163), .B1(n69349), .B2(net113159), 
        .ZN(n80074) );
  AOI22_X1 U65190 ( .A1(IR_in[4]), .A2(n105164), .B1(n69353), .B2(net113155), 
        .ZN(n80075) );
  AOI22_X1 U65191 ( .A1(IR_in[5]), .A2(n105162), .B1(n69354), .B2(net113157), 
        .ZN(n80076) );
  AOI22_X1 U65192 ( .A1(IR_in[8]), .A2(n105165), .B1(n69357), .B2(net113156), 
        .ZN(n80077) );
  AOI22_X1 U65193 ( .A1(IR_in[9]), .A2(n105164), .B1(n69358), .B2(net113155), 
        .ZN(n80078) );
  AOI22_X1 U65194 ( .A1(IR_in[13]), .A2(n105162), .B1(net113155), .B2(
        \DLX_Datapath/IR_IFID[13] ), .ZN(n80079) );
  AOI22_X1 U65195 ( .A1(IR_in[18]), .A2(n105165), .B1(net113155), .B2(n107137), 
        .ZN(n80080) );
  AOI22_X1 U65196 ( .A1(IR_in[20]), .A2(n105163), .B1(net113159), .B2(n107142), 
        .ZN(n80081) );
  AOI22_X1 U65197 ( .A1(IR_in[21]), .A2(n105162), .B1(net113157), .B2(n107144), 
        .ZN(n80082) );
  AOI22_X1 U65198 ( .A1(IR_in[22]), .A2(n105163), .B1(net113159), .B2(n107145), 
        .ZN(n80083) );
  AOI22_X1 U65199 ( .A1(IR_in[23]), .A2(n105164), .B1(net113157), .B2(n105061), 
        .ZN(n80084) );
  AOI22_X1 U65200 ( .A1(n80086), .A2(n105164), .B1(net113157), .B2(
        \DLX_ControlUnit/cw2 [10]), .ZN(n80085) );
  AOI22_X1 U65201 ( .A1(n105164), .A2(IR_in[31]), .B1(n69381), .B2(net113155), 
        .ZN(n80087) );
  AOI22_X1 U65202 ( .A1(n105165), .A2(n80069), .B1(net113155), .B2(n107417), 
        .ZN(n80088) );
  AOI22_X1 U65203 ( .A1(n80056), .A2(n105162), .B1(net113156), .B2(
        \DLX_ControlUnit/cw2 [15]), .ZN(n80089) );
  AOI22_X1 U65204 ( .A1(n105164), .A2(n111119), .B1(net113156), .B2(
        \DLX_ControlUnit/cw2 [0]), .ZN(n80090) );
  NOR3_X1 U65205 ( .A1(n80092), .A2(n111128), .A3(n111137), .ZN(n80091) );
  OAI21_X1 U65206 ( .B1(n80039), .B2(n80093), .A(n80094), .ZN(n103929) );
  NAND2_X1 U65207 ( .A1(net113156), .A2(\DLX_ControlUnit/cw2 [9]), .ZN(n80094)
         );
  NAND2_X1 U65208 ( .A1(n105163), .A2(n111145), .ZN(n80093) );
  AOI22_X1 U65209 ( .A1(n80071), .A2(n105165), .B1(net113159), .B2(
        \DLX_ControlUnit/cw2 [12]), .ZN(n80095) );
  OAI21_X1 U65210 ( .B1(n100770), .B2(net113102), .A(n80096), .ZN(n103930) );
  NOR2_X1 U65211 ( .A1(n80097), .A2(n80098), .ZN(n80096) );
  AOI21_X1 U65212 ( .B1(n80099), .B2(n80100), .A(n105152), .ZN(n80098) );
  OAI21_X1 U65213 ( .B1(n80101), .B2(n104734), .A(n80103), .ZN(n103931) );
  NAND2_X1 U65214 ( .A1(n106346), .A2(n106842), .ZN(n80103) );
  OAI21_X1 U65215 ( .B1(n106786), .B2(n104734), .A(n80105), .ZN(n103932) );
  NAND2_X1 U65216 ( .A1(n62198), .A2(n106346), .ZN(n80105) );
  OAI21_X1 U65217 ( .B1(n80107), .B2(n104734), .A(n80108), .ZN(n103933) );
  NAND2_X1 U65218 ( .A1(n106346), .A2(n109321), .ZN(n80108) );
  OAI21_X1 U65219 ( .B1(n80109), .B2(n104734), .A(n80110), .ZN(n103934) );
  NAND2_X1 U65220 ( .A1(n106346), .A2(n109322), .ZN(n80110) );
  OAI21_X1 U65221 ( .B1(n80111), .B2(n104734), .A(n80112), .ZN(n103935) );
  NAND2_X1 U65222 ( .A1(n106346), .A2(n109323), .ZN(n80112) );
  OAI21_X1 U65223 ( .B1(n80113), .B2(n104736), .A(n80114), .ZN(n103936) );
  NAND2_X1 U65224 ( .A1(n106346), .A2(n109549), .ZN(n80114) );
  OAI21_X1 U65225 ( .B1(n80115), .B2(n104737), .A(n80116), .ZN(n103937) );
  NAND2_X1 U65226 ( .A1(n106346), .A2(n109776), .ZN(n80116) );
  OAI21_X1 U65227 ( .B1(n80117), .B2(n104734), .A(n80118), .ZN(n103938) );
  NAND2_X1 U65228 ( .A1(n106346), .A2(n109777), .ZN(n80118) );
  OAI21_X1 U65229 ( .B1(n80119), .B2(n104737), .A(n80120), .ZN(n103939) );
  NAND2_X1 U65230 ( .A1(n106346), .A2(n109898), .ZN(n80120) );
  OAI21_X1 U65231 ( .B1(n106773), .B2(n104734), .A(n80121), .ZN(n103940) );
  NAND2_X1 U65232 ( .A1(n106346), .A2(n110958), .ZN(n80121) );
  NAND2_X1 U65234 ( .A1(n106346), .A2(n110964), .ZN(n80123) );
  OAI21_X1 U65235 ( .B1(n80125), .B2(n104734), .A(n80126), .ZN(n103942) );
  NAND2_X1 U65236 ( .A1(n106346), .A2(n110965), .ZN(n80126) );
  OAI21_X1 U65237 ( .B1(n106785), .B2(n104734), .A(n80127), .ZN(n103943) );
  NAND2_X1 U65238 ( .A1(n62197), .A2(n106346), .ZN(n80127) );
  OAI21_X1 U65239 ( .B1(n104734), .B2(n80129), .A(n80130), .ZN(n103944) );
  NAND2_X1 U65240 ( .A1(n106346), .A2(n107744), .ZN(n80130) );
  OAI21_X1 U65241 ( .B1(n80131), .B2(n104736), .A(n80132), .ZN(n103945) );
  NAND2_X1 U65242 ( .A1(n106346), .A2(n109547), .ZN(n80132) );
  OAI21_X1 U65243 ( .B1(n104736), .B2(n106791), .A(n80133), .ZN(n103946) );
  NAND2_X1 U65244 ( .A1(n106346), .A2(n109774), .ZN(n80133) );
  OAI21_X1 U65245 ( .B1(n106783), .B2(n104737), .A(n80135), .ZN(n103947) );
  NAND2_X1 U65246 ( .A1(n106346), .A2(n110966), .ZN(n80135) );
  OAI21_X1 U65247 ( .B1(n80137), .B2(n104737), .A(n80138), .ZN(n103948) );
  NAND2_X1 U65248 ( .A1(net2411291), .A2(n106346), .ZN(n80138) );
  OAI21_X1 U65249 ( .B1(n80139), .B2(n104734), .A(n80140), .ZN(n103949) );
  NAND2_X1 U65250 ( .A1(n106346), .A2(n109316), .ZN(n80140) );
  OAI21_X1 U65251 ( .B1(n80141), .B2(n104737), .A(n80142), .ZN(n103950) );
  NAND2_X1 U65252 ( .A1(n106346), .A2(n109548), .ZN(n80142) );
  OAI21_X1 U65253 ( .B1(n80143), .B2(n104734), .A(n80144), .ZN(n103951) );
  NAND2_X1 U65254 ( .A1(n106346), .A2(n109775), .ZN(n80144) );
  OAI21_X1 U65255 ( .B1(n104736), .B2(n106776), .A(n80145), .ZN(n103952) );
  NAND2_X1 U65256 ( .A1(n106347), .A2(n109897), .ZN(n80145) );
  OAI21_X1 U65257 ( .B1(n106787), .B2(n104735), .A(n80147), .ZN(n103953) );
  NAND2_X1 U65258 ( .A1(n66263), .A2(n106346), .ZN(n80147) );
  OAI21_X1 U65259 ( .B1(n104734), .B2(n106784), .A(n80149), .ZN(n103954) );
  NAND2_X1 U65260 ( .A1(net2411318), .A2(n106346), .ZN(n80149) );
  AOI22_X1 U65261 ( .A1(\DLX_Datapath/next_A_IDEX[30] ), .A2(n80152), .B1(
        n106342), .B2(n108043), .ZN(n80151) );
  AOI22_X1 U65262 ( .A1(\DLX_Datapath/next_A_IDEX[29] ), .A2(n80152), .B1(
        n106342), .B2(n107420), .ZN(n80154) );
  AOI22_X1 U65263 ( .A1(\DLX_Datapath/next_A_IDEX[26] ), .A2(n80152), .B1(
        n106342), .B2(n108152), .ZN(n80155) );
  AOI22_X1 U65264 ( .A1(\DLX_Datapath/next_A_IDEX[25] ), .A2(n80152), .B1(
        n106342), .B2(n110850), .ZN(n80156) );
  AOI22_X1 U65265 ( .A1(\DLX_Datapath/next_A_IDEX[22] ), .A2(n106343), .B1(
        n106342), .B2(n110329), .ZN(n80157) );
  AOI22_X1 U65266 ( .A1(\DLX_Datapath/next_A_IDEX[21] ), .A2(n106344), .B1(
        n106342), .B2(n110649), .ZN(n80158) );
  AOI22_X1 U65267 ( .A1(\DLX_Datapath/next_A_IDEX[20] ), .A2(n106343), .B1(
        n106342), .B2(n110438), .ZN(n80159) );
  AOI22_X1 U65268 ( .A1(\DLX_Datapath/next_A_IDEX[19] ), .A2(n106344), .B1(
        n106342), .B2(n110116), .ZN(n80160) );
  AOI22_X1 U65269 ( .A1(\DLX_Datapath/next_A_IDEX[17] ), .A2(n106344), .B1(
        n106342), .B2(n110008), .ZN(n80161) );
  AOI22_X1 U65270 ( .A1(\DLX_Datapath/next_A_IDEX[15] ), .A2(n106344), .B1(
        n106342), .B2(n108265), .ZN(n80162) );
  AOI22_X1 U65271 ( .A1(\DLX_Datapath/next_A_IDEX[12] ), .A2(n106344), .B1(
        n106342), .B2(n107736), .ZN(n80163) );
  AOI22_X1 U65272 ( .A1(\DLX_Datapath/next_A_IDEX[11] ), .A2(n106344), .B1(
        n106342), .B2(n109651), .ZN(n80164) );
  AOI22_X1 U65273 ( .A1(\DLX_Datapath/next_A_IDEX[8] ), .A2(n106344), .B1(
        n106342), .B2(n109543), .ZN(n80165) );
  AOI22_X1 U65274 ( .A1(\DLX_Datapath/next_A_IDEX[6] ), .A2(n106344), .B1(
        n106342), .B2(n109428), .ZN(n80166) );
  AOI22_X1 U65275 ( .A1(\DLX_Datapath/next_A_IDEX[4] ), .A2(n106344), .B1(
        n106342), .B2(n109201), .ZN(n80167) );
  AOI22_X1 U65276 ( .A1(\DLX_Datapath/next_A_IDEX[2] ), .A2(n106344), .B1(
        n106342), .B2(n108964), .ZN(n80168) );
  AOI22_X1 U65277 ( .A1(\DLX_Datapath/next_A_IDEX[31] ), .A2(n106344), .B1(
        n106342), .B2(n107947), .ZN(n80169) );
  AOI22_X1 U65278 ( .A1(\DLX_Datapath/next_A_IDEX[28] ), .A2(n106344), .B1(
        n106342), .B2(n107852), .ZN(n80170) );
  AOI22_X1 U65279 ( .A1(\DLX_Datapath/next_A_IDEX[27] ), .A2(n106344), .B1(
        n106342), .B2(n110747), .ZN(n80171) );
  AOI22_X1 U65280 ( .A1(\DLX_Datapath/next_A_IDEX[24] ), .A2(n106344), .B1(
        n106342), .B2(n110951), .ZN(n80172) );
  AOI22_X1 U65281 ( .A1(\DLX_Datapath/next_A_IDEX[23] ), .A2(n106343), .B1(
        n106342), .B2(n110544), .ZN(n80173) );
  AOI22_X1 U65282 ( .A1(\DLX_Datapath/next_A_IDEX[18] ), .A2(n106343), .B1(
        n106342), .B2(n110223), .ZN(n80174) );
  AOI22_X1 U65283 ( .A1(\DLX_Datapath/next_A_IDEX[16] ), .A2(n106343), .B1(
        n106342), .B2(n109891), .ZN(n80175) );
  AOI22_X1 U65284 ( .A1(\DLX_Datapath/next_A_IDEX[14] ), .A2(n106343), .B1(
        n106342), .B2(n108388), .ZN(n80176) );
  AOI22_X1 U65285 ( .A1(\DLX_Datapath/next_A_IDEX[13] ), .A2(n106343), .B1(
        n106342), .B2(n108499), .ZN(n80177) );
  AOI22_X1 U65286 ( .A1(\DLX_Datapath/next_A_IDEX[10] ), .A2(n106343), .B1(
        n106342), .B2(n108613), .ZN(n80178) );
  AOI22_X1 U65287 ( .A1(\DLX_Datapath/next_A_IDEX[9] ), .A2(n106343), .B1(
        n106342), .B2(n109758), .ZN(n80179) );
  AOI22_X1 U65288 ( .A1(\DLX_Datapath/next_A_IDEX[7] ), .A2(n106343), .B1(
        n106342), .B2(n109081), .ZN(n80180) );
  AOI22_X1 U65289 ( .A1(\DLX_Datapath/next_A_IDEX[5] ), .A2(n106343), .B1(
        n106342), .B2(n109309), .ZN(n80181) );
  AOI22_X1 U65290 ( .A1(\DLX_Datapath/next_A_IDEX[3] ), .A2(n106343), .B1(
        n106342), .B2(n108736), .ZN(n80182) );
  AOI22_X1 U65291 ( .A1(\DLX_Datapath/next_A_IDEX[1] ), .A2(n106343), .B1(
        n106342), .B2(n108853), .ZN(n80183) );
  AOI22_X1 U65292 ( .A1(\DLX_Datapath/next_A_IDEX[0] ), .A2(n106343), .B1(
        n106342), .B2(n107419), .ZN(n80184) );
  NOR2_X1 U65293 ( .A1(net113155), .A2(n80153), .ZN(n80152) );
  OAI21_X1 U65295 ( .B1(n106341), .B2(n107127), .A(n80186), .ZN(n103955) );
  AOI22_X1 U65296 ( .A1(n106340), .A2(n80188), .B1(n106337), .B2(n108824), 
        .ZN(n80186) );
  OAI21_X1 U65297 ( .B1(n106341), .B2(n80190), .A(n80191), .ZN(n103956) );
  AOI22_X1 U65298 ( .A1(n80192), .A2(n106338), .B1(n106337), .B2(n110516), 
        .ZN(n80191) );
  NAND4_X2 U65299 ( .A1(n80193), .A2(n80194), .A3(n80195), .A4(n80196), .ZN(
        n103957) );
  NOR3_X1 U65300 ( .A1(n80197), .A2(n80198), .A3(n80199), .ZN(n80196) );
  NOR2_X1 U65301 ( .A1(n100613), .A2(n80200), .ZN(n80199) );
  AOI21_X1 U65302 ( .B1(n80201), .B2(n80202), .A(n106326), .ZN(n80198) );
  NOR4_X1 U65303 ( .A1(n80204), .A2(n80205), .A3(n80206), .A4(n80207), .ZN(
        n80202) );
  OAI21_X1 U65304 ( .B1(n106322), .B2(n104616), .A(n80209), .ZN(n80207) );
  AOI22_X1 U65305 ( .A1(n72578), .A2(n80210), .B1(n106320), .B2(n109578), .ZN(
        n80209) );
  NAND2_X1 U65306 ( .A1(n80212), .A2(n80213), .ZN(n80206) );
  AOI22_X1 U65307 ( .A1(n72598), .A2(n80214), .B1(n72586), .B2(n106318), .ZN(
        n80213) );
  AOI22_X1 U65308 ( .A1(n72590), .A2(n80216), .B1(n106316), .B2(n109593), .ZN(
        n80212) );
  NAND2_X1 U65309 ( .A1(n80218), .A2(n80219), .ZN(n80205) );
  AOI22_X1 U65310 ( .A1(n80220), .A2(n109613), .B1(n106314), .B2(n109619), 
        .ZN(n80219) );
  AOI22_X1 U65311 ( .A1(n106313), .A2(n109602), .B1(n80223), .B2(n109607), 
        .ZN(n80218) );
  NAND2_X1 U65312 ( .A1(n80224), .A2(n80225), .ZN(n80204) );
  AOI22_X1 U65313 ( .A1(n80226), .A2(n109622), .B1(n72626), .B2(n106310), .ZN(
        n80225) );
  AOI22_X1 U65314 ( .A1(n80228), .A2(n109610), .B1(n72614), .B2(n106308), .ZN(
        n80224) );
  NOR4_X1 U65315 ( .A1(n80230), .A2(n80231), .A3(n80232), .A4(n80233), .ZN(
        n80201) );
  OAI21_X1 U65316 ( .B1(n101857), .B2(n106307), .A(n80235), .ZN(n80233) );
  AOI22_X1 U65317 ( .A1(n72627), .A2(n80236), .B1(n72639), .B2(n80237), .ZN(
        n80235) );
  NAND2_X1 U65318 ( .A1(n80238), .A2(n80239), .ZN(n80232) );
  AOI22_X1 U65319 ( .A1(n80240), .A2(n109554), .B1(n106303), .B2(n109648), 
        .ZN(n80239) );
  AOI22_X1 U65320 ( .A1(n106302), .A2(n109637), .B1(n80243), .B2(n109645), 
        .ZN(n80238) );
  NAND2_X1 U65321 ( .A1(n80244), .A2(n80245), .ZN(n80231) );
  AOI22_X1 U65322 ( .A1(n80246), .A2(n109561), .B1(n72546), .B2(n80247), .ZN(
        n80245) );
  AOI22_X1 U65323 ( .A1(n106298), .A2(n109565), .B1(n80249), .B2(n109552), 
        .ZN(n80244) );
  NAND2_X1 U65324 ( .A1(n80250), .A2(n80251), .ZN(n80230) );
  AOI22_X1 U65325 ( .A1(n106296), .A2(n109584), .B1(n106295), .B2(n109588), 
        .ZN(n80251) );
  AOI22_X1 U65326 ( .A1(n80254), .A2(n109573), .B1(n72558), .B2(n106293), .ZN(
        n80250) );
  NOR2_X1 U65327 ( .A1(n100581), .A2(n80256), .ZN(n80197) );
  AOI22_X1 U65328 ( .A1(n80257), .A2(n109629), .B1(n80258), .B2(n109641), .ZN(
        n80195) );
  AOI22_X1 U65329 ( .A1(n106746), .A2(n72598), .B1(n105172), .B2(n72614), .ZN(
        n80194) );
  AOI22_X1 U65330 ( .A1(n106289), .A2(n109593), .B1(n106282), .B2(n72566), 
        .ZN(n80193) );
  NAND4_X2 U65331 ( .A1(n80261), .A2(n80262), .A3(n80263), .A4(n80264), .ZN(
        n103958) );
  NOR3_X1 U65332 ( .A1(n80265), .A2(n80266), .A3(n80267), .ZN(n80264) );
  NOR2_X1 U65333 ( .A1(n100614), .A2(n106329), .ZN(n80267) );
  AOI21_X1 U65334 ( .B1(n80268), .B2(n80269), .A(n80203), .ZN(n80266) );
  NOR4_X1 U65335 ( .A1(n80270), .A2(n80271), .A3(n80272), .A4(n80273), .ZN(
        n80269) );
  OAI21_X1 U65336 ( .B1(n80208), .B2(n104647), .A(n80274), .ZN(n80273) );
  AOI22_X1 U65337 ( .A1(n71237), .A2(n80210), .B1(n106320), .B2(n108539), .ZN(
        n80274) );
  NAND2_X1 U65338 ( .A1(n80275), .A2(n80276), .ZN(n80272) );
  AOI22_X1 U65339 ( .A1(n71257), .A2(n80214), .B1(n71245), .B2(n106318), .ZN(
        n80276) );
  AOI22_X1 U65340 ( .A1(n71249), .A2(n80216), .B1(n106316), .B2(n108554), .ZN(
        n80275) );
  NAND2_X1 U65341 ( .A1(n80277), .A2(n80278), .ZN(n80271) );
  AOI22_X1 U65342 ( .A1(n80220), .A2(n108575), .B1(n106314), .B2(n108581), 
        .ZN(n80278) );
  AOI22_X1 U65343 ( .A1(n106313), .A2(n108563), .B1(n80223), .B2(n108569), 
        .ZN(n80277) );
  NAND2_X1 U65344 ( .A1(n80279), .A2(n80280), .ZN(n80270) );
  AOI22_X1 U65345 ( .A1(n80226), .A2(n108584), .B1(n71285), .B2(n106310), .ZN(
        n80280) );
  AOI22_X1 U65346 ( .A1(n80228), .A2(n108572), .B1(n71273), .B2(n106308), .ZN(
        n80279) );
  NOR4_X1 U65347 ( .A1(n80281), .A2(n80282), .A3(n80283), .A4(n80284), .ZN(
        n80268) );
  OAI21_X1 U65348 ( .B1(n101841), .B2(n80234), .A(n80285), .ZN(n80284) );
  AOI22_X1 U65349 ( .A1(n71286), .A2(n80236), .B1(n71298), .B2(n80237), .ZN(
        n80285) );
  NAND2_X1 U65350 ( .A1(n80286), .A2(n80287), .ZN(n80283) );
  AOI22_X1 U65351 ( .A1(n80240), .A2(n108515), .B1(n106303), .B2(n108610), 
        .ZN(n80287) );
  AOI22_X1 U65352 ( .A1(n106302), .A2(n108599), .B1(n80243), .B2(n108607), 
        .ZN(n80286) );
  NAND2_X1 U65353 ( .A1(n80288), .A2(n80289), .ZN(n80282) );
  AOI22_X1 U65354 ( .A1(n80246), .A2(n108522), .B1(n71205), .B2(n80247), .ZN(
        n80289) );
  AOI22_X1 U65355 ( .A1(n106298), .A2(n108526), .B1(n80249), .B2(n108513), 
        .ZN(n80288) );
  NAND2_X1 U65356 ( .A1(n80290), .A2(n80291), .ZN(n80281) );
  AOI22_X1 U65357 ( .A1(n106296), .A2(n108545), .B1(n106295), .B2(n108549), 
        .ZN(n80291) );
  AOI22_X1 U65358 ( .A1(n80254), .A2(n108534), .B1(n71217), .B2(n106293), .ZN(
        n80290) );
  NOR2_X1 U65359 ( .A1(n100582), .A2(n106292), .ZN(n80265) );
  AOI22_X1 U65360 ( .A1(n80257), .A2(n108591), .B1(n80258), .B2(n108603), .ZN(
        n80263) );
  AOI22_X1 U65361 ( .A1(n71257), .A2(n105175), .B1(n71273), .B2(n105172), .ZN(
        n80262) );
  AOI22_X1 U65362 ( .A1(n106289), .A2(n108554), .B1(n71225), .B2(n106283), 
        .ZN(n80261) );
  NAND4_X2 U65363 ( .A1(n80292), .A2(n80293), .A3(n80294), .A4(n80295), .ZN(
        n103959) );
  NOR3_X1 U65364 ( .A1(n80296), .A2(n80297), .A3(n80298), .ZN(n80295) );
  NOR2_X1 U65365 ( .A1(n100615), .A2(n80200), .ZN(n80298) );
  AOI21_X1 U65366 ( .B1(n80299), .B2(n80300), .A(n80203), .ZN(n80297) );
  NOR4_X1 U65367 ( .A1(n80301), .A2(n80302), .A3(n80303), .A4(n80304), .ZN(
        n80300) );
  OAI21_X1 U65368 ( .B1(n106322), .B2(n104646), .A(n80305), .ZN(n80304) );
  AOI22_X1 U65369 ( .A1(n72720), .A2(n80210), .B1(n106320), .B2(n109683), .ZN(
        n80305) );
  NAND2_X1 U65370 ( .A1(n80306), .A2(n80307), .ZN(n80303) );
  AOI22_X1 U65371 ( .A1(n72740), .A2(n80214), .B1(n72728), .B2(n106318), .ZN(
        n80307) );
  AOI22_X1 U65372 ( .A1(n72732), .A2(n80216), .B1(n106316), .B2(n109698), .ZN(
        n80306) );
  NAND2_X1 U65373 ( .A1(n80308), .A2(n80309), .ZN(n80302) );
  AOI22_X1 U65374 ( .A1(n80220), .A2(n109720), .B1(n106314), .B2(n109726), 
        .ZN(n80309) );
  AOI22_X1 U65375 ( .A1(n106313), .A2(n109707), .B1(n80223), .B2(n109713), 
        .ZN(n80308) );
  NAND2_X1 U65376 ( .A1(n80310), .A2(n80311), .ZN(n80301) );
  AOI22_X1 U65377 ( .A1(n80226), .A2(n109729), .B1(n72768), .B2(n106310), .ZN(
        n80311) );
  AOI22_X1 U65378 ( .A1(n80228), .A2(n109716), .B1(n72756), .B2(n106308), .ZN(
        n80310) );
  NOR4_X1 U65379 ( .A1(n80312), .A2(n80313), .A3(n80314), .A4(n80315), .ZN(
        n80299) );
  OAI21_X1 U65380 ( .B1(n101823), .B2(n106307), .A(n80316), .ZN(n80315) );
  AOI22_X1 U65381 ( .A1(n72769), .A2(n80236), .B1(n72781), .B2(n80237), .ZN(
        n80316) );
  NAND2_X1 U65382 ( .A1(n80317), .A2(n80318), .ZN(n80314) );
  AOI22_X1 U65383 ( .A1(n80240), .A2(n109659), .B1(n106303), .B2(n109755), 
        .ZN(n80318) );
  AOI22_X1 U65384 ( .A1(n106302), .A2(n109744), .B1(n80243), .B2(n109752), 
        .ZN(n80317) );
  NAND2_X1 U65385 ( .A1(n80319), .A2(n80320), .ZN(n80313) );
  AOI22_X1 U65386 ( .A1(n80246), .A2(n109666), .B1(n72688), .B2(n80247), .ZN(
        n80320) );
  AOI22_X1 U65387 ( .A1(n106298), .A2(n109670), .B1(n80249), .B2(n109657), 
        .ZN(n80319) );
  NAND2_X1 U65388 ( .A1(n80321), .A2(n80322), .ZN(n80312) );
  AOI22_X1 U65389 ( .A1(n106296), .A2(n109689), .B1(n106295), .B2(n109693), 
        .ZN(n80322) );
  AOI22_X1 U65390 ( .A1(n80254), .A2(n109678), .B1(n72700), .B2(n106293), .ZN(
        n80321) );
  NOR2_X1 U65391 ( .A1(n100583), .A2(n80256), .ZN(n80296) );
  AOI22_X1 U65392 ( .A1(n80257), .A2(n109736), .B1(n80258), .B2(n109748), .ZN(
        n80294) );
  AOI22_X1 U65393 ( .A1(n72740), .A2(n105173), .B1(n72756), .B2(n105172), .ZN(
        n80293) );
  AOI22_X1 U65394 ( .A1(n80259), .A2(n109698), .B1(n72708), .B2(n106285), .ZN(
        n80292) );
  NAND4_X2 U65395 ( .A1(n80323), .A2(n80324), .A3(n80325), .A4(n80326), .ZN(
        n103960) );
  NOR3_X1 U65396 ( .A1(n80327), .A2(n80328), .A3(n80329), .ZN(n80326) );
  NOR2_X1 U65397 ( .A1(n100616), .A2(n106329), .ZN(n80329) );
  AOI21_X1 U65398 ( .B1(n80330), .B2(n80331), .A(n106323), .ZN(n80328) );
  NOR4_X1 U65399 ( .A1(n80332), .A2(n80333), .A3(n80334), .A4(n80335), .ZN(
        n80331) );
  OAI21_X1 U65400 ( .B1(n80208), .B2(n104645), .A(n80336), .ZN(n80335) );
  AOI22_X1 U65401 ( .A1(n72430), .A2(n80210), .B1(n106320), .B2(n109467), .ZN(
        n80336) );
  NAND2_X1 U65402 ( .A1(n80337), .A2(n80338), .ZN(n80334) );
  AOI22_X1 U65403 ( .A1(n72450), .A2(n80214), .B1(n72438), .B2(n106318), .ZN(
        n80338) );
  AOI22_X1 U65404 ( .A1(n72442), .A2(n80216), .B1(n106316), .B2(n109482), .ZN(
        n80337) );
  NAND2_X1 U65405 ( .A1(n80339), .A2(n80340), .ZN(n80333) );
  AOI22_X1 U65406 ( .A1(n80220), .A2(n109505), .B1(n106314), .B2(n109511), 
        .ZN(n80340) );
  AOI22_X1 U65407 ( .A1(n106313), .A2(n109491), .B1(n80223), .B2(n109497), 
        .ZN(n80339) );
  NAND2_X1 U65408 ( .A1(n80341), .A2(n80342), .ZN(n80332) );
  AOI22_X1 U65409 ( .A1(n80226), .A2(n109514), .B1(n72478), .B2(n106310), .ZN(
        n80342) );
  AOI22_X1 U65410 ( .A1(n80228), .A2(n109501), .B1(n72466), .B2(n106308), .ZN(
        n80341) );
  NOR4_X1 U65411 ( .A1(n80343), .A2(n80344), .A3(n80345), .A4(n80346), .ZN(
        n80330) );
  OAI21_X1 U65412 ( .B1(n101805), .B2(n80234), .A(n80347), .ZN(n80346) );
  AOI22_X1 U65413 ( .A1(n72479), .A2(n80236), .B1(n72491), .B2(n80237), .ZN(
        n80347) );
  NAND2_X1 U65414 ( .A1(n80348), .A2(n80349), .ZN(n80345) );
  AOI22_X1 U65415 ( .A1(n80240), .A2(n109443), .B1(n106303), .B2(n109540), 
        .ZN(n80349) );
  AOI22_X1 U65416 ( .A1(n106302), .A2(n109529), .B1(n80243), .B2(n109537), 
        .ZN(n80348) );
  NAND2_X1 U65417 ( .A1(n80350), .A2(n80351), .ZN(n80344) );
  AOI22_X1 U65418 ( .A1(n80246), .A2(n109450), .B1(n72398), .B2(n80247), .ZN(
        n80351) );
  AOI22_X1 U65419 ( .A1(n106298), .A2(n109454), .B1(n80249), .B2(n109441), 
        .ZN(n80350) );
  NAND2_X1 U65420 ( .A1(n80352), .A2(n80353), .ZN(n80343) );
  AOI22_X1 U65421 ( .A1(n106296), .A2(n109473), .B1(n106295), .B2(n109477), 
        .ZN(n80353) );
  AOI22_X1 U65422 ( .A1(n80254), .A2(n109462), .B1(n72410), .B2(n106293), .ZN(
        n80352) );
  NOR2_X1 U65423 ( .A1(n100584), .A2(n106292), .ZN(n80327) );
  AOI22_X1 U65424 ( .A1(n80257), .A2(n109521), .B1(n80258), .B2(n109533), .ZN(
        n80325) );
  AOI22_X1 U65425 ( .A1(n72450), .A2(n105174), .B1(n72466), .B2(n105172), .ZN(
        n80324) );
  AOI22_X1 U65426 ( .A1(n80259), .A2(n109482), .B1(n72418), .B2(n106284), .ZN(
        n80323) );
  NAND4_X2 U65427 ( .A1(n80354), .A2(n80355), .A3(n80356), .A4(n80357), .ZN(
        n103961) );
  NOR3_X1 U65428 ( .A1(n80358), .A2(n80359), .A3(n80360), .ZN(n80357) );
  NOR2_X1 U65429 ( .A1(n100617), .A2(n80200), .ZN(n80360) );
  AOI21_X1 U65430 ( .B1(n80361), .B2(n80362), .A(n80203), .ZN(n80359) );
  NOR4_X1 U65431 ( .A1(n80363), .A2(n80364), .A3(n80365), .A4(n80366), .ZN(
        n80362) );
  OAI21_X1 U65432 ( .B1(n106322), .B2(n104644), .A(n80367), .ZN(n80366) );
  AOI22_X1 U65433 ( .A1(n71830), .A2(n80210), .B1(n106320), .B2(n109004), .ZN(
        n80367) );
  NAND2_X1 U65434 ( .A1(n80368), .A2(n80369), .ZN(n80365) );
  AOI22_X1 U65435 ( .A1(n71850), .A2(n80214), .B1(n71838), .B2(n106318), .ZN(
        n80369) );
  AOI22_X1 U65436 ( .A1(n71842), .A2(n80216), .B1(n106316), .B2(n109019), .ZN(
        n80368) );
  NAND2_X1 U65437 ( .A1(n80370), .A2(n80371), .ZN(n80364) );
  AOI22_X1 U65438 ( .A1(n80220), .A2(n109042), .B1(n106314), .B2(n109048), 
        .ZN(n80371) );
  AOI22_X1 U65439 ( .A1(n106313), .A2(n109028), .B1(n80223), .B2(n109034), 
        .ZN(n80370) );
  NAND2_X1 U65440 ( .A1(n80372), .A2(n80373), .ZN(n80363) );
  AOI22_X1 U65441 ( .A1(n80226), .A2(n109051), .B1(n71878), .B2(n106310), .ZN(
        n80373) );
  AOI22_X1 U65442 ( .A1(n80228), .A2(n109038), .B1(n71866), .B2(n106308), .ZN(
        n80372) );
  NOR4_X1 U65443 ( .A1(n80374), .A2(n80375), .A3(n80376), .A4(n80377), .ZN(
        n80361) );
  OAI21_X1 U65444 ( .B1(n101789), .B2(n106307), .A(n80378), .ZN(n80377) );
  AOI22_X1 U65445 ( .A1(n71879), .A2(n80236), .B1(n71891), .B2(n80237), .ZN(
        n80378) );
  NAND2_X1 U65446 ( .A1(n80379), .A2(n80380), .ZN(n80376) );
  AOI22_X1 U65447 ( .A1(n80240), .A2(n108980), .B1(n106303), .B2(n109078), 
        .ZN(n80380) );
  AOI22_X1 U65448 ( .A1(n106302), .A2(n109067), .B1(n80243), .B2(n109075), 
        .ZN(n80379) );
  NAND2_X1 U65449 ( .A1(n80381), .A2(n80382), .ZN(n80375) );
  AOI22_X1 U65450 ( .A1(n80246), .A2(n108987), .B1(n71798), .B2(n80247), .ZN(
        n80382) );
  AOI22_X1 U65451 ( .A1(n106298), .A2(n108991), .B1(n80249), .B2(n108978), 
        .ZN(n80381) );
  NAND2_X1 U65452 ( .A1(n80383), .A2(n80384), .ZN(n80374) );
  AOI22_X1 U65453 ( .A1(n106296), .A2(n109010), .B1(n106295), .B2(n109014), 
        .ZN(n80384) );
  AOI22_X1 U65454 ( .A1(n80254), .A2(n108999), .B1(n71810), .B2(n106293), .ZN(
        n80383) );
  NOR2_X1 U65455 ( .A1(n100585), .A2(n80256), .ZN(n80358) );
  AOI22_X1 U65456 ( .A1(n80257), .A2(n109059), .B1(n80258), .B2(n109071), .ZN(
        n80356) );
  AOI22_X1 U65457 ( .A1(n71850), .A2(n106746), .B1(n71866), .B2(n105172), .ZN(
        n80355) );
  AOI22_X1 U65458 ( .A1(n106286), .A2(n109019), .B1(n71818), .B2(n106282), 
        .ZN(n80354) );
  NAND4_X2 U65459 ( .A1(n80385), .A2(n80386), .A3(n80387), .A4(n80388), .ZN(
        n103962) );
  NOR3_X1 U65460 ( .A1(n80389), .A2(n80390), .A3(n80391), .ZN(n80388) );
  NOR2_X1 U65461 ( .A1(n100618), .A2(n106329), .ZN(n80391) );
  AOI21_X1 U65462 ( .B1(n80392), .B2(n80393), .A(n80203), .ZN(n80390) );
  NOR4_X1 U65463 ( .A1(n80394), .A2(n80395), .A3(n80396), .A4(n80397), .ZN(
        n80393) );
  OAI21_X1 U65464 ( .B1(n80208), .B2(n104643), .A(n80398), .ZN(n80397) );
  AOI22_X1 U65465 ( .A1(n72279), .A2(n80210), .B1(n106320), .B2(n109352), .ZN(
        n80398) );
  NAND2_X1 U65466 ( .A1(n80399), .A2(n80400), .ZN(n80396) );
  AOI22_X1 U65467 ( .A1(n72299), .A2(n80214), .B1(n72287), .B2(n106318), .ZN(
        n80400) );
  AOI22_X1 U65468 ( .A1(n72291), .A2(n80216), .B1(n106316), .B2(n109367), .ZN(
        n80399) );
  NAND2_X1 U65469 ( .A1(n80401), .A2(n80402), .ZN(n80395) );
  AOI22_X1 U65470 ( .A1(n80220), .A2(n109390), .B1(n106314), .B2(n109396), 
        .ZN(n80402) );
  AOI22_X1 U65471 ( .A1(n106313), .A2(n109376), .B1(n80223), .B2(n109382), 
        .ZN(n80401) );
  NAND2_X1 U65472 ( .A1(n80403), .A2(n80404), .ZN(n80394) );
  AOI22_X1 U65473 ( .A1(n80226), .A2(n109399), .B1(n72327), .B2(n106310), .ZN(
        n80404) );
  AOI22_X1 U65474 ( .A1(n80228), .A2(n109386), .B1(n72315), .B2(n106308), .ZN(
        n80403) );
  NOR4_X1 U65475 ( .A1(n80405), .A2(n80406), .A3(n80407), .A4(n80408), .ZN(
        n80392) );
  OAI21_X1 U65476 ( .B1(n101771), .B2(n80234), .A(n80409), .ZN(n80408) );
  AOI22_X1 U65477 ( .A1(n72328), .A2(n80236), .B1(n72340), .B2(n80237), .ZN(
        n80409) );
  NAND2_X1 U65478 ( .A1(n80410), .A2(n80411), .ZN(n80407) );
  AOI22_X1 U65479 ( .A1(n80240), .A2(n109328), .B1(n106303), .B2(n109425), 
        .ZN(n80411) );
  AOI22_X1 U65480 ( .A1(n106302), .A2(n109414), .B1(n80243), .B2(n109422), 
        .ZN(n80410) );
  NAND2_X1 U65481 ( .A1(n80412), .A2(n80413), .ZN(n80406) );
  AOI22_X1 U65482 ( .A1(n80246), .A2(n109335), .B1(n72247), .B2(n80247), .ZN(
        n80413) );
  AOI22_X1 U65483 ( .A1(n106298), .A2(n109339), .B1(n80249), .B2(n109326), 
        .ZN(n80412) );
  NAND2_X1 U65484 ( .A1(n80414), .A2(n80415), .ZN(n80405) );
  AOI22_X1 U65485 ( .A1(n106296), .A2(n109358), .B1(n106295), .B2(n109362), 
        .ZN(n80415) );
  AOI22_X1 U65486 ( .A1(n80254), .A2(n109347), .B1(n72259), .B2(n106293), .ZN(
        n80414) );
  NOR2_X1 U65487 ( .A1(n100586), .A2(n106292), .ZN(n80389) );
  AOI22_X1 U65488 ( .A1(n80257), .A2(n109406), .B1(n80258), .B2(n109418), .ZN(
        n80387) );
  AOI22_X1 U65489 ( .A1(n72299), .A2(n105175), .B1(n72315), .B2(n105172), .ZN(
        n80386) );
  AOI22_X1 U65490 ( .A1(n106286), .A2(n109367), .B1(n72267), .B2(n106283), 
        .ZN(n80385) );
  NAND4_X2 U65491 ( .A1(n80416), .A2(n80417), .A3(n80418), .A4(n80419), .ZN(
        n103963) );
  NOR3_X1 U65492 ( .A1(n80420), .A2(n80421), .A3(n80422), .ZN(n80419) );
  NOR2_X1 U65493 ( .A1(n100619), .A2(n80200), .ZN(n80422) );
  AOI21_X1 U65494 ( .B1(n80423), .B2(n80424), .A(n106323), .ZN(n80421) );
  NOR4_X1 U65495 ( .A1(n80425), .A2(n80426), .A3(n80427), .A4(n80428), .ZN(
        n80424) );
  OAI21_X1 U65496 ( .B1(n106322), .B2(n104642), .A(n80429), .ZN(n80428) );
  AOI22_X1 U65497 ( .A1(n72128), .A2(n80210), .B1(n106320), .B2(n109234), .ZN(
        n80429) );
  NAND2_X1 U65498 ( .A1(n80430), .A2(n80431), .ZN(n80427) );
  AOI22_X1 U65499 ( .A1(n72148), .A2(n80214), .B1(n72136), .B2(n106318), .ZN(
        n80431) );
  AOI22_X1 U65500 ( .A1(n72140), .A2(n80216), .B1(n106316), .B2(n109249), .ZN(
        n80430) );
  NAND2_X1 U65501 ( .A1(n80432), .A2(n80433), .ZN(n80426) );
  AOI22_X1 U65502 ( .A1(n80220), .A2(n109272), .B1(n106314), .B2(n109278), 
        .ZN(n80433) );
  AOI22_X1 U65503 ( .A1(n106313), .A2(n109258), .B1(n80223), .B2(n109264), 
        .ZN(n80432) );
  NAND2_X1 U65504 ( .A1(n80434), .A2(n80435), .ZN(n80425) );
  AOI22_X1 U65505 ( .A1(n80226), .A2(n109280), .B1(n72176), .B2(n106310), .ZN(
        n80435) );
  AOI22_X1 U65506 ( .A1(n80228), .A2(n109268), .B1(n72164), .B2(n106308), .ZN(
        n80434) );
  NOR4_X1 U65507 ( .A1(n80436), .A2(n80437), .A3(n80438), .A4(n80439), .ZN(
        n80423) );
  OAI21_X1 U65508 ( .B1(n101755), .B2(n106307), .A(n80440), .ZN(n80439) );
  AOI22_X1 U65509 ( .A1(n72177), .A2(n80236), .B1(n72189), .B2(n80237), .ZN(
        n80440) );
  NAND2_X1 U65510 ( .A1(n80441), .A2(n80442), .ZN(n80438) );
  AOI22_X1 U65511 ( .A1(n80240), .A2(n109210), .B1(n106303), .B2(n109306), 
        .ZN(n80442) );
  AOI22_X1 U65512 ( .A1(n106302), .A2(n109295), .B1(n80243), .B2(n109303), 
        .ZN(n80441) );
  NAND2_X1 U65513 ( .A1(n80443), .A2(n80444), .ZN(n80437) );
  AOI22_X1 U65514 ( .A1(n80246), .A2(n109217), .B1(n72096), .B2(n80247), .ZN(
        n80444) );
  AOI22_X1 U65515 ( .A1(n106298), .A2(n109221), .B1(n80249), .B2(n109208), 
        .ZN(n80443) );
  NAND2_X1 U65516 ( .A1(n80445), .A2(n80446), .ZN(n80436) );
  AOI22_X1 U65517 ( .A1(n106296), .A2(n109240), .B1(n106295), .B2(n109244), 
        .ZN(n80446) );
  AOI22_X1 U65518 ( .A1(n80254), .A2(n109229), .B1(n72108), .B2(n106293), .ZN(
        n80445) );
  NOR2_X1 U65519 ( .A1(n100587), .A2(n80256), .ZN(n80420) );
  AOI22_X1 U65520 ( .A1(n80257), .A2(n109287), .B1(n80258), .B2(n109299), .ZN(
        n80418) );
  AOI22_X1 U65521 ( .A1(n72148), .A2(n105174), .B1(n72164), .B2(n105172), .ZN(
        n80417) );
  AOI22_X1 U65522 ( .A1(n106286), .A2(n109249), .B1(n72116), .B2(n106283), 
        .ZN(n80416) );
  NAND4_X2 U65523 ( .A1(n80447), .A2(n80448), .A3(n80449), .A4(n80450), .ZN(
        n103964) );
  NOR3_X1 U65524 ( .A1(n80451), .A2(n80452), .A3(n80453), .ZN(n80450) );
  NOR2_X1 U65525 ( .A1(n100620), .A2(n106329), .ZN(n80453) );
  AOI21_X1 U65526 ( .B1(n80454), .B2(n80455), .A(n106323), .ZN(n80452) );
  NOR4_X1 U65527 ( .A1(n80456), .A2(n80457), .A3(n80458), .A4(n80459), .ZN(
        n80455) );
  OAI21_X1 U65528 ( .B1(n80208), .B2(n104641), .A(n80460), .ZN(n80459) );
  AOI22_X1 U65529 ( .A1(n71984), .A2(n80210), .B1(n106320), .B2(n109126), .ZN(
        n80460) );
  NAND2_X1 U65530 ( .A1(n80461), .A2(n80462), .ZN(n80458) );
  AOI22_X1 U65531 ( .A1(n72004), .A2(n80214), .B1(n71992), .B2(n106318), .ZN(
        n80462) );
  AOI22_X1 U65532 ( .A1(n71996), .A2(n80216), .B1(n106316), .B2(n109141), .ZN(
        n80461) );
  NAND2_X1 U65533 ( .A1(n80463), .A2(n80464), .ZN(n80457) );
  AOI22_X1 U65534 ( .A1(n80220), .A2(n109163), .B1(n106314), .B2(n109169), 
        .ZN(n80464) );
  AOI22_X1 U65535 ( .A1(n106313), .A2(n109149), .B1(n80223), .B2(n109155), 
        .ZN(n80463) );
  NAND2_X1 U65536 ( .A1(n80465), .A2(n80466), .ZN(n80456) );
  AOI22_X1 U65537 ( .A1(n80226), .A2(n109172), .B1(n72032), .B2(n106310), .ZN(
        n80466) );
  AOI22_X1 U65538 ( .A1(n80228), .A2(n109159), .B1(n72020), .B2(n106308), .ZN(
        n80465) );
  NOR4_X1 U65539 ( .A1(n80467), .A2(n80468), .A3(n80469), .A4(n80470), .ZN(
        n80454) );
  OAI21_X1 U65540 ( .B1(n101737), .B2(n80234), .A(n80471), .ZN(n80470) );
  AOI22_X1 U65541 ( .A1(n72033), .A2(n80236), .B1(n72045), .B2(n80237), .ZN(
        n80471) );
  NAND2_X1 U65542 ( .A1(n80472), .A2(n80473), .ZN(n80469) );
  AOI22_X1 U65543 ( .A1(n80240), .A2(n109102), .B1(n106303), .B2(n109198), 
        .ZN(n80473) );
  AOI22_X1 U65544 ( .A1(n106302), .A2(n109187), .B1(n80243), .B2(n109195), 
        .ZN(n80472) );
  NAND2_X1 U65545 ( .A1(n80474), .A2(n80475), .ZN(n80468) );
  AOI22_X1 U65546 ( .A1(n80246), .A2(n109109), .B1(n71952), .B2(n80247), .ZN(
        n80475) );
  AOI22_X1 U65547 ( .A1(n106298), .A2(n109113), .B1(n80249), .B2(n109100), 
        .ZN(n80474) );
  NAND2_X1 U65548 ( .A1(n80476), .A2(n80477), .ZN(n80467) );
  AOI22_X1 U65549 ( .A1(n106296), .A2(n109132), .B1(n106295), .B2(n109136), 
        .ZN(n80477) );
  AOI22_X1 U65550 ( .A1(n80254), .A2(n109121), .B1(n71964), .B2(n106293), .ZN(
        n80476) );
  NOR2_X1 U65551 ( .A1(n100588), .A2(n106292), .ZN(n80451) );
  AOI22_X1 U65552 ( .A1(n80257), .A2(n109179), .B1(n80258), .B2(n109191), .ZN(
        n80449) );
  AOI22_X1 U65553 ( .A1(n72004), .A2(n105173), .B1(n72020), .B2(n105172), .ZN(
        n80448) );
  AOI22_X1 U65554 ( .A1(n106286), .A2(n109141), .B1(n71972), .B2(n106284), 
        .ZN(n80447) );
  NAND4_X2 U65555 ( .A1(n80478), .A2(n80479), .A3(n80480), .A4(n80481), .ZN(
        n103965) );
  NOR3_X1 U65556 ( .A1(n80482), .A2(n80483), .A3(n80484), .ZN(n80481) );
  NOR2_X1 U65557 ( .A1(n100621), .A2(n106329), .ZN(n80484) );
  AOI21_X1 U65558 ( .B1(n80485), .B2(n80486), .A(n106324), .ZN(n80483) );
  NOR4_X1 U65559 ( .A1(n80487), .A2(n80488), .A3(n80489), .A4(n80490), .ZN(
        n80486) );
  OAI21_X1 U65560 ( .B1(n106322), .B2(n104640), .A(n80491), .ZN(n80490) );
  AOI22_X1 U65561 ( .A1(n71386), .A2(n80210), .B1(n106320), .B2(n108661), .ZN(
        n80491) );
  NAND2_X1 U65562 ( .A1(n80492), .A2(n80493), .ZN(n80489) );
  AOI22_X1 U65563 ( .A1(n71406), .A2(n80214), .B1(n71394), .B2(n106318), .ZN(
        n80493) );
  AOI22_X1 U65564 ( .A1(n71398), .A2(n80216), .B1(n106316), .B2(n108676), .ZN(
        n80492) );
  NAND2_X1 U65565 ( .A1(n80494), .A2(n80495), .ZN(n80488) );
  AOI22_X1 U65566 ( .A1(n80220), .A2(n108699), .B1(n80221), .B2(n108705), .ZN(
        n80495) );
  AOI22_X1 U65567 ( .A1(n80222), .A2(n108685), .B1(n106312), .B2(n108691), 
        .ZN(n80494) );
  NAND2_X1 U65568 ( .A1(n80496), .A2(n80497), .ZN(n80487) );
  AOI22_X1 U65569 ( .A1(n80226), .A2(n108707), .B1(n71434), .B2(n80227), .ZN(
        n80497) );
  AOI22_X1 U65570 ( .A1(n80228), .A2(n108695), .B1(n71422), .B2(n106308), .ZN(
        n80496) );
  NOR4_X1 U65571 ( .A1(n80498), .A2(n80499), .A3(n80500), .A4(n80501), .ZN(
        n80485) );
  OAI21_X1 U65572 ( .B1(n101719), .B2(n106307), .A(n80502), .ZN(n80501) );
  AOI22_X1 U65573 ( .A1(n71435), .A2(n80236), .B1(n71447), .B2(n80237), .ZN(
        n80502) );
  NAND2_X1 U65574 ( .A1(n80503), .A2(n80504), .ZN(n80500) );
  AOI22_X1 U65575 ( .A1(n80240), .A2(n108637), .B1(n80241), .B2(n108733), .ZN(
        n80504) );
  AOI22_X1 U65576 ( .A1(n106302), .A2(n108722), .B1(n80243), .B2(n108730), 
        .ZN(n80503) );
  NAND2_X1 U65577 ( .A1(n80505), .A2(n80506), .ZN(n80499) );
  AOI22_X1 U65578 ( .A1(n80246), .A2(n108644), .B1(n71354), .B2(n80247), .ZN(
        n80506) );
  AOI22_X1 U65579 ( .A1(n80248), .A2(n108648), .B1(n80249), .B2(n108635), .ZN(
        n80505) );
  NAND2_X1 U65580 ( .A1(n80507), .A2(n80508), .ZN(n80498) );
  AOI22_X1 U65581 ( .A1(n106296), .A2(n108667), .B1(n106295), .B2(n108671), 
        .ZN(n80508) );
  AOI22_X1 U65582 ( .A1(n80254), .A2(n108656), .B1(n71366), .B2(n80255), .ZN(
        n80507) );
  NOR2_X1 U65583 ( .A1(n100589), .A2(n106292), .ZN(n80482) );
  AOI22_X1 U65584 ( .A1(n80257), .A2(n108714), .B1(n80258), .B2(n108726), .ZN(
        n80480) );
  AOI22_X1 U65585 ( .A1(n71406), .A2(n105174), .B1(n71422), .B2(n105172), .ZN(
        n80479) );
  AOI22_X1 U65586 ( .A1(n106286), .A2(n108676), .B1(n71374), .B2(n80260), .ZN(
        n80478) );
  NAND4_X2 U65587 ( .A1(n80509), .A2(n80510), .A3(n80511), .A4(n80512), .ZN(
        n103966) );
  NOR3_X1 U65588 ( .A1(n80513), .A2(n80514), .A3(n80515), .ZN(n80512) );
  NOR2_X1 U65589 ( .A1(n100622), .A2(n80200), .ZN(n80515) );
  AOI21_X1 U65590 ( .B1(n80516), .B2(n80517), .A(n106325), .ZN(n80514) );
  NOR4_X1 U65591 ( .A1(n80518), .A2(n80519), .A3(n80520), .A4(n80521), .ZN(
        n80517) );
  OAI21_X1 U65592 ( .B1(n106322), .B2(n104639), .A(n80522), .ZN(n80521) );
  AOI22_X1 U65593 ( .A1(n71681), .A2(n80210), .B1(n106320), .B2(n108888), .ZN(
        n80522) );
  NAND2_X1 U65594 ( .A1(n80523), .A2(n80524), .ZN(n80520) );
  AOI22_X1 U65595 ( .A1(n71701), .A2(n80214), .B1(n71689), .B2(n106318), .ZN(
        n80524) );
  AOI22_X1 U65596 ( .A1(n71693), .A2(n80216), .B1(n106316), .B2(n108903), .ZN(
        n80523) );
  NAND2_X1 U65597 ( .A1(n80525), .A2(n80526), .ZN(n80519) );
  AOI22_X1 U65598 ( .A1(n80220), .A2(n108926), .B1(n80221), .B2(n108932), .ZN(
        n80526) );
  AOI22_X1 U65599 ( .A1(n80222), .A2(n108912), .B1(n106312), .B2(n108918), 
        .ZN(n80525) );
  NAND2_X1 U65600 ( .A1(n80527), .A2(n80528), .ZN(n80518) );
  AOI22_X1 U65601 ( .A1(n80226), .A2(n108935), .B1(n71729), .B2(n80227), .ZN(
        n80528) );
  AOI22_X1 U65602 ( .A1(n80228), .A2(n108922), .B1(n71717), .B2(n106308), .ZN(
        n80527) );
  NOR4_X1 U65603 ( .A1(n80529), .A2(n80530), .A3(n80531), .A4(n80532), .ZN(
        n80516) );
  OAI21_X1 U65604 ( .B1(n101701), .B2(n106307), .A(n80533), .ZN(n80532) );
  AOI22_X1 U65605 ( .A1(n71730), .A2(n80236), .B1(n71742), .B2(n80237), .ZN(
        n80533) );
  NAND2_X1 U65606 ( .A1(n80534), .A2(n80535), .ZN(n80531) );
  AOI22_X1 U65607 ( .A1(n80240), .A2(n108864), .B1(n80241), .B2(n108961), .ZN(
        n80535) );
  AOI22_X1 U65608 ( .A1(n106302), .A2(n108950), .B1(n80243), .B2(n108958), 
        .ZN(n80534) );
  NAND2_X1 U65609 ( .A1(n80536), .A2(n80537), .ZN(n80530) );
  AOI22_X1 U65610 ( .A1(n80246), .A2(n108871), .B1(n71649), .B2(n80247), .ZN(
        n80537) );
  AOI22_X1 U65611 ( .A1(n80248), .A2(n108875), .B1(n106297), .B2(n108862), 
        .ZN(n80536) );
  NAND2_X1 U65612 ( .A1(n80538), .A2(n80539), .ZN(n80529) );
  AOI22_X1 U65613 ( .A1(n106296), .A2(n108894), .B1(n106295), .B2(n108898), 
        .ZN(n80539) );
  AOI22_X1 U65614 ( .A1(n80254), .A2(n108883), .B1(n71661), .B2(n80255), .ZN(
        n80538) );
  NOR2_X1 U65615 ( .A1(n100590), .A2(n80256), .ZN(n80513) );
  AOI22_X1 U65616 ( .A1(n80257), .A2(n108942), .B1(n80258), .B2(n108954), .ZN(
        n80511) );
  AOI22_X1 U65617 ( .A1(n71701), .A2(n106746), .B1(n71717), .B2(n105172), .ZN(
        n80510) );
  AOI22_X1 U65618 ( .A1(n106289), .A2(n108903), .B1(n71669), .B2(n106282), 
        .ZN(n80509) );
  NAND4_X2 U65619 ( .A1(n80540), .A2(n80541), .A3(n80542), .A4(n80543), .ZN(
        n103967) );
  NOR3_X1 U65620 ( .A1(n80544), .A2(n80545), .A3(n80546), .ZN(n80543) );
  NOR2_X1 U65621 ( .A1(n100623), .A2(n106329), .ZN(n80546) );
  AOI21_X1 U65622 ( .B1(n80547), .B2(n80548), .A(n106326), .ZN(n80545) );
  NOR4_X1 U65623 ( .A1(n80549), .A2(n80550), .A3(n80551), .A4(n80552), .ZN(
        n80548) );
  OAI21_X1 U65624 ( .B1(n106322), .B2(n104638), .A(n80553), .ZN(n80552) );
  AOI22_X1 U65625 ( .A1(n71537), .A2(n80210), .B1(n106320), .B2(n108776), .ZN(
        n80553) );
  NAND2_X1 U65626 ( .A1(n80554), .A2(n80555), .ZN(n80551) );
  AOI22_X1 U65627 ( .A1(n71557), .A2(n80214), .B1(n71545), .B2(n106318), .ZN(
        n80555) );
  AOI22_X1 U65628 ( .A1(n71549), .A2(n80216), .B1(n106316), .B2(n108791), .ZN(
        n80554) );
  NAND2_X1 U65629 ( .A1(n80556), .A2(n80557), .ZN(n80550) );
  AOI22_X1 U65630 ( .A1(n80220), .A2(n108814), .B1(n106314), .B2(n108820), 
        .ZN(n80557) );
  AOI22_X1 U65631 ( .A1(n106313), .A2(n108800), .B1(n80223), .B2(n108806), 
        .ZN(n80556) );
  NAND2_X1 U65632 ( .A1(n80558), .A2(n80559), .ZN(n80549) );
  AOI22_X1 U65633 ( .A1(n80226), .A2(n108823), .B1(n71585), .B2(n80227), .ZN(
        n80559) );
  AOI22_X1 U65634 ( .A1(n80228), .A2(n108810), .B1(n71573), .B2(n106308), .ZN(
        n80558) );
  NOR4_X1 U65635 ( .A1(n80560), .A2(n80561), .A3(n80562), .A4(n80563), .ZN(
        n80547) );
  OAI21_X1 U65636 ( .B1(n101683), .B2(n106307), .A(n80564), .ZN(n80563) );
  AOI22_X1 U65637 ( .A1(n71586), .A2(n80236), .B1(n71598), .B2(n80237), .ZN(
        n80564) );
  NAND2_X1 U65638 ( .A1(n80565), .A2(n80566), .ZN(n80562) );
  AOI22_X1 U65639 ( .A1(n80240), .A2(n108752), .B1(n80241), .B2(n108849), .ZN(
        n80566) );
  AOI22_X1 U65640 ( .A1(n106302), .A2(n108838), .B1(n80243), .B2(n108846), 
        .ZN(n80565) );
  NAND2_X1 U65641 ( .A1(n80567), .A2(n80568), .ZN(n80561) );
  AOI22_X1 U65642 ( .A1(n80246), .A2(n108759), .B1(n71505), .B2(n80247), .ZN(
        n80568) );
  AOI22_X1 U65643 ( .A1(n80248), .A2(n108763), .B1(n106297), .B2(n108750), 
        .ZN(n80567) );
  NAND2_X1 U65644 ( .A1(n80569), .A2(n80570), .ZN(n80560) );
  AOI22_X1 U65645 ( .A1(n106296), .A2(n108782), .B1(n106295), .B2(n108786), 
        .ZN(n80570) );
  AOI22_X1 U65646 ( .A1(n80254), .A2(n108771), .B1(n71517), .B2(n80255), .ZN(
        n80569) );
  NOR2_X1 U65647 ( .A1(n100591), .A2(n106292), .ZN(n80544) );
  AOI22_X1 U65648 ( .A1(n80257), .A2(n108830), .B1(n80258), .B2(n108842), .ZN(
        n80542) );
  AOI22_X1 U65649 ( .A1(n71557), .A2(n105173), .B1(n71573), .B2(n105172), .ZN(
        n80541) );
  AOI22_X1 U65650 ( .A1(n80259), .A2(n108791), .B1(n71525), .B2(n80260), .ZN(
        n80540) );
  NAND4_X2 U65651 ( .A1(n80571), .A2(n80572), .A3(n80573), .A4(n80574), .ZN(
        n103968) );
  NOR3_X1 U65652 ( .A1(n80575), .A2(n80576), .A3(n80577), .ZN(n80574) );
  NOR2_X1 U65653 ( .A1(n100624), .A2(n80200), .ZN(n80577) );
  AOI21_X1 U65654 ( .B1(n80578), .B2(n80579), .A(n106324), .ZN(n80576) );
  NOR4_X1 U65655 ( .A1(n80580), .A2(n80581), .A3(n80582), .A4(n80583), .ZN(
        n80579) );
  OAI21_X1 U65656 ( .B1(n106322), .B2(n104637), .A(n80584), .ZN(n80583) );
  AOI22_X1 U65657 ( .A1(n69646), .A2(n106321), .B1(n106320), .B2(n107316), 
        .ZN(n80584) );
  NAND2_X1 U65658 ( .A1(n80585), .A2(n80586), .ZN(n80582) );
  AOI22_X1 U65659 ( .A1(n69666), .A2(n106319), .B1(n69654), .B2(n106318), .ZN(
        n80586) );
  AOI22_X1 U65660 ( .A1(n69658), .A2(n106317), .B1(n106316), .B2(n107331), 
        .ZN(n80585) );
  NAND2_X1 U65661 ( .A1(n80587), .A2(n80588), .ZN(n80581) );
  AOI22_X1 U65662 ( .A1(n106315), .A2(n107354), .B1(n106314), .B2(n107360), 
        .ZN(n80588) );
  AOI22_X1 U65663 ( .A1(n106313), .A2(n107340), .B1(n80223), .B2(n107346), 
        .ZN(n80587) );
  NAND2_X1 U65664 ( .A1(n80589), .A2(n80590), .ZN(n80580) );
  AOI22_X1 U65665 ( .A1(n106311), .A2(n107362), .B1(n69694), .B2(n80227), .ZN(
        n80590) );
  AOI22_X1 U65666 ( .A1(n106309), .A2(n107350), .B1(n69682), .B2(n106308), 
        .ZN(n80589) );
  NOR4_X1 U65667 ( .A1(n80591), .A2(n80592), .A3(n80593), .A4(n80594), .ZN(
        n80578) );
  OAI21_X1 U65668 ( .B1(n101665), .B2(n106307), .A(n80595), .ZN(n80594) );
  AOI22_X1 U65669 ( .A1(n69484), .A2(n106306), .B1(n69460), .B2(n106305), .ZN(
        n80595) );
  NAND2_X1 U65670 ( .A1(n80596), .A2(n80597), .ZN(n80593) );
  AOI22_X1 U65671 ( .A1(n106304), .A2(n107292), .B1(n80241), .B2(n107169), 
        .ZN(n80597) );
  AOI22_X1 U65672 ( .A1(n106302), .A2(n107191), .B1(n80243), .B2(n107175), 
        .ZN(n80596) );
  NAND2_X1 U65673 ( .A1(n80598), .A2(n80599), .ZN(n80592) );
  AOI22_X1 U65674 ( .A1(n106300), .A2(n107299), .B1(n69614), .B2(n106299), 
        .ZN(n80599) );
  AOI22_X1 U65675 ( .A1(n80248), .A2(n107303), .B1(n106297), .B2(n107290), 
        .ZN(n80598) );
  NAND2_X1 U65676 ( .A1(n80600), .A2(n80601), .ZN(n80591) );
  AOI22_X1 U65677 ( .A1(n106296), .A2(n107322), .B1(n106295), .B2(n107326), 
        .ZN(n80601) );
  AOI22_X1 U65678 ( .A1(n106294), .A2(n107311), .B1(n69626), .B2(n80255), .ZN(
        n80600) );
  NOR2_X1 U65679 ( .A1(n100592), .A2(n80256), .ZN(n80575) );
  AOI22_X1 U65680 ( .A1(n106291), .A2(n107207), .B1(n106290), .B2(n107183), 
        .ZN(n80573) );
  AOI22_X1 U65681 ( .A1(n69666), .A2(n106746), .B1(n69682), .B2(n105172), .ZN(
        n80572) );
  AOI22_X1 U65682 ( .A1(n106286), .A2(n107331), .B1(n69634), .B2(n106283), 
        .ZN(n80571) );
  NAND4_X2 U65683 ( .A1(n80602), .A2(n80603), .A3(n80604), .A4(n80605), .ZN(
        n103969) );
  NOR3_X1 U65684 ( .A1(n80606), .A2(n80607), .A3(n80608), .ZN(n80605) );
  NOR2_X1 U65685 ( .A1(n100593), .A2(n106329), .ZN(n80608) );
  AOI21_X1 U65686 ( .B1(n80609), .B2(n80610), .A(n106327), .ZN(n80607) );
  NOR4_X1 U65687 ( .A1(n80611), .A2(n80612), .A3(n80613), .A4(n80614), .ZN(
        n80610) );
  OAI21_X1 U65688 ( .B1(n106322), .B2(n104636), .A(n80615), .ZN(n80614) );
  AOI22_X1 U65689 ( .A1(n70346), .A2(n106321), .B1(n70330), .B2(n106320), .ZN(
        n80615) );
  NAND2_X1 U65690 ( .A1(n80616), .A2(n80617), .ZN(n80613) );
  AOI22_X1 U65691 ( .A1(n70366), .A2(n106319), .B1(n70354), .B2(n106318), .ZN(
        n80617) );
  AOI22_X1 U65692 ( .A1(n70358), .A2(n106317), .B1(n70350), .B2(n106316), .ZN(
        n80616) );
  NAND2_X1 U65693 ( .A1(n80618), .A2(n80619), .ZN(n80612) );
  AOI22_X1 U65694 ( .A1(n106315), .A2(n107909), .B1(n70386), .B2(n106314), 
        .ZN(n80619) );
  AOI22_X1 U65695 ( .A1(n106313), .A2(n107900), .B1(n80223), .B2(n107902), 
        .ZN(n80618) );
  NAND2_X1 U65696 ( .A1(n80620), .A2(n80621), .ZN(n80611) );
  AOI22_X1 U65697 ( .A1(n106311), .A2(n107917), .B1(n70394), .B2(n80227), .ZN(
        n80621) );
  AOI22_X1 U65698 ( .A1(n106309), .A2(n107906), .B1(n70382), .B2(n106308), 
        .ZN(n80620) );
  NOR4_X1 U65699 ( .A1(n80622), .A2(n80623), .A3(n80624), .A4(n80625), .ZN(
        n80609) );
  OAI21_X1 U65700 ( .B1(n102178), .B2(n106307), .A(n80626), .ZN(n80625) );
  AOI22_X1 U65701 ( .A1(n70395), .A2(n106306), .B1(n70407), .B2(n106305), .ZN(
        n80626) );
  NAND2_X1 U65702 ( .A1(n80627), .A2(n80628), .ZN(n80624) );
  AOI22_X1 U65703 ( .A1(n106304), .A2(n107859), .B1(n80241), .B2(n107944), 
        .ZN(n80628) );
  AOI22_X1 U65704 ( .A1(n106302), .A2(n107933), .B1(n106301), .B2(n107941), 
        .ZN(n80627) );
  NAND2_X1 U65705 ( .A1(n80629), .A2(n80630), .ZN(n80623) );
  AOI22_X1 U65706 ( .A1(n106300), .A2(n107865), .B1(n70314), .B2(n106299), 
        .ZN(n80630) );
  AOI22_X1 U65707 ( .A1(n80248), .A2(n107869), .B1(n106297), .B2(n107857), 
        .ZN(n80629) );
  NAND2_X1 U65708 ( .A1(n80631), .A2(n80632), .ZN(n80622) );
  AOI22_X1 U65709 ( .A1(n106296), .A2(n107885), .B1(n70342), .B2(n106295), 
        .ZN(n80632) );
  AOI22_X1 U65710 ( .A1(n106294), .A2(n107875), .B1(n70326), .B2(n80255), .ZN(
        n80631) );
  NOR2_X1 U65711 ( .A1(n100561), .A2(n106292), .ZN(n80606) );
  AOI22_X1 U65712 ( .A1(n106291), .A2(n107925), .B1(n106290), .B2(n107937), 
        .ZN(n80604) );
  AOI22_X1 U65713 ( .A1(n70366), .A2(n106746), .B1(n70382), .B2(n105171), .ZN(
        n80603) );
  AOI22_X1 U65714 ( .A1(n70350), .A2(n106286), .B1(n70334), .B2(n106282), .ZN(
        n80602) );
  NAND4_X2 U65715 ( .A1(n80633), .A2(n80634), .A3(n80635), .A4(n80636), .ZN(
        n103970) );
  NOR3_X1 U65716 ( .A1(n80637), .A2(n80638), .A3(n80639), .ZN(n80636) );
  NOR2_X1 U65717 ( .A1(n100594), .A2(n80200), .ZN(n80639) );
  AOI21_X1 U65718 ( .B1(n80640), .B2(n80641), .A(n106323), .ZN(n80638) );
  NOR4_X1 U65719 ( .A1(n80642), .A2(n80643), .A3(n80644), .A4(n80645), .ZN(
        n80641) );
  OAI21_X1 U65720 ( .B1(n106322), .B2(n104635), .A(n80646), .ZN(n80645) );
  AOI22_X1 U65721 ( .A1(n70488), .A2(n106321), .B1(n70472), .B2(n106320), .ZN(
        n80646) );
  NAND2_X1 U65722 ( .A1(n80647), .A2(n80648), .ZN(n80644) );
  AOI22_X1 U65723 ( .A1(n70508), .A2(n106319), .B1(n70496), .B2(n106318), .ZN(
        n80648) );
  AOI22_X1 U65724 ( .A1(n70500), .A2(n106317), .B1(n70492), .B2(n106316), .ZN(
        n80647) );
  NAND2_X1 U65725 ( .A1(n80649), .A2(n80650), .ZN(n80643) );
  AOI22_X1 U65726 ( .A1(n106315), .A2(n108005), .B1(n106314), .B2(n108011), 
        .ZN(n80650) );
  AOI22_X1 U65727 ( .A1(n106313), .A2(n107994), .B1(n80223), .B2(n107998), 
        .ZN(n80649) );
  NAND2_X1 U65728 ( .A1(n80651), .A2(n80652), .ZN(n80642) );
  AOI22_X1 U65729 ( .A1(n106311), .A2(n108014), .B1(n70536), .B2(n80227), .ZN(
        n80652) );
  AOI22_X1 U65730 ( .A1(n106309), .A2(n108002), .B1(n70524), .B2(n106308), 
        .ZN(n80651) );
  NOR4_X1 U65731 ( .A1(n80653), .A2(n80654), .A3(n80655), .A4(n80656), .ZN(
        n80640) );
  OAI21_X1 U65732 ( .B1(n102164), .B2(n106307), .A(n80657), .ZN(n80656) );
  AOI22_X1 U65733 ( .A1(n70537), .A2(n106306), .B1(n70549), .B2(n106305), .ZN(
        n80657) );
  NAND2_X1 U65734 ( .A1(n80658), .A2(n80659), .ZN(n80655) );
  AOI22_X1 U65735 ( .A1(n106304), .A2(n107956), .B1(n80241), .B2(n108040), 
        .ZN(n80659) );
  AOI22_X1 U65736 ( .A1(n106302), .A2(n108029), .B1(n106301), .B2(n108037), 
        .ZN(n80658) );
  NAND2_X1 U65737 ( .A1(n80660), .A2(n80661), .ZN(n80654) );
  AOI22_X1 U65738 ( .A1(n106300), .A2(n107962), .B1(n70456), .B2(n106299), 
        .ZN(n80661) );
  AOI22_X1 U65739 ( .A1(n80248), .A2(n107966), .B1(n106297), .B2(n107954), 
        .ZN(n80660) );
  NAND2_X1 U65740 ( .A1(n80662), .A2(n80663), .ZN(n80653) );
  AOI22_X1 U65741 ( .A1(n106296), .A2(n107980), .B1(n70484), .B2(n106295), 
        .ZN(n80663) );
  AOI22_X1 U65742 ( .A1(n106294), .A2(n107972), .B1(n70468), .B2(n80255), .ZN(
        n80662) );
  NOR2_X1 U65743 ( .A1(n100562), .A2(n80256), .ZN(n80637) );
  AOI22_X1 U65744 ( .A1(n106291), .A2(n108021), .B1(n106290), .B2(n108033), 
        .ZN(n80635) );
  AOI22_X1 U65745 ( .A1(n70508), .A2(n105173), .B1(n70524), .B2(n105171), .ZN(
        n80634) );
  AOI22_X1 U65746 ( .A1(n70492), .A2(n80259), .B1(n70476), .B2(n106282), .ZN(
        n80633) );
  NAND4_X2 U65747 ( .A1(n80664), .A2(n80665), .A3(n80666), .A4(n80667), .ZN(
        n103971) );
  NOR3_X1 U65748 ( .A1(n80668), .A2(n80669), .A3(n80670), .ZN(n80667) );
  NOR2_X1 U65749 ( .A1(n100595), .A2(n106329), .ZN(n80670) );
  AOI21_X1 U65750 ( .B1(n80671), .B2(n80672), .A(n106323), .ZN(n80669) );
  NOR4_X1 U65751 ( .A1(n80673), .A2(n80674), .A3(n80675), .A4(n80676), .ZN(
        n80672) );
  OAI21_X1 U65752 ( .B1(n106322), .B2(n104634), .A(n80677), .ZN(n80676) );
  AOI22_X1 U65753 ( .A1(n69541), .A2(n106321), .B1(n106320), .B2(n107241), 
        .ZN(n80677) );
  NAND2_X1 U65754 ( .A1(n80678), .A2(n80679), .ZN(n80675) );
  AOI22_X1 U65755 ( .A1(n69561), .A2(n106319), .B1(n69549), .B2(n106318), .ZN(
        n80679) );
  AOI22_X1 U65756 ( .A1(n69553), .A2(n106317), .B1(n69545), .B2(n106316), .ZN(
        n80678) );
  NAND2_X1 U65757 ( .A1(n80680), .A2(n80681), .ZN(n80674) );
  AOI22_X1 U65758 ( .A1(n106315), .A2(n107276), .B1(n69581), .B2(n106314), 
        .ZN(n80681) );
  AOI22_X1 U65759 ( .A1(n106313), .A2(n107264), .B1(n106312), .B2(n107269), 
        .ZN(n80680) );
  NAND2_X1 U65760 ( .A1(n80682), .A2(n80683), .ZN(n80673) );
  AOI22_X1 U65761 ( .A1(n106311), .A2(n107284), .B1(n69589), .B2(n80227), .ZN(
        n80683) );
  AOI22_X1 U65762 ( .A1(n106309), .A2(n107273), .B1(n69577), .B2(n106308), 
        .ZN(n80682) );
  NOR4_X1 U65763 ( .A1(n80684), .A2(n80685), .A3(n80686), .A4(n80687), .ZN(
        n80671) );
  OAI21_X1 U65764 ( .B1(n102149), .B2(n106307), .A(n80688), .ZN(n80687) );
  AOI22_X1 U65765 ( .A1(n69483), .A2(n106306), .B1(n69459), .B2(n106305), .ZN(
        n80688) );
  NAND2_X1 U65766 ( .A1(n80689), .A2(n80690), .ZN(n80686) );
  AOI22_X1 U65767 ( .A1(n106304), .A2(n107218), .B1(n80241), .B2(n107168), 
        .ZN(n80690) );
  AOI22_X1 U65768 ( .A1(n106302), .A2(n107190), .B1(n106301), .B2(n107174), 
        .ZN(n80689) );
  NAND2_X1 U65769 ( .A1(n80691), .A2(n80692), .ZN(n80685) );
  AOI22_X1 U65770 ( .A1(n106300), .A2(n107225), .B1(n69509), .B2(n106299), 
        .ZN(n80692) );
  AOI22_X1 U65771 ( .A1(n80248), .A2(n107229), .B1(n106297), .B2(n107216), 
        .ZN(n80691) );
  NAND2_X1 U65772 ( .A1(n80693), .A2(n80694), .ZN(n80684) );
  AOI22_X1 U65773 ( .A1(n106296), .A2(n107247), .B1(n106295), .B2(n107251), 
        .ZN(n80694) );
  AOI22_X1 U65774 ( .A1(n106294), .A2(n107236), .B1(n69521), .B2(n80255), .ZN(
        n80693) );
  NOR2_X1 U65775 ( .A1(n100563), .A2(n106292), .ZN(n80668) );
  AOI22_X1 U65776 ( .A1(n106291), .A2(n107206), .B1(n106290), .B2(n107182), 
        .ZN(n80666) );
  AOI22_X1 U65777 ( .A1(n69561), .A2(n106746), .B1(n69577), .B2(n105171), .ZN(
        n80665) );
  AOI22_X1 U65778 ( .A1(n69545), .A2(n80259), .B1(n69529), .B2(n106284), .ZN(
        n80664) );
  NAND4_X2 U65779 ( .A1(n80695), .A2(n80696), .A3(n80697), .A4(n80698), .ZN(
        n103972) );
  NOR3_X1 U65780 ( .A1(n80699), .A2(n80700), .A3(n80701), .ZN(n80698) );
  NOR2_X1 U65781 ( .A1(n100596), .A2(n80200), .ZN(n80701) );
  AOI21_X1 U65782 ( .B1(n80702), .B2(n80703), .A(n106324), .ZN(n80700) );
  NOR4_X1 U65783 ( .A1(n80704), .A2(n80705), .A3(n80706), .A4(n80707), .ZN(
        n80703) );
  OAI21_X1 U65784 ( .B1(n106322), .B2(n104633), .A(n80708), .ZN(n80707) );
  AOI22_X1 U65785 ( .A1(n70202), .A2(n106321), .B1(n106320), .B2(n107780), 
        .ZN(n80708) );
  NAND2_X1 U65786 ( .A1(n80709), .A2(n80710), .ZN(n80706) );
  AOI22_X1 U65787 ( .A1(n70222), .A2(n106319), .B1(n70210), .B2(n106318), .ZN(
        n80710) );
  AOI22_X1 U65788 ( .A1(n70214), .A2(n106317), .B1(n70206), .B2(n106316), .ZN(
        n80709) );
  NAND2_X1 U65789 ( .A1(n80711), .A2(n80712), .ZN(n80705) );
  AOI22_X1 U65790 ( .A1(n106315), .A2(n107814), .B1(n70242), .B2(n106314), 
        .ZN(n80712) );
  AOI22_X1 U65791 ( .A1(n106313), .A2(n107801), .B1(n106312), .B2(n107806), 
        .ZN(n80711) );
  NAND2_X1 U65792 ( .A1(n80713), .A2(n80714), .ZN(n80704) );
  AOI22_X1 U65793 ( .A1(n106311), .A2(n107822), .B1(n70250), .B2(n106310), 
        .ZN(n80714) );
  AOI22_X1 U65794 ( .A1(n106309), .A2(n107810), .B1(n70238), .B2(n106308), 
        .ZN(n80713) );
  NOR4_X1 U65795 ( .A1(n80715), .A2(n80716), .A3(n80717), .A4(n80718), .ZN(
        n80702) );
  OAI21_X1 U65796 ( .B1(n102133), .B2(n106307), .A(n80719), .ZN(n80718) );
  AOI22_X1 U65797 ( .A1(n70251), .A2(n106306), .B1(n70263), .B2(n106305), .ZN(
        n80719) );
  NAND2_X1 U65798 ( .A1(n80720), .A2(n80721), .ZN(n80717) );
  AOI22_X1 U65799 ( .A1(n106304), .A2(n107756), .B1(n106303), .B2(n107849), 
        .ZN(n80721) );
  AOI22_X1 U65800 ( .A1(n106302), .A2(n107838), .B1(n106301), .B2(n107846), 
        .ZN(n80720) );
  NAND2_X1 U65801 ( .A1(n80722), .A2(n80723), .ZN(n80716) );
  AOI22_X1 U65802 ( .A1(n106300), .A2(n107763), .B1(n70170), .B2(n106299), 
        .ZN(n80723) );
  AOI22_X1 U65803 ( .A1(n106298), .A2(n107767), .B1(n80249), .B2(n107754), 
        .ZN(n80722) );
  NAND2_X1 U65804 ( .A1(n80724), .A2(n80725), .ZN(n80715) );
  AOI22_X1 U65805 ( .A1(n106296), .A2(n107786), .B1(n106295), .B2(n107790), 
        .ZN(n80725) );
  AOI22_X1 U65806 ( .A1(n106294), .A2(n107775), .B1(n70182), .B2(n106293), 
        .ZN(n80724) );
  NOR2_X1 U65807 ( .A1(n100564), .A2(n80256), .ZN(n80699) );
  AOI22_X1 U65808 ( .A1(n106291), .A2(n107829), .B1(n106290), .B2(n107842), 
        .ZN(n80697) );
  AOI22_X1 U65809 ( .A1(n70222), .A2(n105175), .B1(n70238), .B2(n105171), .ZN(
        n80696) );
  AOI22_X1 U65810 ( .A1(n70206), .A2(n106286), .B1(n70190), .B2(n106283), .ZN(
        n80695) );
  NAND4_X2 U65811 ( .A1(n80726), .A2(n80727), .A3(n80728), .A4(n80729), .ZN(
        n103973) );
  NOR3_X1 U65812 ( .A1(n80730), .A2(n80731), .A3(n80732), .ZN(n80729) );
  NOR2_X1 U65813 ( .A1(n100597), .A2(n106329), .ZN(n80732) );
  AOI21_X1 U65814 ( .B1(n80733), .B2(n80734), .A(n106325), .ZN(n80731) );
  NOR4_X1 U65815 ( .A1(n80735), .A2(n80736), .A3(n80737), .A4(n80738), .ZN(
        n80734) );
  OAI21_X1 U65816 ( .B1(n106322), .B2(n104632), .A(n80739), .ZN(n80738) );
  AOI22_X1 U65817 ( .A1(n74048), .A2(n106321), .B1(n74032), .B2(n106320), .ZN(
        n80739) );
  NAND2_X1 U65818 ( .A1(n80740), .A2(n80741), .ZN(n80737) );
  AOI22_X1 U65819 ( .A1(n74068), .A2(n106319), .B1(n74056), .B2(n106318), .ZN(
        n80741) );
  AOI22_X1 U65820 ( .A1(n74060), .A2(n106317), .B1(n74052), .B2(n106316), .ZN(
        n80740) );
  NAND2_X1 U65821 ( .A1(n80742), .A2(n80743), .ZN(n80736) );
  AOI22_X1 U65822 ( .A1(n106315), .A2(n110710), .B1(n74088), .B2(n106314), 
        .ZN(n80743) );
  AOI22_X1 U65823 ( .A1(n106313), .A2(n110700), .B1(n106312), .B2(n110703), 
        .ZN(n80742) );
  NAND2_X1 U65824 ( .A1(n80744), .A2(n80745), .ZN(n80735) );
  AOI22_X1 U65825 ( .A1(n106311), .A2(n110718), .B1(n74096), .B2(n80227), .ZN(
        n80745) );
  AOI22_X1 U65826 ( .A1(n106309), .A2(n110707), .B1(n74084), .B2(n106308), 
        .ZN(n80744) );
  NOR4_X1 U65827 ( .A1(n80746), .A2(n80747), .A3(n80748), .A4(n80749), .ZN(
        n80733) );
  OAI21_X1 U65828 ( .B1(n102119), .B2(n106307), .A(n80750), .ZN(n80749) );
  AOI22_X1 U65829 ( .A1(n74097), .A2(n106306), .B1(n74109), .B2(n106305), .ZN(
        n80750) );
  NAND2_X1 U65830 ( .A1(n80751), .A2(n80752), .ZN(n80748) );
  AOI22_X1 U65831 ( .A1(n106304), .A2(n110659), .B1(n80241), .B2(n110744), 
        .ZN(n80752) );
  AOI22_X1 U65832 ( .A1(n106302), .A2(n110733), .B1(n106301), .B2(n110741), 
        .ZN(n80751) );
  NAND2_X1 U65833 ( .A1(n80753), .A2(n80754), .ZN(n80747) );
  AOI22_X1 U65834 ( .A1(n106300), .A2(n110666), .B1(n74016), .B2(n106299), 
        .ZN(n80754) );
  AOI22_X1 U65835 ( .A1(n80248), .A2(n110670), .B1(n106297), .B2(n110657), 
        .ZN(n80753) );
  NAND2_X1 U65836 ( .A1(n80755), .A2(n80756), .ZN(n80746) );
  AOI22_X1 U65837 ( .A1(n106296), .A2(n110687), .B1(n74044), .B2(n106295), 
        .ZN(n80756) );
  AOI22_X1 U65838 ( .A1(n106294), .A2(n110677), .B1(n74028), .B2(n80255), .ZN(
        n80755) );
  NOR2_X1 U65839 ( .A1(n100565), .A2(n106292), .ZN(n80730) );
  AOI22_X1 U65840 ( .A1(n106291), .A2(n110725), .B1(n106290), .B2(n110737), 
        .ZN(n80728) );
  AOI22_X1 U65841 ( .A1(n74068), .A2(n105175), .B1(n74084), .B2(n105171), .ZN(
        n80727) );
  AOI22_X1 U65842 ( .A1(n74052), .A2(n80259), .B1(n74036), .B2(n106285), .ZN(
        n80726) );
  NAND4_X2 U65843 ( .A1(n80757), .A2(n80758), .A3(n80759), .A4(n80760), .ZN(
        n103974) );
  NOR3_X1 U65844 ( .A1(n80761), .A2(n80762), .A3(n80763), .ZN(n80760) );
  NOR2_X1 U65845 ( .A1(n100598), .A2(n80200), .ZN(n80763) );
  AOI21_X1 U65846 ( .B1(n80764), .B2(n80765), .A(n106326), .ZN(n80762) );
  NOR4_X1 U65847 ( .A1(n80766), .A2(n80767), .A3(n80768), .A4(n80769), .ZN(
        n80765) );
  OAI21_X1 U65848 ( .B1(n106322), .B2(n104631), .A(n80770), .ZN(n80769) );
  AOI22_X1 U65849 ( .A1(n70635), .A2(n106321), .B1(n70619), .B2(n106320), .ZN(
        n80770) );
  NAND2_X1 U65850 ( .A1(n80771), .A2(n80772), .ZN(n80768) );
  AOI22_X1 U65851 ( .A1(n70655), .A2(n106319), .B1(n70643), .B2(n106318), .ZN(
        n80772) );
  AOI22_X1 U65852 ( .A1(n70647), .A2(n106317), .B1(n70639), .B2(n106316), .ZN(
        n80771) );
  NAND2_X1 U65853 ( .A1(n80773), .A2(n80774), .ZN(n80767) );
  AOI22_X1 U65854 ( .A1(n106315), .A2(n108113), .B1(n70675), .B2(n106314), 
        .ZN(n80774) );
  AOI22_X1 U65855 ( .A1(n106313), .A2(n108103), .B1(n106312), .B2(n108106), 
        .ZN(n80773) );
  NAND2_X1 U65856 ( .A1(n80775), .A2(n80776), .ZN(n80766) );
  AOI22_X1 U65857 ( .A1(n106311), .A2(n108121), .B1(n70683), .B2(n106310), 
        .ZN(n80776) );
  AOI22_X1 U65858 ( .A1(n106309), .A2(n108110), .B1(n70671), .B2(n106308), 
        .ZN(n80775) );
  NOR4_X1 U65859 ( .A1(n80777), .A2(n80778), .A3(n80779), .A4(n80780), .ZN(
        n80764) );
  OAI21_X1 U65860 ( .B1(n102105), .B2(n106307), .A(n80781), .ZN(n80780) );
  AOI22_X1 U65861 ( .A1(n70684), .A2(n106306), .B1(n70696), .B2(n106305), .ZN(
        n80781) );
  NAND2_X1 U65862 ( .A1(n80782), .A2(n80783), .ZN(n80779) );
  AOI22_X1 U65863 ( .A1(n106304), .A2(n108058), .B1(n106303), .B2(n108149), 
        .ZN(n80783) );
  AOI22_X1 U65864 ( .A1(n106302), .A2(n108138), .B1(n106301), .B2(n108146), 
        .ZN(n80782) );
  NAND2_X1 U65865 ( .A1(n80784), .A2(n80785), .ZN(n80778) );
  AOI22_X1 U65866 ( .A1(n106300), .A2(n108065), .B1(n70603), .B2(n106299), 
        .ZN(n80785) );
  AOI22_X1 U65867 ( .A1(n106298), .A2(n108069), .B1(n80249), .B2(n108056), 
        .ZN(n80784) );
  NAND2_X1 U65868 ( .A1(n80786), .A2(n80787), .ZN(n80777) );
  AOI22_X1 U65869 ( .A1(n106296), .A2(n108087), .B1(n70631), .B2(n106295), 
        .ZN(n80787) );
  AOI22_X1 U65870 ( .A1(n106294), .A2(n108077), .B1(n70615), .B2(n106293), 
        .ZN(n80786) );
  NOR2_X1 U65871 ( .A1(n100566), .A2(n80256), .ZN(n80761) );
  AOI22_X1 U65872 ( .A1(n106291), .A2(n108129), .B1(n106290), .B2(n108142), 
        .ZN(n80759) );
  AOI22_X1 U65873 ( .A1(n70655), .A2(n105174), .B1(n70671), .B2(n105171), .ZN(
        n80758) );
  AOI22_X1 U65874 ( .A1(n70639), .A2(n106286), .B1(n70623), .B2(n106284), .ZN(
        n80757) );
  NAND4_X2 U65875 ( .A1(n80788), .A2(n80789), .A3(n80790), .A4(n80791), .ZN(
        n103975) );
  NOR3_X1 U65876 ( .A1(n80792), .A2(n80793), .A3(n80794), .ZN(n80791) );
  NOR2_X1 U65877 ( .A1(n100599), .A2(n106329), .ZN(n80794) );
  AOI21_X1 U65878 ( .B1(n80795), .B2(n80796), .A(n106324), .ZN(n80793) );
  NOR4_X1 U65879 ( .A1(n80797), .A2(n80798), .A3(n80799), .A4(n80800), .ZN(
        n80796) );
  OAI21_X1 U65880 ( .B1(n106322), .B2(n104630), .A(n80801), .ZN(n80800) );
  AOI22_X1 U65881 ( .A1(n74189), .A2(n106321), .B1(n106320), .B2(n110779), 
        .ZN(n80801) );
  NAND2_X1 U65882 ( .A1(n80802), .A2(n80803), .ZN(n80799) );
  AOI22_X1 U65883 ( .A1(n74209), .A2(n106319), .B1(n74197), .B2(n106318), .ZN(
        n80803) );
  AOI22_X1 U65884 ( .A1(n74201), .A2(n106317), .B1(n106316), .B2(n110794), 
        .ZN(n80802) );
  NAND2_X1 U65885 ( .A1(n80804), .A2(n80805), .ZN(n80798) );
  AOI22_X1 U65886 ( .A1(n106315), .A2(n110812), .B1(n74229), .B2(n106314), 
        .ZN(n80805) );
  AOI22_X1 U65887 ( .A1(n106313), .A2(n110802), .B1(n106312), .B2(n110805), 
        .ZN(n80804) );
  NAND2_X1 U65888 ( .A1(n80806), .A2(n80807), .ZN(n80797) );
  AOI22_X1 U65889 ( .A1(n106311), .A2(n110820), .B1(n74237), .B2(n80227), .ZN(
        n80807) );
  AOI22_X1 U65890 ( .A1(n106309), .A2(n110809), .B1(n74225), .B2(n106308), 
        .ZN(n80806) );
  NOR4_X1 U65891 ( .A1(n80808), .A2(n80809), .A3(n80810), .A4(n80811), .ZN(
        n80795) );
  OAI21_X1 U65892 ( .B1(n102091), .B2(n106307), .A(n80812), .ZN(n80811) );
  AOI22_X1 U65893 ( .A1(n74238), .A2(n106306), .B1(n74250), .B2(n106305), .ZN(
        n80812) );
  NAND2_X1 U65894 ( .A1(n80813), .A2(n80814), .ZN(n80810) );
  AOI22_X1 U65895 ( .A1(n106304), .A2(n110756), .B1(n80241), .B2(n110847), 
        .ZN(n80814) );
  AOI22_X1 U65896 ( .A1(n106302), .A2(n110836), .B1(n106301), .B2(n110844), 
        .ZN(n80813) );
  NAND2_X1 U65897 ( .A1(n80815), .A2(n80816), .ZN(n80809) );
  AOI22_X1 U65898 ( .A1(n106300), .A2(n110763), .B1(n74157), .B2(n106299), 
        .ZN(n80816) );
  AOI22_X1 U65899 ( .A1(n80248), .A2(n110767), .B1(n106297), .B2(n110754), 
        .ZN(n80815) );
  NAND2_X1 U65900 ( .A1(n80817), .A2(n80818), .ZN(n80808) );
  AOI22_X1 U65901 ( .A1(n80252), .A2(n110785), .B1(n106295), .B2(n110789), 
        .ZN(n80818) );
  AOI22_X1 U65902 ( .A1(n106294), .A2(n110774), .B1(n74169), .B2(n80255), .ZN(
        n80817) );
  NOR2_X1 U65903 ( .A1(n100567), .A2(n106292), .ZN(n80792) );
  AOI22_X1 U65904 ( .A1(n106291), .A2(n110828), .B1(n106290), .B2(n110840), 
        .ZN(n80790) );
  AOI22_X1 U65905 ( .A1(n74209), .A2(n105173), .B1(n74225), .B2(n105171), .ZN(
        n80789) );
  AOI22_X1 U65906 ( .A1(n106286), .A2(n110794), .B1(n74177), .B2(n106282), 
        .ZN(n80788) );
  NAND4_X2 U65907 ( .A1(n80819), .A2(n80820), .A3(n80821), .A4(n80822), .ZN(
        n103976) );
  NOR3_X1 U65908 ( .A1(n80823), .A2(n80824), .A3(n80825), .ZN(n80822) );
  NOR2_X1 U65909 ( .A1(n100600), .A2(n80200), .ZN(n80825) );
  AOI21_X1 U65910 ( .B1(n80826), .B2(n80827), .A(n106325), .ZN(n80824) );
  NOR4_X1 U65911 ( .A1(n80828), .A2(n80829), .A3(n80830), .A4(n80831), .ZN(
        n80827) );
  OAI21_X1 U65912 ( .B1(n106322), .B2(n104629), .A(n80832), .ZN(n80831) );
  AOI22_X1 U65913 ( .A1(n74329), .A2(n106321), .B1(n80211), .B2(n110880), .ZN(
        n80832) );
  NAND2_X1 U65914 ( .A1(n80833), .A2(n80834), .ZN(n80830) );
  AOI22_X1 U65915 ( .A1(n74349), .A2(n106319), .B1(n74337), .B2(n106318), .ZN(
        n80834) );
  AOI22_X1 U65916 ( .A1(n74341), .A2(n106317), .B1(n80217), .B2(n110893), .ZN(
        n80833) );
  NAND2_X1 U65917 ( .A1(n80835), .A2(n80836), .ZN(n80829) );
  AOI22_X1 U65918 ( .A1(n106315), .A2(n110912), .B1(n106314), .B2(n110918), 
        .ZN(n80836) );
  AOI22_X1 U65919 ( .A1(n106313), .A2(n110899), .B1(n106312), .B2(n110904), 
        .ZN(n80835) );
  NAND2_X1 U65920 ( .A1(n80837), .A2(n80838), .ZN(n80828) );
  AOI22_X1 U65921 ( .A1(n106311), .A2(n110921), .B1(n74377), .B2(n106310), 
        .ZN(n80838) );
  AOI22_X1 U65922 ( .A1(n106309), .A2(n110908), .B1(n74365), .B2(n106308), 
        .ZN(n80837) );
  NOR4_X1 U65923 ( .A1(n80839), .A2(n80840), .A3(n80841), .A4(n80842), .ZN(
        n80826) );
  OAI21_X1 U65924 ( .B1(n102074), .B2(n106307), .A(n80843), .ZN(n80842) );
  AOI22_X1 U65925 ( .A1(n74378), .A2(n106306), .B1(n74390), .B2(n106305), .ZN(
        n80843) );
  NAND2_X1 U65926 ( .A1(n80844), .A2(n80845), .ZN(n80841) );
  AOI22_X1 U65927 ( .A1(n106304), .A2(n110857), .B1(n106303), .B2(n110948), 
        .ZN(n80845) );
  AOI22_X1 U65928 ( .A1(n106302), .A2(n110937), .B1(n106301), .B2(n110945), 
        .ZN(n80844) );
  NAND2_X1 U65929 ( .A1(n80846), .A2(n80847), .ZN(n80840) );
  AOI22_X1 U65930 ( .A1(n106300), .A2(n110864), .B1(n74297), .B2(n106299), 
        .ZN(n80847) );
  AOI22_X1 U65931 ( .A1(n106298), .A2(n110868), .B1(n80249), .B2(n110855), 
        .ZN(n80846) );
  NAND2_X1 U65932 ( .A1(n80848), .A2(n80849), .ZN(n80839) );
  AOI22_X1 U65933 ( .A1(n80252), .A2(n110885), .B1(n80253), .B2(n110889), .ZN(
        n80849) );
  AOI22_X1 U65934 ( .A1(n106294), .A2(n110875), .B1(n74309), .B2(n106293), 
        .ZN(n80848) );
  NOR2_X1 U65935 ( .A1(n100568), .A2(n80256), .ZN(n80823) );
  AOI22_X1 U65936 ( .A1(n106291), .A2(n110929), .B1(n106290), .B2(n110941), 
        .ZN(n80821) );
  AOI22_X1 U65937 ( .A1(n74349), .A2(n105175), .B1(n74365), .B2(n105171), .ZN(
        n80820) );
  AOI22_X1 U65938 ( .A1(n80259), .A2(n110893), .B1(n74317), .B2(n106285), .ZN(
        n80819) );
  NAND4_X2 U65939 ( .A1(n80850), .A2(n80851), .A3(n80852), .A4(n80853), .ZN(
        n103977) );
  NOR3_X1 U65940 ( .A1(n80854), .A2(n80855), .A3(n80856), .ZN(n80853) );
  NOR2_X1 U65941 ( .A1(n100601), .A2(n106329), .ZN(n80856) );
  AOI21_X1 U65942 ( .B1(n80857), .B2(n80858), .A(n106326), .ZN(n80855) );
  NOR4_X1 U65943 ( .A1(n80859), .A2(n80860), .A3(n80861), .A4(n80862), .ZN(
        n80858) );
  OAI21_X1 U65944 ( .B1(n80208), .B2(n104628), .A(n80863), .ZN(n80862) );
  AOI22_X1 U65945 ( .A1(n73765), .A2(n106321), .B1(n80211), .B2(n110474), .ZN(
        n80863) );
  NAND2_X1 U65946 ( .A1(n80864), .A2(n80865), .ZN(n80861) );
  AOI22_X1 U65947 ( .A1(n73785), .A2(n106319), .B1(n73773), .B2(n80215), .ZN(
        n80865) );
  AOI22_X1 U65948 ( .A1(n73777), .A2(n106317), .B1(n80217), .B2(n110487), .ZN(
        n80864) );
  NAND2_X1 U65949 ( .A1(n80866), .A2(n80867), .ZN(n80860) );
  AOI22_X1 U65950 ( .A1(n106315), .A2(n110507), .B1(n73805), .B2(n106314), 
        .ZN(n80867) );
  AOI22_X1 U65951 ( .A1(n80222), .A2(n110494), .B1(n106312), .B2(n110499), 
        .ZN(n80866) );
  NAND2_X1 U65952 ( .A1(n80868), .A2(n80869), .ZN(n80859) );
  AOI22_X1 U65953 ( .A1(n106311), .A2(n110515), .B1(n73813), .B2(n80227), .ZN(
        n80869) );
  AOI22_X1 U65954 ( .A1(n106309), .A2(n110503), .B1(n73801), .B2(n80229), .ZN(
        n80868) );
  NOR4_X1 U65955 ( .A1(n80870), .A2(n80871), .A3(n80872), .A4(n80873), .ZN(
        n80857) );
  OAI21_X1 U65956 ( .B1(n102056), .B2(n80234), .A(n80874), .ZN(n80873) );
  AOI22_X1 U65957 ( .A1(n73814), .A2(n106306), .B1(n73826), .B2(n106305), .ZN(
        n80874) );
  NAND2_X1 U65958 ( .A1(n80875), .A2(n80876), .ZN(n80872) );
  AOI22_X1 U65959 ( .A1(n106304), .A2(n110452), .B1(n80241), .B2(n110541), 
        .ZN(n80876) );
  AOI22_X1 U65960 ( .A1(n80242), .A2(n110530), .B1(n106301), .B2(n110538), 
        .ZN(n80875) );
  NAND2_X1 U65961 ( .A1(n80877), .A2(n80878), .ZN(n80871) );
  AOI22_X1 U65962 ( .A1(n106300), .A2(n110459), .B1(n73733), .B2(n106299), 
        .ZN(n80878) );
  AOI22_X1 U65963 ( .A1(n80248), .A2(n110463), .B1(n106297), .B2(n110450), 
        .ZN(n80877) );
  NAND2_X1 U65964 ( .A1(n80879), .A2(n80880), .ZN(n80870) );
  AOI22_X1 U65965 ( .A1(n73757), .A2(n106296), .B1(n80253), .B2(n110483), .ZN(
        n80880) );
  AOI22_X1 U65966 ( .A1(n106294), .A2(n110470), .B1(n73745), .B2(n80255), .ZN(
        n80879) );
  NOR2_X1 U65967 ( .A1(n100569), .A2(n106292), .ZN(n80854) );
  AOI22_X1 U65968 ( .A1(n106291), .A2(n110522), .B1(n106290), .B2(n110534), 
        .ZN(n80852) );
  AOI22_X1 U65969 ( .A1(n73785), .A2(n106746), .B1(n73801), .B2(n105171), .ZN(
        n80851) );
  AOI22_X1 U65970 ( .A1(n106287), .A2(n110487), .B1(n73753), .B2(n106282), 
        .ZN(n80850) );
  NAND4_X2 U65971 ( .A1(n80881), .A2(n80882), .A3(n80883), .A4(n80884), .ZN(
        n103978) );
  NOR3_X1 U65972 ( .A1(n80885), .A2(n80886), .A3(n80887), .ZN(n80884) );
  NOR2_X1 U65973 ( .A1(n100602), .A2(n80200), .ZN(n80887) );
  AOI21_X1 U65974 ( .B1(n80888), .B2(n80889), .A(n106326), .ZN(n80886) );
  NOR4_X1 U65975 ( .A1(n80890), .A2(n80891), .A3(n80892), .A4(n80893), .ZN(
        n80889) );
  OAI21_X1 U65976 ( .B1(n80208), .B2(n104627), .A(n80894), .ZN(n80893) );
  AOI22_X1 U65977 ( .A1(n73469), .A2(n106321), .B1(n80211), .B2(n110256), .ZN(
        n80894) );
  NAND2_X1 U65978 ( .A1(n80895), .A2(n80896), .ZN(n80892) );
  AOI22_X1 U65979 ( .A1(n73489), .A2(n106319), .B1(n73477), .B2(n80215), .ZN(
        n80896) );
  AOI22_X1 U65980 ( .A1(n73481), .A2(n106317), .B1(n80217), .B2(n110270), .ZN(
        n80895) );
  NAND2_X1 U65981 ( .A1(n80897), .A2(n80898), .ZN(n80891) );
  AOI22_X1 U65982 ( .A1(n106315), .A2(n110290), .B1(n80221), .B2(n110296), 
        .ZN(n80898) );
  AOI22_X1 U65983 ( .A1(n80222), .A2(n110277), .B1(n106312), .B2(n110282), 
        .ZN(n80897) );
  NAND2_X1 U65984 ( .A1(n80899), .A2(n80900), .ZN(n80890) );
  AOI22_X1 U65985 ( .A1(n106311), .A2(n110299), .B1(n73517), .B2(n80227), .ZN(
        n80900) );
  AOI22_X1 U65986 ( .A1(n106309), .A2(n110286), .B1(n73505), .B2(n80229), .ZN(
        n80899) );
  NOR4_X1 U65987 ( .A1(n80901), .A2(n80902), .A3(n80903), .A4(n80904), .ZN(
        n80888) );
  OAI21_X1 U65988 ( .B1(n102040), .B2(n80234), .A(n80905), .ZN(n80904) );
  AOI22_X1 U65989 ( .A1(n73518), .A2(n106306), .B1(n73530), .B2(n106305), .ZN(
        n80905) );
  NAND2_X1 U65990 ( .A1(n80906), .A2(n80907), .ZN(n80903) );
  AOI22_X1 U65991 ( .A1(n106304), .A2(n110234), .B1(n80241), .B2(n110326), 
        .ZN(n80907) );
  AOI22_X1 U65992 ( .A1(n80242), .A2(n110315), .B1(n106301), .B2(n110323), 
        .ZN(n80906) );
  NAND2_X1 U65993 ( .A1(n80908), .A2(n80909), .ZN(n80902) );
  AOI22_X1 U65994 ( .A1(n106300), .A2(n110241), .B1(n73437), .B2(n106299), 
        .ZN(n80909) );
  AOI22_X1 U65995 ( .A1(n80248), .A2(n110245), .B1(n106297), .B2(n110232), 
        .ZN(n80908) );
  NAND2_X1 U65996 ( .A1(n80910), .A2(n80911), .ZN(n80901) );
  AOI22_X1 U65997 ( .A1(n73461), .A2(n106296), .B1(n80253), .B2(n110265), .ZN(
        n80911) );
  AOI22_X1 U65998 ( .A1(n106294), .A2(n110252), .B1(n73449), .B2(n80255), .ZN(
        n80910) );
  NOR2_X1 U65999 ( .A1(n100570), .A2(n80256), .ZN(n80885) );
  AOI22_X1 U66000 ( .A1(n106291), .A2(n110307), .B1(n106290), .B2(n110319), 
        .ZN(n80883) );
  AOI22_X1 U66001 ( .A1(n73489), .A2(n106746), .B1(n73505), .B2(n105171), .ZN(
        n80882) );
  AOI22_X1 U66002 ( .A1(n106286), .A2(n110270), .B1(n73457), .B2(n106285), 
        .ZN(n80881) );
  NAND4_X2 U66003 ( .A1(n80912), .A2(n80913), .A3(n80914), .A4(n80915), .ZN(
        n103979) );
  NOR3_X1 U66004 ( .A1(n80916), .A2(n80917), .A3(n80918), .ZN(n80915) );
  NOR2_X1 U66005 ( .A1(n100603), .A2(n106329), .ZN(n80918) );
  AOI21_X1 U66006 ( .B1(n80919), .B2(n80920), .A(n106325), .ZN(n80917) );
  NOR4_X1 U66007 ( .A1(n80921), .A2(n80922), .A3(n80923), .A4(n80924), .ZN(
        n80920) );
  OAI21_X1 U66008 ( .B1(n80208), .B2(n104626), .A(n80925), .ZN(n80924) );
  AOI22_X1 U66009 ( .A1(n73906), .A2(n106321), .B1(n80211), .B2(n110573), .ZN(
        n80925) );
  NAND2_X1 U66010 ( .A1(n80926), .A2(n80927), .ZN(n80923) );
  AOI22_X1 U66011 ( .A1(n73926), .A2(n106319), .B1(n73914), .B2(n80215), .ZN(
        n80927) );
  AOI22_X1 U66012 ( .A1(n73918), .A2(n106317), .B1(n80217), .B2(n110588), .ZN(
        n80926) );
  NAND2_X1 U66013 ( .A1(n80928), .A2(n80929), .ZN(n80922) );
  AOI22_X1 U66014 ( .A1(n106315), .A2(n110610), .B1(n80221), .B2(n110616), 
        .ZN(n80929) );
  AOI22_X1 U66015 ( .A1(n80222), .A2(n110596), .B1(n106312), .B2(n110602), 
        .ZN(n80928) );
  NAND2_X1 U66016 ( .A1(n80930), .A2(n80931), .ZN(n80921) );
  AOI22_X1 U66017 ( .A1(n106311), .A2(n110620), .B1(n73954), .B2(n106310), 
        .ZN(n80931) );
  AOI22_X1 U66018 ( .A1(n106309), .A2(n110606), .B1(n73942), .B2(n80229), .ZN(
        n80930) );
  NOR4_X1 U66019 ( .A1(n80932), .A2(n80933), .A3(n80934), .A4(n80935), .ZN(
        n80919) );
  OAI21_X1 U66020 ( .B1(n102023), .B2(n80234), .A(n80936), .ZN(n80935) );
  AOI22_X1 U66021 ( .A1(n73955), .A2(n106306), .B1(n73967), .B2(n106305), .ZN(
        n80936) );
  NAND2_X1 U66022 ( .A1(n80937), .A2(n80938), .ZN(n80934) );
  AOI22_X1 U66023 ( .A1(n106304), .A2(n110551), .B1(n106303), .B2(n110646), 
        .ZN(n80938) );
  AOI22_X1 U66024 ( .A1(n80242), .A2(n110635), .B1(n106301), .B2(n110643), 
        .ZN(n80937) );
  NAND2_X1 U66025 ( .A1(n80939), .A2(n80940), .ZN(n80933) );
  AOI22_X1 U66026 ( .A1(n106300), .A2(n110558), .B1(n73874), .B2(n106299), 
        .ZN(n80940) );
  AOI22_X1 U66027 ( .A1(n106298), .A2(n110562), .B1(n106297), .B2(n110549), 
        .ZN(n80939) );
  NAND2_X1 U66028 ( .A1(n80941), .A2(n80942), .ZN(n80932) );
  AOI22_X1 U66029 ( .A1(n80252), .A2(n110579), .B1(n80253), .B2(n110583), .ZN(
        n80942) );
  AOI22_X1 U66030 ( .A1(n106294), .A2(n110569), .B1(n73886), .B2(n106293), 
        .ZN(n80941) );
  NOR2_X1 U66031 ( .A1(n100571), .A2(n106292), .ZN(n80916) );
  AOI22_X1 U66032 ( .A1(n106291), .A2(n110627), .B1(n106290), .B2(n110639), 
        .ZN(n80914) );
  AOI22_X1 U66033 ( .A1(n73926), .A2(n105175), .B1(n73942), .B2(n105171), .ZN(
        n80913) );
  AOI22_X1 U66034 ( .A1(n106288), .A2(n110588), .B1(n73894), .B2(n106285), 
        .ZN(n80912) );
  NAND4_X2 U66035 ( .A1(n80943), .A2(n80944), .A3(n80945), .A4(n80946), .ZN(
        n103980) );
  NOR3_X1 U66036 ( .A1(n80947), .A2(n80948), .A3(n80949), .ZN(n80946) );
  NOR2_X1 U66037 ( .A1(n100604), .A2(n106329), .ZN(n80949) );
  AOI21_X1 U66038 ( .B1(n80950), .B2(n80951), .A(n106323), .ZN(n80948) );
  NOR4_X1 U66039 ( .A1(n80952), .A2(n80953), .A3(n80954), .A4(n80955), .ZN(
        n80951) );
  OAI21_X1 U66040 ( .B1(n80208), .B2(n104625), .A(n80956), .ZN(n80955) );
  AOI22_X1 U66041 ( .A1(n73618), .A2(n106321), .B1(n80211), .B2(n110364), .ZN(
        n80956) );
  NAND2_X1 U66042 ( .A1(n80957), .A2(n80958), .ZN(n80954) );
  AOI22_X1 U66043 ( .A1(n73638), .A2(n106319), .B1(n73626), .B2(n80215), .ZN(
        n80958) );
  AOI22_X1 U66044 ( .A1(n73630), .A2(n106317), .B1(n80217), .B2(n110379), .ZN(
        n80957) );
  NAND2_X1 U66045 ( .A1(n80959), .A2(n80960), .ZN(n80953) );
  AOI22_X1 U66046 ( .A1(n106315), .A2(n110399), .B1(n80221), .B2(n110405), 
        .ZN(n80960) );
  AOI22_X1 U66047 ( .A1(n80222), .A2(n110386), .B1(n106312), .B2(n110391), 
        .ZN(n80959) );
  NAND2_X1 U66048 ( .A1(n80961), .A2(n80962), .ZN(n80952) );
  AOI22_X1 U66049 ( .A1(n106311), .A2(n110408), .B1(n73666), .B2(n106310), 
        .ZN(n80962) );
  AOI22_X1 U66050 ( .A1(n106309), .A2(n110395), .B1(n73654), .B2(n80229), .ZN(
        n80961) );
  NOR4_X1 U66051 ( .A1(n80963), .A2(n80964), .A3(n80965), .A4(n80966), .ZN(
        n80950) );
  OAI21_X1 U66052 ( .B1(n102005), .B2(n80234), .A(n80967), .ZN(n80966) );
  AOI22_X1 U66053 ( .A1(n73667), .A2(n106306), .B1(n73679), .B2(n106305), .ZN(
        n80967) );
  NAND2_X1 U66054 ( .A1(n80968), .A2(n80969), .ZN(n80965) );
  AOI22_X1 U66055 ( .A1(n106304), .A2(n110342), .B1(n80241), .B2(n110435), 
        .ZN(n80969) );
  AOI22_X1 U66056 ( .A1(n80242), .A2(n110424), .B1(n106301), .B2(n110432), 
        .ZN(n80968) );
  NAND2_X1 U66057 ( .A1(n80970), .A2(n80971), .ZN(n80964) );
  AOI22_X1 U66058 ( .A1(n106300), .A2(n110349), .B1(n73586), .B2(n106299), 
        .ZN(n80971) );
  AOI22_X1 U66059 ( .A1(n106298), .A2(n110353), .B1(n106297), .B2(n110340), 
        .ZN(n80970) );
  NAND2_X1 U66060 ( .A1(n80972), .A2(n80973), .ZN(n80963) );
  AOI22_X1 U66061 ( .A1(n80252), .A2(n110370), .B1(n80253), .B2(n110374), .ZN(
        n80973) );
  AOI22_X1 U66062 ( .A1(n106294), .A2(n110360), .B1(n73598), .B2(n106293), 
        .ZN(n80972) );
  NOR2_X1 U66063 ( .A1(n100572), .A2(n106292), .ZN(n80947) );
  AOI22_X1 U66064 ( .A1(n106291), .A2(n110416), .B1(n106290), .B2(n110428), 
        .ZN(n80945) );
  AOI22_X1 U66065 ( .A1(n73638), .A2(n105174), .B1(n73654), .B2(n105171), .ZN(
        n80944) );
  AOI22_X1 U66066 ( .A1(n80259), .A2(n110379), .B1(n73606), .B2(n106282), .ZN(
        n80943) );
  NAND4_X2 U66067 ( .A1(n80974), .A2(n80975), .A3(n80976), .A4(n80977), .ZN(
        n103981) );
  NOR3_X1 U66068 ( .A1(n80978), .A2(n80979), .A3(n80980), .ZN(n80977) );
  NOR2_X1 U66069 ( .A1(n100605), .A2(n106329), .ZN(n80980) );
  AOI21_X1 U66070 ( .B1(n80981), .B2(n80982), .A(n106324), .ZN(n80979) );
  NOR4_X1 U66071 ( .A1(n80983), .A2(n80984), .A3(n80985), .A4(n80986), .ZN(
        n80982) );
  OAI21_X1 U66072 ( .B1(n80208), .B2(n104624), .A(n80987), .ZN(n80986) );
  AOI22_X1 U66073 ( .A1(n73180), .A2(n106321), .B1(n80211), .B2(n110040), .ZN(
        n80987) );
  NAND2_X1 U66074 ( .A1(n80988), .A2(n80989), .ZN(n80985) );
  AOI22_X1 U66075 ( .A1(n73200), .A2(n106319), .B1(n73188), .B2(n80215), .ZN(
        n80989) );
  AOI22_X1 U66076 ( .A1(n73192), .A2(n106317), .B1(n80217), .B2(n110055), .ZN(
        n80988) );
  NAND2_X1 U66077 ( .A1(n80990), .A2(n80991), .ZN(n80984) );
  AOI22_X1 U66078 ( .A1(n106315), .A2(n110077), .B1(n80221), .B2(n110083), 
        .ZN(n80991) );
  AOI22_X1 U66079 ( .A1(n80222), .A2(n110064), .B1(n106312), .B2(n110069), 
        .ZN(n80990) );
  NAND2_X1 U66080 ( .A1(n80992), .A2(n80993), .ZN(n80983) );
  AOI22_X1 U66081 ( .A1(n106311), .A2(n110086), .B1(n73228), .B2(n106310), 
        .ZN(n80993) );
  AOI22_X1 U66082 ( .A1(n106309), .A2(n110073), .B1(n73216), .B2(n80229), .ZN(
        n80992) );
  NOR4_X1 U66083 ( .A1(n80994), .A2(n80995), .A3(n80996), .A4(n80997), .ZN(
        n80981) );
  OAI21_X1 U66084 ( .B1(n101987), .B2(n80234), .A(n80998), .ZN(n80997) );
  AOI22_X1 U66085 ( .A1(n73229), .A2(n106306), .B1(n73241), .B2(n106305), .ZN(
        n80998) );
  NAND2_X1 U66086 ( .A1(n80999), .A2(n81000), .ZN(n80996) );
  AOI22_X1 U66087 ( .A1(n106304), .A2(n110017), .B1(n106303), .B2(n110113), 
        .ZN(n81000) );
  AOI22_X1 U66088 ( .A1(n80242), .A2(n110102), .B1(n106301), .B2(n110110), 
        .ZN(n80999) );
  NAND2_X1 U66089 ( .A1(n81001), .A2(n81002), .ZN(n80995) );
  AOI22_X1 U66090 ( .A1(n106300), .A2(n110024), .B1(n73148), .B2(n106299), 
        .ZN(n81002) );
  AOI22_X1 U66091 ( .A1(n106298), .A2(n110028), .B1(n106297), .B2(n110015), 
        .ZN(n81001) );
  NAND2_X1 U66092 ( .A1(n81003), .A2(n81004), .ZN(n80994) );
  AOI22_X1 U66093 ( .A1(n80252), .A2(n110046), .B1(n80253), .B2(n110050), .ZN(
        n81004) );
  AOI22_X1 U66094 ( .A1(n106294), .A2(n110036), .B1(n73160), .B2(n106293), 
        .ZN(n81003) );
  NOR2_X1 U66095 ( .A1(n100573), .A2(n106292), .ZN(n80978) );
  AOI22_X1 U66096 ( .A1(n106291), .A2(n110094), .B1(n106290), .B2(n110106), 
        .ZN(n80976) );
  AOI22_X1 U66097 ( .A1(n73200), .A2(n105173), .B1(n73216), .B2(n105171), .ZN(
        n80975) );
  AOI22_X1 U66098 ( .A1(n80259), .A2(n110055), .B1(n73168), .B2(n80260), .ZN(
        n80974) );
  NAND4_X2 U66099 ( .A1(n81005), .A2(n81006), .A3(n81007), .A4(n81008), .ZN(
        n103982) );
  NOR3_X1 U66100 ( .A1(n81009), .A2(n81010), .A3(n81011), .ZN(n81008) );
  NOR2_X1 U66101 ( .A1(n100606), .A2(n106329), .ZN(n81011) );
  AOI21_X1 U66102 ( .B1(n81012), .B2(n81013), .A(n106325), .ZN(n81010) );
  NOR4_X1 U66103 ( .A1(n81014), .A2(n81015), .A3(n81016), .A4(n81017), .ZN(
        n81013) );
  OAI21_X1 U66104 ( .B1(n80208), .B2(n104623), .A(n81018), .ZN(n81017) );
  AOI22_X1 U66105 ( .A1(n73322), .A2(n106321), .B1(n80211), .B2(n110147), .ZN(
        n81018) );
  NAND2_X1 U66106 ( .A1(n81019), .A2(n81020), .ZN(n81016) );
  AOI22_X1 U66107 ( .A1(n73342), .A2(n106319), .B1(n73330), .B2(n80215), .ZN(
        n81020) );
  AOI22_X1 U66108 ( .A1(n73334), .A2(n106317), .B1(n80217), .B2(n110162), .ZN(
        n81019) );
  NAND2_X1 U66109 ( .A1(n81021), .A2(n81022), .ZN(n81015) );
  AOI22_X1 U66110 ( .A1(n106315), .A2(n110184), .B1(n80221), .B2(n110190), 
        .ZN(n81022) );
  AOI22_X1 U66111 ( .A1(n80222), .A2(n110171), .B1(n106312), .B2(n110176), 
        .ZN(n81021) );
  NAND2_X1 U66112 ( .A1(n81023), .A2(n81024), .ZN(n81014) );
  AOI22_X1 U66113 ( .A1(n106311), .A2(n110193), .B1(n73370), .B2(n106310), 
        .ZN(n81024) );
  AOI22_X1 U66114 ( .A1(n106309), .A2(n110180), .B1(n73358), .B2(n80229), .ZN(
        n81023) );
  NOR4_X1 U66115 ( .A1(n81025), .A2(n81026), .A3(n81027), .A4(n81028), .ZN(
        n81012) );
  OAI21_X1 U66116 ( .B1(n101971), .B2(n80234), .A(n81029), .ZN(n81028) );
  AOI22_X1 U66117 ( .A1(n73371), .A2(n106306), .B1(n73383), .B2(n106305), .ZN(
        n81029) );
  NAND2_X1 U66118 ( .A1(n81030), .A2(n81031), .ZN(n81027) );
  AOI22_X1 U66119 ( .A1(n106304), .A2(n110124), .B1(n106303), .B2(n110220), 
        .ZN(n81031) );
  AOI22_X1 U66120 ( .A1(n80242), .A2(n110209), .B1(n106301), .B2(n110217), 
        .ZN(n81030) );
  NAND2_X1 U66121 ( .A1(n81032), .A2(n81033), .ZN(n81026) );
  AOI22_X1 U66122 ( .A1(n106300), .A2(n110131), .B1(n73290), .B2(n106299), 
        .ZN(n81033) );
  AOI22_X1 U66123 ( .A1(n106298), .A2(n110135), .B1(n106297), .B2(n110122), 
        .ZN(n81032) );
  NAND2_X1 U66124 ( .A1(n81034), .A2(n81035), .ZN(n81025) );
  AOI22_X1 U66125 ( .A1(n80252), .A2(n110153), .B1(n80253), .B2(n110157), .ZN(
        n81035) );
  AOI22_X1 U66126 ( .A1(n106294), .A2(n110143), .B1(n73302), .B2(n106293), 
        .ZN(n81034) );
  NOR2_X1 U66127 ( .A1(n100574), .A2(n106292), .ZN(n81009) );
  AOI22_X1 U66128 ( .A1(n106291), .A2(n110201), .B1(n106290), .B2(n110213), 
        .ZN(n81007) );
  AOI22_X1 U66129 ( .A1(n73342), .A2(n106746), .B1(n73358), .B2(n106745), .ZN(
        n81006) );
  AOI22_X1 U66130 ( .A1(n106287), .A2(n110162), .B1(n73310), .B2(n106282), 
        .ZN(n81005) );
  NAND4_X2 U66131 ( .A1(n81036), .A2(n81037), .A3(n81038), .A4(n81039), .ZN(
        n103983) );
  NOR3_X1 U66132 ( .A1(n81040), .A2(n81041), .A3(n81042), .ZN(n81039) );
  NOR2_X1 U66133 ( .A1(n100607), .A2(n106329), .ZN(n81042) );
  AOI21_X1 U66134 ( .B1(n81043), .B2(n81044), .A(n106326), .ZN(n81041) );
  NOR4_X1 U66135 ( .A1(n81045), .A2(n81046), .A3(n81047), .A4(n81048), .ZN(
        n81044) );
  OAI21_X1 U66136 ( .B1(n80208), .B2(n104622), .A(n81049), .ZN(n81048) );
  AOI22_X1 U66137 ( .A1(n73038), .A2(n106321), .B1(n80211), .B2(n109931), .ZN(
        n81049) );
  NAND2_X1 U66138 ( .A1(n81050), .A2(n81051), .ZN(n81047) );
  AOI22_X1 U66139 ( .A1(n73058), .A2(n106319), .B1(n73046), .B2(n80215), .ZN(
        n81051) );
  AOI22_X1 U66140 ( .A1(n73050), .A2(n106317), .B1(n80217), .B2(n109946), .ZN(
        n81050) );
  NAND2_X1 U66141 ( .A1(n81052), .A2(n81053), .ZN(n81046) );
  AOI22_X1 U66142 ( .A1(n106315), .A2(n109969), .B1(n80221), .B2(n109975), 
        .ZN(n81053) );
  AOI22_X1 U66143 ( .A1(n80222), .A2(n109955), .B1(n106312), .B2(n109961), 
        .ZN(n81052) );
  NAND2_X1 U66144 ( .A1(n81054), .A2(n81055), .ZN(n81045) );
  AOI22_X1 U66145 ( .A1(n106311), .A2(n109978), .B1(n73086), .B2(n106310), 
        .ZN(n81055) );
  AOI22_X1 U66146 ( .A1(n106309), .A2(n109965), .B1(n73074), .B2(n80229), .ZN(
        n81054) );
  NOR4_X1 U66147 ( .A1(n81056), .A2(n81057), .A3(n81058), .A4(n81059), .ZN(
        n81043) );
  OAI21_X1 U66148 ( .B1(n101955), .B2(n80234), .A(n81060), .ZN(n81059) );
  AOI22_X1 U66149 ( .A1(n73087), .A2(n106306), .B1(n73099), .B2(n106305), .ZN(
        n81060) );
  NAND2_X1 U66150 ( .A1(n81061), .A2(n81062), .ZN(n81058) );
  AOI22_X1 U66151 ( .A1(n106304), .A2(n109908), .B1(n106303), .B2(n110005), 
        .ZN(n81062) );
  AOI22_X1 U66152 ( .A1(n80242), .A2(n109994), .B1(n106301), .B2(n110002), 
        .ZN(n81061) );
  NAND2_X1 U66153 ( .A1(n81063), .A2(n81064), .ZN(n81057) );
  AOI22_X1 U66154 ( .A1(n106300), .A2(n109915), .B1(n73006), .B2(n106299), 
        .ZN(n81064) );
  AOI22_X1 U66155 ( .A1(n106298), .A2(n109919), .B1(n106297), .B2(n109906), 
        .ZN(n81063) );
  NAND2_X1 U66156 ( .A1(n81065), .A2(n81066), .ZN(n81056) );
  AOI22_X1 U66157 ( .A1(n80252), .A2(n109937), .B1(n80253), .B2(n109941), .ZN(
        n81066) );
  AOI22_X1 U66158 ( .A1(n106294), .A2(n109927), .B1(n73018), .B2(n106293), 
        .ZN(n81065) );
  NOR2_X1 U66159 ( .A1(n100575), .A2(n106292), .ZN(n81040) );
  AOI22_X1 U66160 ( .A1(n106291), .A2(n109986), .B1(n106290), .B2(n109998), 
        .ZN(n81038) );
  AOI22_X1 U66161 ( .A1(n73058), .A2(n105173), .B1(n73074), .B2(n105172), .ZN(
        n81037) );
  AOI22_X1 U66162 ( .A1(n106287), .A2(n109946), .B1(n73026), .B2(n106282), 
        .ZN(n81036) );
  NAND4_X2 U66163 ( .A1(n81067), .A2(n81068), .A3(n81069), .A4(n81070), .ZN(
        n103984) );
  NOR3_X1 U66164 ( .A1(n81071), .A2(n81072), .A3(n81073), .ZN(n81070) );
  NOR2_X1 U66165 ( .A1(n100608), .A2(n106329), .ZN(n81073) );
  AOI21_X1 U66166 ( .B1(n81074), .B2(n81075), .A(n106323), .ZN(n81072) );
  NOR4_X1 U66167 ( .A1(n81076), .A2(n81077), .A3(n81078), .A4(n81079), .ZN(
        n81075) );
  OAI21_X1 U66168 ( .B1(n80208), .B2(n104621), .A(n81080), .ZN(n81079) );
  AOI22_X1 U66169 ( .A1(n72888), .A2(n106321), .B1(n80211), .B2(n109814), .ZN(
        n81080) );
  NAND2_X1 U66170 ( .A1(n81081), .A2(n81082), .ZN(n81078) );
  AOI22_X1 U66171 ( .A1(n72908), .A2(n106319), .B1(n72896), .B2(n80215), .ZN(
        n81082) );
  AOI22_X1 U66172 ( .A1(n72900), .A2(n106317), .B1(n80217), .B2(n109829), .ZN(
        n81081) );
  NAND2_X1 U66173 ( .A1(n81083), .A2(n81084), .ZN(n81077) );
  AOI22_X1 U66174 ( .A1(n106315), .A2(n109852), .B1(n80221), .B2(n109858), 
        .ZN(n81084) );
  AOI22_X1 U66175 ( .A1(n106313), .A2(n109838), .B1(n106312), .B2(n109844), 
        .ZN(n81083) );
  NAND2_X1 U66176 ( .A1(n81085), .A2(n81086), .ZN(n81076) );
  AOI22_X1 U66177 ( .A1(n106311), .A2(n109861), .B1(n72936), .B2(n106310), 
        .ZN(n81086) );
  AOI22_X1 U66178 ( .A1(n106309), .A2(n109848), .B1(n72924), .B2(n80229), .ZN(
        n81085) );
  NOR4_X1 U66179 ( .A1(n81087), .A2(n81088), .A3(n81089), .A4(n81090), .ZN(
        n81074) );
  OAI21_X1 U66180 ( .B1(n101939), .B2(n80234), .A(n81091), .ZN(n81090) );
  AOI22_X1 U66181 ( .A1(n72937), .A2(n106306), .B1(n72949), .B2(n106305), .ZN(
        n81091) );
  NAND2_X1 U66182 ( .A1(n81092), .A2(n81093), .ZN(n81089) );
  AOI22_X1 U66183 ( .A1(n106304), .A2(n109790), .B1(n106303), .B2(n109888), 
        .ZN(n81093) );
  AOI22_X1 U66184 ( .A1(n80242), .A2(n109877), .B1(n106301), .B2(n109885), 
        .ZN(n81092) );
  NAND2_X1 U66185 ( .A1(n81094), .A2(n81095), .ZN(n81088) );
  AOI22_X1 U66186 ( .A1(n106300), .A2(n109797), .B1(n72856), .B2(n106299), 
        .ZN(n81095) );
  AOI22_X1 U66187 ( .A1(n106298), .A2(n109801), .B1(n106297), .B2(n109788), 
        .ZN(n81094) );
  NAND2_X1 U66188 ( .A1(n81096), .A2(n81097), .ZN(n81087) );
  AOI22_X1 U66189 ( .A1(n80252), .A2(n109820), .B1(n80253), .B2(n109824), .ZN(
        n81097) );
  AOI22_X1 U66190 ( .A1(n106294), .A2(n109809), .B1(n72868), .B2(n106293), 
        .ZN(n81096) );
  NOR2_X1 U66191 ( .A1(n100576), .A2(n106292), .ZN(n81071) );
  AOI22_X1 U66192 ( .A1(n106291), .A2(n109869), .B1(n106290), .B2(n109881), 
        .ZN(n81069) );
  AOI22_X1 U66193 ( .A1(n72908), .A2(n105175), .B1(n72924), .B2(n106745), .ZN(
        n81068) );
  AOI22_X1 U66194 ( .A1(n106287), .A2(n109829), .B1(n72876), .B2(n106282), 
        .ZN(n81067) );
  NAND4_X2 U66195 ( .A1(n81098), .A2(n81099), .A3(n81100), .A4(n81101), .ZN(
        n103985) );
  NOR3_X1 U66196 ( .A1(n81102), .A2(n81103), .A3(n81104), .ZN(n81101) );
  NOR2_X1 U66197 ( .A1(n100609), .A2(n106329), .ZN(n81104) );
  AOI21_X1 U66198 ( .B1(n81105), .B2(n81106), .A(n106326), .ZN(n81103) );
  NOR4_X1 U66199 ( .A1(n81107), .A2(n81108), .A3(n81109), .A4(n81110), .ZN(
        n81106) );
  OAI21_X1 U66200 ( .B1(n80208), .B2(n104620), .A(n81111), .ZN(n81110) );
  AOI22_X1 U66201 ( .A1(n70784), .A2(n106321), .B1(n80211), .B2(n108188), .ZN(
        n81111) );
  NAND2_X1 U66202 ( .A1(n81112), .A2(n81113), .ZN(n81109) );
  AOI22_X1 U66203 ( .A1(n70804), .A2(n106319), .B1(n70792), .B2(n80215), .ZN(
        n81113) );
  AOI22_X1 U66204 ( .A1(n70796), .A2(n106317), .B1(n80217), .B2(n108203), .ZN(
        n81112) );
  NAND2_X1 U66205 ( .A1(n81114), .A2(n81115), .ZN(n81108) );
  AOI22_X1 U66206 ( .A1(n106315), .A2(n108226), .B1(n80221), .B2(n108232), 
        .ZN(n81115) );
  AOI22_X1 U66207 ( .A1(n80222), .A2(n108212), .B1(n106312), .B2(n108218), 
        .ZN(n81114) );
  NAND2_X1 U66208 ( .A1(n81116), .A2(n81117), .ZN(n81107) );
  AOI22_X1 U66209 ( .A1(n106311), .A2(n108235), .B1(n70832), .B2(n106310), 
        .ZN(n81117) );
  AOI22_X1 U66210 ( .A1(n106309), .A2(n108222), .B1(n70820), .B2(n80229), .ZN(
        n81116) );
  NOR4_X1 U66211 ( .A1(n81118), .A2(n81119), .A3(n81120), .A4(n81121), .ZN(
        n81105) );
  OAI21_X1 U66212 ( .B1(n101923), .B2(n80234), .A(n81122), .ZN(n81121) );
  AOI22_X1 U66213 ( .A1(n70833), .A2(n106306), .B1(n70845), .B2(n106305), .ZN(
        n81122) );
  NAND2_X1 U66214 ( .A1(n81123), .A2(n81124), .ZN(n81120) );
  AOI22_X1 U66215 ( .A1(n106304), .A2(n108164), .B1(n106303), .B2(n108262), 
        .ZN(n81124) );
  AOI22_X1 U66216 ( .A1(n80242), .A2(n108251), .B1(n106301), .B2(n108259), 
        .ZN(n81123) );
  NAND2_X1 U66217 ( .A1(n81125), .A2(n81126), .ZN(n81119) );
  AOI22_X1 U66218 ( .A1(n106300), .A2(n108171), .B1(n70752), .B2(n106299), 
        .ZN(n81126) );
  AOI22_X1 U66219 ( .A1(n106298), .A2(n108175), .B1(n106297), .B2(n108162), 
        .ZN(n81125) );
  NAND2_X1 U66220 ( .A1(n81127), .A2(n81128), .ZN(n81118) );
  AOI22_X1 U66221 ( .A1(n80252), .A2(n108194), .B1(n80253), .B2(n108198), .ZN(
        n81128) );
  AOI22_X1 U66222 ( .A1(n106294), .A2(n108183), .B1(n70764), .B2(n106293), 
        .ZN(n81127) );
  NOR2_X1 U66223 ( .A1(n100577), .A2(n106292), .ZN(n81102) );
  AOI22_X1 U66224 ( .A1(n106291), .A2(n108243), .B1(n106290), .B2(n108255), 
        .ZN(n81100) );
  AOI22_X1 U66225 ( .A1(n70804), .A2(n106746), .B1(n70820), .B2(n105170), .ZN(
        n81099) );
  AOI22_X1 U66226 ( .A1(n106287), .A2(n108203), .B1(n70772), .B2(n80260), .ZN(
        n81098) );
  NAND4_X2 U66227 ( .A1(n81129), .A2(n81130), .A3(n81131), .A4(n81132), .ZN(
        n103986) );
  NOR3_X1 U66228 ( .A1(n81133), .A2(n81134), .A3(n81135), .ZN(n81132) );
  NOR2_X1 U66229 ( .A1(n100610), .A2(n106329), .ZN(n81135) );
  AOI21_X1 U66230 ( .B1(n81136), .B2(n81137), .A(n106323), .ZN(n81134) );
  NOR4_X1 U66231 ( .A1(n81138), .A2(n81139), .A3(n81140), .A4(n81141), .ZN(
        n81137) );
  OAI21_X1 U66232 ( .B1(n80208), .B2(n104619), .A(n81142), .ZN(n81141) );
  AOI22_X1 U66233 ( .A1(n70943), .A2(n106321), .B1(n80211), .B2(n108311), .ZN(
        n81142) );
  NAND2_X1 U66234 ( .A1(n81143), .A2(n81144), .ZN(n81140) );
  AOI22_X1 U66235 ( .A1(n70963), .A2(n106319), .B1(n70951), .B2(n80215), .ZN(
        n81144) );
  AOI22_X1 U66236 ( .A1(n70955), .A2(n106317), .B1(n80217), .B2(n108326), .ZN(
        n81143) );
  NAND2_X1 U66237 ( .A1(n81145), .A2(n81146), .ZN(n81139) );
  AOI22_X1 U66238 ( .A1(n106315), .A2(n108349), .B1(n80221), .B2(n108355), 
        .ZN(n81146) );
  AOI22_X1 U66239 ( .A1(n106313), .A2(n108335), .B1(n106312), .B2(n108341), 
        .ZN(n81145) );
  NAND2_X1 U66240 ( .A1(n81147), .A2(n81148), .ZN(n81138) );
  AOI22_X1 U66241 ( .A1(n106311), .A2(n108358), .B1(n70991), .B2(n106310), 
        .ZN(n81148) );
  AOI22_X1 U66242 ( .A1(n106309), .A2(n108345), .B1(n70979), .B2(n80229), .ZN(
        n81147) );
  NOR4_X1 U66243 ( .A1(n81149), .A2(n81150), .A3(n81151), .A4(n81152), .ZN(
        n81136) );
  OAI21_X1 U66244 ( .B1(n101907), .B2(n80234), .A(n81153), .ZN(n81152) );
  AOI22_X1 U66245 ( .A1(n70992), .A2(n106306), .B1(n71004), .B2(n106305), .ZN(
        n81153) );
  NAND2_X1 U66246 ( .A1(n81154), .A2(n81155), .ZN(n81151) );
  AOI22_X1 U66247 ( .A1(n106304), .A2(n108287), .B1(n106303), .B2(n108385), 
        .ZN(n81155) );
  AOI22_X1 U66248 ( .A1(n80242), .A2(n108374), .B1(n106301), .B2(n108382), 
        .ZN(n81154) );
  NAND2_X1 U66249 ( .A1(n81156), .A2(n81157), .ZN(n81150) );
  AOI22_X1 U66250 ( .A1(n106300), .A2(n108294), .B1(n70911), .B2(n106299), 
        .ZN(n81157) );
  AOI22_X1 U66251 ( .A1(n106298), .A2(n108298), .B1(n106297), .B2(n108285), 
        .ZN(n81156) );
  NAND2_X1 U66252 ( .A1(n81158), .A2(n81159), .ZN(n81149) );
  AOI22_X1 U66253 ( .A1(n80252), .A2(n108317), .B1(n80253), .B2(n108321), .ZN(
        n81159) );
  AOI22_X1 U66254 ( .A1(n106294), .A2(n108306), .B1(n70923), .B2(n106293), 
        .ZN(n81158) );
  NOR2_X1 U66255 ( .A1(n100578), .A2(n106292), .ZN(n81133) );
  AOI22_X1 U66256 ( .A1(n106291), .A2(n108366), .B1(n106290), .B2(n108378), 
        .ZN(n81131) );
  AOI22_X1 U66257 ( .A1(n70963), .A2(n105173), .B1(n70979), .B2(n105171), .ZN(
        n81130) );
  AOI22_X1 U66258 ( .A1(n106287), .A2(n108326), .B1(n70931), .B2(n106283), 
        .ZN(n81129) );
  NAND4_X2 U66259 ( .A1(n81160), .A2(n81161), .A3(n81162), .A4(n81163), .ZN(
        n103987) );
  NOR3_X1 U66260 ( .A1(n81164), .A2(n81165), .A3(n81166), .ZN(n81163) );
  NOR2_X1 U66261 ( .A1(n100611), .A2(n106329), .ZN(n81166) );
  AOI21_X1 U66262 ( .B1(n81167), .B2(n81168), .A(n106324), .ZN(n81165) );
  NOR4_X1 U66263 ( .A1(n81169), .A2(n81170), .A3(n81171), .A4(n81172), .ZN(
        n81168) );
  OAI21_X1 U66264 ( .B1(n80208), .B2(n104618), .A(n81173), .ZN(n81172) );
  AOI22_X1 U66265 ( .A1(n71088), .A2(n106321), .B1(n80211), .B2(n108422), .ZN(
        n81173) );
  NAND2_X1 U66266 ( .A1(n81174), .A2(n81175), .ZN(n81171) );
  AOI22_X1 U66267 ( .A1(n71108), .A2(n106319), .B1(n71096), .B2(n80215), .ZN(
        n81175) );
  AOI22_X1 U66268 ( .A1(n71100), .A2(n106317), .B1(n80217), .B2(n108437), .ZN(
        n81174) );
  NAND2_X1 U66269 ( .A1(n81176), .A2(n81177), .ZN(n81170) );
  AOI22_X1 U66270 ( .A1(n106315), .A2(n108460), .B1(n80221), .B2(n108466), 
        .ZN(n81177) );
  AOI22_X1 U66271 ( .A1(n80222), .A2(n108446), .B1(n106312), .B2(n108452), 
        .ZN(n81176) );
  NAND2_X1 U66272 ( .A1(n81178), .A2(n81179), .ZN(n81169) );
  AOI22_X1 U66273 ( .A1(n106311), .A2(n108469), .B1(n71136), .B2(n106310), 
        .ZN(n81179) );
  AOI22_X1 U66274 ( .A1(n106309), .A2(n108456), .B1(n71124), .B2(n80229), .ZN(
        n81178) );
  NOR4_X1 U66275 ( .A1(n81180), .A2(n81181), .A3(n81182), .A4(n81183), .ZN(
        n81167) );
  OAI21_X1 U66276 ( .B1(n101891), .B2(n80234), .A(n81184), .ZN(n81183) );
  AOI22_X1 U66277 ( .A1(n71137), .A2(n106306), .B1(n71149), .B2(n106305), .ZN(
        n81184) );
  NAND2_X1 U66278 ( .A1(n81185), .A2(n81186), .ZN(n81182) );
  AOI22_X1 U66279 ( .A1(n106304), .A2(n108398), .B1(n106303), .B2(n108496), 
        .ZN(n81186) );
  AOI22_X1 U66280 ( .A1(n80242), .A2(n108485), .B1(n106301), .B2(n108493), 
        .ZN(n81185) );
  NAND2_X1 U66281 ( .A1(n81187), .A2(n81188), .ZN(n81181) );
  AOI22_X1 U66282 ( .A1(n106300), .A2(n108405), .B1(n71056), .B2(n106299), 
        .ZN(n81188) );
  AOI22_X1 U66283 ( .A1(n106298), .A2(n108409), .B1(n106297), .B2(n108396), 
        .ZN(n81187) );
  NAND2_X1 U66284 ( .A1(n81189), .A2(n81190), .ZN(n81180) );
  AOI22_X1 U66285 ( .A1(n80252), .A2(n108428), .B1(n80253), .B2(n108432), .ZN(
        n81190) );
  AOI22_X1 U66286 ( .A1(n106294), .A2(n108417), .B1(n71068), .B2(n106293), 
        .ZN(n81189) );
  NOR2_X1 U66287 ( .A1(n100579), .A2(n106292), .ZN(n81164) );
  AOI22_X1 U66288 ( .A1(n106291), .A2(n108477), .B1(n106290), .B2(n108489), 
        .ZN(n81162) );
  AOI22_X1 U66289 ( .A1(n71108), .A2(n105174), .B1(n71124), .B2(n105172), .ZN(
        n81161) );
  AOI22_X1 U66290 ( .A1(n106287), .A2(n108437), .B1(n71076), .B2(n106282), 
        .ZN(n81160) );
  NAND4_X2 U66291 ( .A1(n81191), .A2(n81192), .A3(n81193), .A4(n81194), .ZN(
        n103988) );
  NOR3_X1 U66292 ( .A1(n81195), .A2(n81196), .A3(n81197), .ZN(n81194) );
  NOR2_X1 U66293 ( .A1(n100612), .A2(n106329), .ZN(n81197) );
  AOI21_X1 U66294 ( .B1(n106744), .B2(n81198), .A(n105100), .ZN(n80200) );
  AOI21_X1 U66295 ( .B1(n81200), .B2(n81201), .A(n106325), .ZN(n81196) );
  NOR4_X1 U66296 ( .A1(n81202), .A2(n81203), .A3(n81204), .A4(n81205), .ZN(
        n81201) );
  OAI21_X1 U66297 ( .B1(n80208), .B2(n104617), .A(n81206), .ZN(n81205) );
  AOI22_X1 U66298 ( .A1(n70049), .A2(n106321), .B1(n106320), .B2(n107660), 
        .ZN(n81206) );
  NOR2_X1 U66299 ( .A1(n81207), .A2(n81208), .ZN(n80211) );
  NOR2_X1 U66300 ( .A1(n81207), .A2(n106278), .ZN(n80210) );
  NAND2_X1 U66301 ( .A1(n81210), .A2(n81211), .ZN(n80208) );
  NAND2_X1 U66302 ( .A1(n81212), .A2(n81213), .ZN(n81204) );
  AOI22_X1 U66303 ( .A1(n70069), .A2(n106319), .B1(n70057), .B2(n106318), .ZN(
        n81213) );
  NOR2_X1 U66304 ( .A1(n81207), .A2(n107026), .ZN(n80215) );
  NOR2_X1 U66305 ( .A1(n107024), .A2(n81214), .ZN(n80214) );
  AOI22_X1 U66306 ( .A1(n70061), .A2(n106317), .B1(n106316), .B2(n107675), 
        .ZN(n81212) );
  NOR2_X1 U66307 ( .A1(n106742), .A2(n107026), .ZN(n80217) );
  NOR2_X1 U66308 ( .A1(n81208), .A2(n81214), .ZN(n80216) );
  NAND2_X1 U66309 ( .A1(n81215), .A2(n81216), .ZN(n81203) );
  AOI22_X1 U66310 ( .A1(n106315), .A2(n107698), .B1(n106314), .B2(n107704), 
        .ZN(n81216) );
  NOR2_X1 U66311 ( .A1(n81217), .A2(n107026), .ZN(n80221) );
  NOR2_X1 U66312 ( .A1(n81217), .A2(n106278), .ZN(n80220) );
  AOI22_X1 U66313 ( .A1(n106313), .A2(n107684), .B1(n106312), .B2(n107690), 
        .ZN(n81215) );
  NOR2_X1 U66314 ( .A1(n107024), .A2(n81217), .ZN(n80223) );
  NOR2_X1 U66315 ( .A1(n81208), .A2(n81217), .ZN(n80222) );
  NAND2_X1 U66316 ( .A1(n81218), .A2(n105056), .ZN(n81217) );
  NOR2_X1 U66317 ( .A1(n62190), .A2(n106697), .ZN(n81218) );
  NAND2_X1 U66318 ( .A1(n81219), .A2(n81220), .ZN(n81202) );
  AOI22_X1 U66319 ( .A1(n106311), .A2(n107707), .B1(n70097), .B2(n106310), 
        .ZN(n81220) );
  NOR2_X1 U66320 ( .A1(n81221), .A2(n62190), .ZN(n80227) );
  NOR2_X1 U66321 ( .A1(n81221), .A2(n104582), .ZN(n80226) );
  AOI22_X1 U66322 ( .A1(n106309), .A2(n107694), .B1(n70085), .B2(n106308), 
        .ZN(n81219) );
  NOR2_X1 U66323 ( .A1(n107026), .A2(n81214), .ZN(n80229) );
  NOR2_X1 U66324 ( .A1(n81214), .A2(n106278), .ZN(n80228) );
  NAND2_X1 U66325 ( .A1(n81222), .A2(n105056), .ZN(n81214) );
  NOR2_X1 U66326 ( .A1(n104582), .A2(n106697), .ZN(n81222) );
  NOR4_X1 U66327 ( .A1(n81223), .A2(n81224), .A3(n81225), .A4(n81226), .ZN(
        n81200) );
  OAI21_X1 U66328 ( .B1(n101875), .B2(n80234), .A(n81227), .ZN(n81226) );
  AOI22_X1 U66329 ( .A1(n70098), .A2(n106306), .B1(n70110), .B2(n106305), .ZN(
        n81227) );
  NOR2_X1 U66330 ( .A1(n81228), .A2(n106743), .ZN(n80237) );
  NOR2_X1 U66331 ( .A1(n81229), .A2(n106743), .ZN(n80236) );
  NAND2_X1 U66332 ( .A1(n104582), .A2(n81230), .ZN(n81229) );
  NAND2_X1 U66333 ( .A1(n81231), .A2(n81232), .ZN(n80234) );
  NOR2_X1 U66334 ( .A1(n62190), .A2(n106278), .ZN(n81231) );
  NAND2_X1 U66335 ( .A1(n81233), .A2(n81234), .ZN(n81225) );
  AOI22_X1 U66336 ( .A1(n106304), .A2(n107636), .B1(n106303), .B2(n107733), 
        .ZN(n81234) );
  NOR2_X1 U66337 ( .A1(n81235), .A2(n104582), .ZN(n80241) );
  NOR2_X1 U66338 ( .A1(n81236), .A2(n81208), .ZN(n80240) );
  AOI22_X1 U66339 ( .A1(n106302), .A2(n107722), .B1(n106301), .B2(n107730), 
        .ZN(n81233) );
  NOR2_X1 U66340 ( .A1(n81235), .A2(n62190), .ZN(n80243) );
  NAND2_X1 U66343 ( .A1(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ), 
        .A2(n81238), .ZN(n81221) );
  NOR2_X1 U66344 ( .A1(n81239), .A2(n106743), .ZN(n80242) );
  NAND2_X1 U66345 ( .A1(n104582), .A2(n81211), .ZN(n81239) );
  NAND2_X1 U66346 ( .A1(n81240), .A2(n81241), .ZN(n81224) );
  AOI22_X1 U66347 ( .A1(n106300), .A2(n107643), .B1(n70017), .B2(n106299), 
        .ZN(n81241) );
  NOR2_X1 U66348 ( .A1(n81236), .A2(n106278), .ZN(n80247) );
  NOR2_X1 U66349 ( .A1(n81236), .A2(n107024), .ZN(n80246) );
  AOI22_X1 U66350 ( .A1(n106298), .A2(n107647), .B1(n106297), .B2(n107634), 
        .ZN(n81240) );
  NOR2_X1 U66351 ( .A1(n81242), .A2(n81208), .ZN(n80249) );
  NOR2_X1 U66352 ( .A1(n81242), .A2(n106278), .ZN(n80248) );
  NAND2_X1 U66353 ( .A1(n81243), .A2(n81244), .ZN(n81223) );
  AOI22_X1 U66354 ( .A1(n106296), .A2(n107666), .B1(n106295), .B2(n107670), 
        .ZN(n81244) );
  NOR2_X1 U66355 ( .A1(n106742), .A2(n106278), .ZN(n80253) );
  NOR2_X1 U66356 ( .A1(n81207), .A2(n107024), .ZN(n80252) );
  AOI22_X1 U66359 ( .A1(n106294), .A2(n107655), .B1(n70029), .B2(n106293), 
        .ZN(n81243) );
  NOR2_X1 U66360 ( .A1(n106742), .A2(n81208), .ZN(n80255) );
  NOR2_X1 U66363 ( .A1(n81236), .A2(n107026), .ZN(n80254) );
  NAND2_X1 U66364 ( .A1(n81248), .A2(n105056), .ZN(n81236) );
  NOR2_X1 U66365 ( .A1(n62190), .A2(n81247), .ZN(n81248) );
  NOR2_X1 U66366 ( .A1(n100580), .A2(n106292), .ZN(n81195) );
  AOI21_X1 U66367 ( .B1(n106744), .B2(n81249), .A(n106275), .ZN(n80256) );
  NAND2_X1 U66368 ( .A1(n81251), .A2(n105056), .ZN(n81242) );
  NOR2_X1 U66369 ( .A1(n81247), .A2(n104582), .ZN(n81251) );
  AOI22_X1 U66370 ( .A1(n106291), .A2(n107714), .B1(n106290), .B2(n107726), 
        .ZN(n81193) );
  OAI21_X1 U66371 ( .B1(n106743), .B2(n81252), .A(n81253), .ZN(n80258) );
  OAI21_X1 U66372 ( .B1(n106743), .B2(n81254), .A(n106761), .ZN(n80257) );
  NOR2_X1 U66373 ( .A1(n81247), .A2(n105056), .ZN(n81232) );
  XOR2_X1 U66374 ( .A(n81238), .B(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ), 
        .Z(n81247) );
  AOI22_X1 U66375 ( .A1(n70069), .A2(n106746), .B1(n70085), .B2(n106745), .ZN(
        n81192) );
  AOI22_X1 U66376 ( .A1(n106287), .A2(n107675), .B1(n70037), .B2(n80260), .ZN(
        n81191) );
  OAI21_X1 U66377 ( .B1(n109055), .B2(n81256), .A(n81257), .ZN(n103989) );
  AOI22_X1 U66378 ( .A1(n81258), .A2(n81259), .B1(n106012), .B2(n81260), .ZN(
        n81257) );
  OAI21_X1 U66379 ( .B1(n106271), .B2(n81262), .A(n81263), .ZN(n103990) );
  AOI22_X1 U66380 ( .A1(n106265), .A2(n107355), .B1(n81265), .B2(n104879), 
        .ZN(n81263) );
  OAI21_X1 U66381 ( .B1(n106271), .B2(n81267), .A(n81268), .ZN(n103991) );
  AOI22_X1 U66382 ( .A1(n106265), .A2(n109391), .B1(n81269), .B2(n104879), 
        .ZN(n81268) );
  OAI21_X1 U66383 ( .B1(n106272), .B2(n81270), .A(n81271), .ZN(n103992) );
  AOI22_X1 U66384 ( .A1(n106265), .A2(n110813), .B1(n81272), .B2(n104880), 
        .ZN(n81271) );
  OAI21_X1 U66385 ( .B1(n106266), .B2(n106253), .A(n81274), .ZN(n103993) );
  AOI22_X1 U66386 ( .A1(n69683), .A2(n106251), .B1(n106249), .B2(n81265), .ZN(
        n81274) );
  OAI21_X1 U66387 ( .B1(n106261), .B2(n106253), .A(n81277), .ZN(n103994) );
  AOI22_X1 U66388 ( .A1(n72316), .A2(n106250), .B1(n106249), .B2(n81269), .ZN(
        n81277) );
  OAI21_X1 U66389 ( .B1(n106253), .B2(n81278), .A(n81279), .ZN(n103995) );
  AOI22_X1 U66390 ( .A1(n71274), .A2(n106250), .B1(n106242), .B2(n106249), 
        .ZN(n81279) );
  OAI21_X1 U66391 ( .B1(n106252), .B2(n81281), .A(n81282), .ZN(n103996) );
  AOI22_X1 U66392 ( .A1(n71125), .A2(n106251), .B1(n81283), .B2(n106248), .ZN(
        n81282) );
  OAI21_X1 U66393 ( .B1(n106253), .B2(n81284), .A(n81285), .ZN(n103997) );
  AOI22_X1 U66394 ( .A1(n70821), .A2(n106250), .B1(n81286), .B2(n106249), .ZN(
        n81285) );
  OAI21_X1 U66395 ( .B1(n107127), .B2(n106253), .A(n81287), .ZN(n103998) );
  AOI22_X1 U66396 ( .A1(n71574), .A2(n106251), .B1(n106249), .B2(n80188), .ZN(
        n81287) );
  OAI21_X1 U66397 ( .B1(n81267), .B2(n106229), .A(n81289), .ZN(n103999) );
  AOI22_X1 U66398 ( .A1(n106228), .A2(n81269), .B1(n106225), .B2(n109383), 
        .ZN(n81289) );
  OAI21_X1 U66399 ( .B1(n106235), .B2(n106229), .A(n81292), .ZN(n104000) );
  AOI22_X1 U66400 ( .A1(n106227), .A2(n81283), .B1(n106224), .B2(n108453), 
        .ZN(n81292) );
  OAI21_X1 U66401 ( .B1(n106223), .B2(n106219), .A(n81295), .ZN(n104001) );
  AOI22_X1 U66402 ( .A1(n106217), .A2(n109966), .B1(n81297), .B2(n106214), 
        .ZN(n81295) );
  OAI21_X1 U66403 ( .B1(n106223), .B2(n106209), .A(n81300), .ZN(n104002) );
  AOI22_X1 U66404 ( .A1(n106216), .A2(n107811), .B1(n81301), .B2(n106214), 
        .ZN(n81300) );
  OAI21_X1 U66405 ( .B1(n107127), .B2(n106229), .A(n81302), .ZN(n104003) );
  AOI22_X1 U66406 ( .A1(n106227), .A2(n80188), .B1(n106224), .B2(n108807), 
        .ZN(n81302) );
  OAI21_X1 U66407 ( .B1(n81278), .B2(n106229), .A(n81303), .ZN(n104004) );
  AOI22_X1 U66408 ( .A1(n106228), .A2(n106240), .B1(n71262), .B2(n106224), 
        .ZN(n81303) );
  OAI21_X1 U66409 ( .B1(n81284), .B2(n106229), .A(n81304), .ZN(n104005) );
  AOI22_X1 U66410 ( .A1(n106227), .A2(n81286), .B1(n106224), .B2(n108219), 
        .ZN(n81304) );
  OAI21_X1 U66411 ( .B1(n106254), .B2(n106229), .A(n81305), .ZN(n104006) );
  AOI22_X1 U66412 ( .A1(n106228), .A2(n81272), .B1(n106224), .B2(n110806), 
        .ZN(n81305) );
  OAI21_X1 U66413 ( .B1(n106229), .B2(n106205), .A(n81307), .ZN(n104007) );
  AOI22_X1 U66414 ( .A1(n81308), .A2(n106227), .B1(n106224), .B2(n110704), 
        .ZN(n81307) );
  OAI21_X1 U66415 ( .B1(n106202), .B2(n81310), .A(n81311), .ZN(n104008) );
  AOI22_X1 U66416 ( .A1(n106195), .A2(n81313), .B1(n81314), .B2(n109612), .ZN(
        n81311) );
  OAI21_X1 U66417 ( .B1(n106202), .B2(n81315), .A(n81316), .ZN(n104009) );
  AOI22_X1 U66418 ( .A1(n81317), .A2(n106196), .B1(n81314), .B2(n110289), .ZN(
        n81316) );
  OAI21_X1 U66419 ( .B1(n106202), .B2(n81318), .A(n81319), .ZN(n104010) );
  AOI22_X1 U66420 ( .A1(n81320), .A2(n106195), .B1(n81314), .B2(n110398), .ZN(
        n81319) );
  OAI21_X1 U66421 ( .B1(n106235), .B2(n106202), .A(n81321), .ZN(n104011) );
  AOI22_X1 U66422 ( .A1(n81322), .A2(n106196), .B1(n81314), .B2(n108459), .ZN(
        n81321) );
  OAI21_X1 U66423 ( .B1(n106266), .B2(n106183), .A(n81324), .ZN(n104012) );
  AOI22_X1 U66424 ( .A1(n106182), .A2(n107357), .B1(n104882), .B2(n81327), 
        .ZN(n81324) );
  OAI21_X1 U66425 ( .B1(n106235), .B2(n106184), .A(n81328), .ZN(n104013) );
  AOI22_X1 U66426 ( .A1(n81325), .A2(n108463), .B1(n104881), .B2(n81322), .ZN(
        n81328) );
  OAI21_X1 U66427 ( .B1(n106244), .B2(n106184), .A(n81329), .ZN(n104014) );
  AOI22_X1 U66428 ( .A1(n81325), .A2(n108578), .B1(n81330), .B2(n104882), .ZN(
        n81329) );
  OAI21_X1 U66429 ( .B1(n81284), .B2(n106184), .A(n81331), .ZN(n104015) );
  AOI22_X1 U66430 ( .A1(n106182), .A2(n108229), .B1(n81332), .B2(n104881), 
        .ZN(n81331) );
  OAI21_X1 U66431 ( .B1(n81318), .B2(n106184), .A(n81333), .ZN(n104016) );
  AOI22_X1 U66432 ( .A1(n106182), .A2(n110402), .B1(n81326), .B2(n81320), .ZN(
        n81333) );
  OAI21_X1 U66433 ( .B1(n107127), .B2(n106184), .A(n81334), .ZN(n104017) );
  AOI22_X1 U66434 ( .A1(n81325), .A2(n108817), .B1(n81335), .B2(n81326), .ZN(
        n81334) );
  OAI21_X1 U66435 ( .B1(n106235), .B2(n106180), .A(n81337), .ZN(n104018) );
  AOI22_X1 U66436 ( .A1(n106178), .A2(n81283), .B1(n106175), .B2(n108441), 
        .ZN(n81337) );
  OAI21_X1 U66437 ( .B1(n106179), .B2(n106173), .A(n81341), .ZN(n104019) );
  AOI22_X1 U66438 ( .A1(n106167), .A2(n106178), .B1(n81339), .B2(n108330), 
        .ZN(n81341) );
  OAI21_X1 U66439 ( .B1(n106230), .B2(n106180), .A(n81343), .ZN(n104020) );
  AOI22_X1 U66440 ( .A1(n106178), .A2(n81286), .B1(n106176), .B2(n108207), 
        .ZN(n81343) );
  OAI21_X1 U66441 ( .B1(n106218), .B2(n106180), .A(n81344), .ZN(n104021) );
  AOI22_X1 U66442 ( .A1(n106178), .A2(n81297), .B1(n106175), .B2(n109950), 
        .ZN(n81344) );
  OAI21_X1 U66443 ( .B1(n106180), .B2(n106164), .A(n81346), .ZN(n104022) );
  AOI22_X1 U66444 ( .A1(n81347), .A2(n106177), .B1(n81339), .B2(n110059), .ZN(
        n81346) );
  OAI21_X1 U66445 ( .B1(n107127), .B2(n106180), .A(n81348), .ZN(n104023) );
  AOI22_X1 U66446 ( .A1(n106178), .A2(n80188), .B1(n81339), .B2(n108795), .ZN(
        n81348) );
  OAI21_X1 U66447 ( .B1(n106179), .B2(n106159), .A(n81350), .ZN(n104024) );
  AOI22_X1 U66448 ( .A1(n81351), .A2(n106178), .B1(n81339), .B2(n109702), .ZN(
        n81350) );
  OAI21_X1 U66449 ( .B1(n81299), .B2(n106180), .A(n81352), .ZN(n104025) );
  AOI22_X1 U66450 ( .A1(n106178), .A2(n81301), .B1(n106175), .B2(n107796), 
        .ZN(n81352) );
  OAI21_X1 U66451 ( .B1(n106259), .B2(n106156), .A(n81354), .ZN(n104026) );
  AOI22_X1 U66452 ( .A1(n106153), .A2(n109377), .B1(n106151), .B2(n81269), 
        .ZN(n81354) );
  OAI21_X1 U66453 ( .B1(n106243), .B2(n106156), .A(n81357), .ZN(n104027) );
  AOI22_X1 U66454 ( .A1(n81355), .A2(n108564), .B1(n106152), .B2(n106242), 
        .ZN(n81357) );
  OAI21_X1 U66455 ( .B1(n106155), .B2(n106148), .A(n81359), .ZN(n104028) );
  AOI22_X1 U66456 ( .A1(n70363), .A2(n106154), .B1(n81360), .B2(n81356), .ZN(
        n81359) );
  OAI21_X1 U66457 ( .B1(n106235), .B2(n106156), .A(n81361), .ZN(n104029) );
  AOI22_X1 U66458 ( .A1(n81355), .A2(n108447), .B1(n106152), .B2(n81283), .ZN(
        n81361) );
  OAI21_X1 U66459 ( .B1(n81340), .B2(n106156), .A(n81362), .ZN(n104030) );
  AOI22_X1 U66460 ( .A1(n106153), .A2(n108336), .B1(n106152), .B2(n106168), 
        .ZN(n81362) );
  OAI21_X1 U66461 ( .B1(n106231), .B2(n106156), .A(n81363), .ZN(n104031) );
  AOI22_X1 U66462 ( .A1(n81355), .A2(n108213), .B1(n106152), .B2(n81286), .ZN(
        n81363) );
  OAI21_X1 U66463 ( .B1(n107127), .B2(n106156), .A(n81364), .ZN(n104032) );
  AOI22_X1 U66464 ( .A1(n81355), .A2(n108801), .B1(n106152), .B2(n80188), .ZN(
        n81364) );
  OAI21_X1 U66465 ( .B1(n81349), .B2(n106156), .A(n81365), .ZN(n104033) );
  AOI22_X1 U66466 ( .A1(n106153), .A2(n109708), .B1(n106152), .B2(n81351), 
        .ZN(n81365) );
  OAI21_X1 U66467 ( .B1(n106208), .B2(n106156), .A(n81366), .ZN(n104034) );
  AOI22_X1 U66468 ( .A1(n81355), .A2(n107802), .B1(n106152), .B2(n81301), .ZN(
        n81366) );
  OAI21_X1 U66469 ( .B1(n106235), .B2(n106144), .A(n81368), .ZN(n104035) );
  AOI22_X1 U66470 ( .A1(n106143), .A2(n108443), .B1(n106141), .B2(n81322), 
        .ZN(n81368) );
  OAI21_X1 U66471 ( .B1(n81284), .B2(n106144), .A(n81371), .ZN(n104036) );
  AOI22_X1 U66472 ( .A1(n106143), .A2(n108209), .B1(n106140), .B2(n81332), 
        .ZN(n81371) );
  OAI21_X1 U66473 ( .B1(n81340), .B2(n106144), .A(n81372), .ZN(n104037) );
  AOI22_X1 U66474 ( .A1(n106143), .A2(n108332), .B1(n81373), .B2(n106140), 
        .ZN(n81372) );
  OAI21_X1 U66475 ( .B1(n106245), .B2(n106144), .A(n81374), .ZN(n104038) );
  AOI22_X1 U66476 ( .A1(n106143), .A2(n108560), .B1(n106141), .B2(n81330), 
        .ZN(n81374) );
  OAI21_X1 U66477 ( .B1(n81310), .B2(n106144), .A(n81375), .ZN(n104039) );
  AOI22_X1 U66478 ( .A1(n106143), .A2(n109599), .B1(n106140), .B2(n81313), 
        .ZN(n81375) );
  OAI21_X1 U66479 ( .B1(n81299), .B2(n106144), .A(n81376), .ZN(n104040) );
  AOI22_X1 U66480 ( .A1(n106143), .A2(n107798), .B1(n81377), .B2(n106141), 
        .ZN(n81376) );
  OAI21_X1 U66481 ( .B1(n106145), .B2(n81378), .A(n81379), .ZN(n104041) );
  AOI22_X1 U66482 ( .A1(n106143), .A2(n107261), .B1(n81380), .B2(n106140), 
        .ZN(n81379) );
  OAI21_X1 U66483 ( .B1(n105220), .B2(n106144), .A(n81381), .ZN(n104042) );
  AOI22_X1 U66484 ( .A1(n106143), .A2(n108797), .B1(n106140), .B2(n81335), 
        .ZN(n81381) );
  OAI21_X1 U66485 ( .B1(n106134), .B2(n81383), .A(n81384), .ZN(n104043) );
  AOI22_X1 U66486 ( .A1(n106127), .A2(n81386), .B1(n106124), .B2(n110595), 
        .ZN(n81384) );
  OAI21_X1 U66487 ( .B1(n106235), .B2(n106122), .A(n81389), .ZN(n104044) );
  AOI22_X1 U66488 ( .A1(n71107), .A2(n106121), .B1(n106118), .B2(n81322), .ZN(
        n81389) );
  OAI21_X1 U66489 ( .B1(n81284), .B2(n106122), .A(n81392), .ZN(n104045) );
  AOI22_X1 U66490 ( .A1(n70803), .A2(n106121), .B1(n106118), .B2(n81332), .ZN(
        n81392) );
  OAI21_X1 U66491 ( .B1(n81340), .B2(n106122), .A(n81393), .ZN(n104046) );
  AOI22_X1 U66492 ( .A1(n70962), .A2(n106121), .B1(n106119), .B2(n81373), .ZN(
        n81393) );
  OAI21_X1 U66493 ( .B1(n106122), .B2(n106114), .A(n81395), .ZN(n104047) );
  AOI22_X1 U66494 ( .A1(n72449), .A2(n106121), .B1(n81396), .B2(n106118), .ZN(
        n81395) );
  OAI21_X1 U66495 ( .B1(n81310), .B2(n106122), .A(n81397), .ZN(n104048) );
  AOI22_X1 U66496 ( .A1(n72597), .A2(n106121), .B1(n106118), .B2(n81313), .ZN(
        n81397) );
  OAI21_X1 U66497 ( .B1(n106123), .B2(n106110), .A(n81399), .ZN(n104049) );
  AOI22_X1 U66498 ( .A1(n72907), .A2(n106121), .B1(n81400), .B2(n106119), .ZN(
        n81399) );
  OAI21_X1 U66499 ( .B1(n81294), .B2(n106122), .A(n81401), .ZN(n104050) );
  AOI22_X1 U66500 ( .A1(n73057), .A2(n106121), .B1(n81402), .B2(n106119), .ZN(
        n81401) );
  OAI21_X1 U66501 ( .B1(n106122), .B2(n81403), .A(n81404), .ZN(n104051) );
  AOI22_X1 U66502 ( .A1(n73341), .A2(n106121), .B1(n81405), .B2(n106118), .ZN(
        n81404) );
  OAI21_X1 U66503 ( .B1(n81278), .B2(n106122), .A(n81406), .ZN(n104052) );
  AOI22_X1 U66504 ( .A1(n71256), .A2(n106120), .B1(n106118), .B2(n81330), .ZN(
        n81406) );
  OAI21_X1 U66505 ( .B1(n81299), .B2(n106122), .A(n81407), .ZN(n104053) );
  AOI22_X1 U66506 ( .A1(n70221), .A2(n106120), .B1(n106119), .B2(n81377), .ZN(
        n81407) );
  OAI21_X1 U66507 ( .B1(n106123), .B2(n106099), .A(n81409), .ZN(n104054) );
  AOI22_X1 U66508 ( .A1(n70654), .A2(n106120), .B1(n81410), .B2(n106119), .ZN(
        n81409) );
  OAI21_X1 U66509 ( .B1(n81318), .B2(n106122), .A(n81411), .ZN(n104055) );
  AOI22_X1 U66510 ( .A1(n73637), .A2(n106120), .B1(n106118), .B2(n81320), .ZN(
        n81411) );
  OAI21_X1 U66511 ( .B1(n81383), .B2(n106122), .A(n81412), .ZN(n104056) );
  AOI22_X1 U66512 ( .A1(n73925), .A2(n106120), .B1(n106119), .B2(n81386), .ZN(
        n81412) );
  OAI21_X1 U66513 ( .B1(n106332), .B2(n106122), .A(n81413), .ZN(n104057) );
  AOI22_X1 U66514 ( .A1(n73784), .A2(n106120), .B1(n81414), .B2(n81391), .ZN(
        n81413) );
  OAI21_X1 U66515 ( .B1(n106122), .B2(n106096), .A(n81416), .ZN(n104058) );
  AOI22_X1 U66516 ( .A1(n71405), .A2(n106120), .B1(n81417), .B2(n106118), .ZN(
        n81416) );
  OAI21_X1 U66517 ( .B1(n105220), .B2(n106122), .A(n81418), .ZN(n104059) );
  AOI22_X1 U66518 ( .A1(n71556), .A2(n106120), .B1(n106119), .B2(n81335), .ZN(
        n81418) );
  OAI21_X1 U66519 ( .B1(n106259), .B2(n106091), .A(n81420), .ZN(n104060) );
  AOI22_X1 U66520 ( .A1(n106089), .A2(n109381), .B1(n106087), .B2(n81423), 
        .ZN(n81420) );
  OAI21_X1 U66521 ( .B1(n81349), .B2(n106092), .A(n81424), .ZN(n104061) );
  AOI22_X1 U66522 ( .A1(n81421), .A2(n109712), .B1(n81425), .B2(n81422), .ZN(
        n81424) );
  OAI21_X1 U66523 ( .B1(n106333), .B2(n106091), .A(n81426), .ZN(n104062) );
  AOI22_X1 U66524 ( .A1(n81421), .A2(n110498), .B1(n106087), .B2(n81414), .ZN(
        n81426) );
  OAI21_X1 U66525 ( .B1(n81306), .B2(n106092), .A(n81427), .ZN(n104063) );
  AOI22_X1 U66526 ( .A1(n74071), .A2(n106090), .B1(n81428), .B2(n81422), .ZN(
        n81427) );
  OAI21_X1 U66527 ( .B1(n81310), .B2(n106092), .A(n81429), .ZN(n104064) );
  AOI22_X1 U66528 ( .A1(n81421), .A2(n109606), .B1(n106087), .B2(n81313), .ZN(
        n81429) );
  OAI21_X1 U66529 ( .B1(n81284), .B2(n106091), .A(n81430), .ZN(n104065) );
  AOI22_X1 U66530 ( .A1(n81421), .A2(n108217), .B1(n106087), .B2(n81332), .ZN(
        n81430) );
  OAI21_X1 U66531 ( .B1(n106235), .B2(n106091), .A(n81431), .ZN(n104066) );
  AOI22_X1 U66532 ( .A1(n106089), .A2(n108451), .B1(n106087), .B2(n81322), 
        .ZN(n81431) );
  OAI21_X1 U66533 ( .B1(n106105), .B2(n106091), .A(n81432), .ZN(n104067) );
  AOI22_X1 U66534 ( .A1(n81421), .A2(n110175), .B1(n106087), .B2(n81405), .ZN(
        n81432) );
  OAI21_X1 U66535 ( .B1(n81318), .B2(n106091), .A(n81433), .ZN(n104068) );
  AOI22_X1 U66536 ( .A1(n106089), .A2(n110390), .B1(n106087), .B2(n81320), 
        .ZN(n81433) );
  OAI21_X1 U66537 ( .B1(n81340), .B2(n106091), .A(n81434), .ZN(n104069) );
  AOI22_X1 U66538 ( .A1(n106089), .A2(n108340), .B1(n106087), .B2(n81373), 
        .ZN(n81434) );
  OAI21_X1 U66539 ( .B1(n81383), .B2(n106091), .A(n81435), .ZN(n104070) );
  AOI22_X1 U66540 ( .A1(n106089), .A2(n110601), .B1(n106087), .B2(n81386), 
        .ZN(n81435) );
  OAI21_X1 U66541 ( .B1(n105220), .B2(n106091), .A(n81436), .ZN(n104071) );
  AOI22_X1 U66542 ( .A1(n106089), .A2(n108805), .B1(n106087), .B2(n81335), 
        .ZN(n81436) );
  OAI21_X1 U66543 ( .B1(n81278), .B2(n106091), .A(n81437), .ZN(n104072) );
  AOI22_X1 U66544 ( .A1(n106089), .A2(n108568), .B1(n106087), .B2(n81330), 
        .ZN(n81437) );
  OAI21_X1 U66545 ( .B1(n106094), .B2(n106091), .A(n81438), .ZN(n104073) );
  AOI22_X1 U66546 ( .A1(n106089), .A2(n108690), .B1(n106088), .B2(n81417), 
        .ZN(n81438) );
  OAI21_X1 U66547 ( .B1(n81284), .B2(n106086), .A(n81440), .ZN(n104074) );
  AOI22_X1 U66548 ( .A1(n106083), .A2(n81286), .B1(n106082), .B2(n108195), 
        .ZN(n81440) );
  OAI21_X1 U66549 ( .B1(n106262), .B2(n106078), .A(n81444), .ZN(n104075) );
  AOI22_X1 U66550 ( .A1(n106077), .A2(n109365), .B1(n106074), .B2(n81269), 
        .ZN(n81444) );
  OAI21_X1 U66551 ( .B1(n81278), .B2(n106079), .A(n81447), .ZN(n104076) );
  AOI22_X1 U66552 ( .A1(n106076), .A2(n108552), .B1(n106075), .B2(n106242), 
        .ZN(n81447) );
  OAI21_X1 U66553 ( .B1(n106254), .B2(n106078), .A(n81448), .ZN(n104077) );
  AOI22_X1 U66554 ( .A1(n106077), .A2(n110792), .B1(n106075), .B2(n81272), 
        .ZN(n81448) );
  OAI21_X1 U66555 ( .B1(n106203), .B2(n106079), .A(n81449), .ZN(n104078) );
  AOI22_X1 U66556 ( .A1(n106077), .A2(n110693), .B1(n106075), .B2(n81308), 
        .ZN(n81449) );
  OAI21_X1 U66557 ( .B1(n106146), .B2(n106078), .A(n81450), .ZN(n104079) );
  AOI22_X1 U66558 ( .A1(n106076), .A2(n107891), .B1(n106075), .B2(n81360), 
        .ZN(n81450) );
  OAI21_X1 U66559 ( .B1(n106079), .B2(n106072), .A(n81452), .ZN(n104080) );
  AOI22_X1 U66560 ( .A1(n106077), .A2(n107673), .B1(n81453), .B2(n81446), .ZN(
        n81452) );
  OAI21_X1 U66561 ( .B1(n106235), .B2(n106079), .A(n81454), .ZN(n104081) );
  AOI22_X1 U66562 ( .A1(n106076), .A2(n108435), .B1(n106075), .B2(n81283), 
        .ZN(n81454) );
  OAI21_X1 U66563 ( .B1(n81340), .B2(n106078), .A(n81455), .ZN(n104082) );
  AOI22_X1 U66564 ( .A1(n106076), .A2(n108324), .B1(n106075), .B2(n106169), 
        .ZN(n81455) );
  OAI21_X1 U66565 ( .B1(n81284), .B2(n106078), .A(n81456), .ZN(n104083) );
  AOI22_X1 U66566 ( .A1(n81445), .A2(n108201), .B1(n106075), .B2(n81286), .ZN(
        n81456) );
  OAI21_X1 U66567 ( .B1(n81345), .B2(n106078), .A(n81457), .ZN(n104084) );
  AOI22_X1 U66568 ( .A1(n81445), .A2(n110053), .B1(n106074), .B2(n81347), .ZN(
        n81457) );
  OAI21_X1 U66569 ( .B1(n105220), .B2(n106078), .A(n81458), .ZN(n104085) );
  AOI22_X1 U66570 ( .A1(n106076), .A2(n108789), .B1(n106074), .B2(n80188), 
        .ZN(n81458) );
  OAI21_X1 U66571 ( .B1(n81267), .B2(n106068), .A(n81460), .ZN(n104086) );
  AOI22_X1 U66572 ( .A1(n106066), .A2(n109368), .B1(n106063), .B2(n81269), 
        .ZN(n81460) );
  OAI21_X1 U66573 ( .B1(n81278), .B2(n106068), .A(n81463), .ZN(n104087) );
  AOI22_X1 U66574 ( .A1(n106065), .A2(n108555), .B1(n106064), .B2(n106241), 
        .ZN(n81463) );
  OAI21_X1 U66575 ( .B1(n106254), .B2(n106068), .A(n81464), .ZN(n104088) );
  AOI22_X1 U66576 ( .A1(n81461), .A2(n110795), .B1(n106064), .B2(n81272), .ZN(
        n81464) );
  OAI21_X1 U66577 ( .B1(n81306), .B2(n106068), .A(n81465), .ZN(n104089) );
  AOI22_X1 U66578 ( .A1(n81461), .A2(n110695), .B1(n106064), .B2(n81308), .ZN(
        n81465) );
  OAI21_X1 U66579 ( .B1(n106148), .B2(n106068), .A(n81466), .ZN(n104090) );
  AOI22_X1 U66580 ( .A1(n81461), .A2(n107893), .B1(n106064), .B2(n81360), .ZN(
        n81466) );
  OAI21_X1 U66581 ( .B1(n81451), .B2(n106068), .A(n81467), .ZN(n104091) );
  AOI22_X1 U66582 ( .A1(n81461), .A2(n107676), .B1(n106064), .B2(n81453), .ZN(
        n81467) );
  OAI21_X1 U66583 ( .B1(n106235), .B2(n106068), .A(n81468), .ZN(n104092) );
  AOI22_X1 U66584 ( .A1(n81461), .A2(n108438), .B1(n106064), .B2(n81283), .ZN(
        n81468) );
  OAI21_X1 U66585 ( .B1(n81284), .B2(n106068), .A(n81469), .ZN(n104093) );
  AOI22_X1 U66586 ( .A1(n81461), .A2(n108204), .B1(n106064), .B2(n81286), .ZN(
        n81469) );
  OAI21_X1 U66587 ( .B1(n81345), .B2(n106068), .A(n81470), .ZN(n104094) );
  AOI22_X1 U66588 ( .A1(n106066), .A2(n110056), .B1(n106063), .B2(n81347), 
        .ZN(n81470) );
  OAI21_X1 U66589 ( .B1(n81318), .B2(n106067), .A(n81471), .ZN(n104095) );
  AOI22_X1 U66590 ( .A1(n106066), .A2(n110380), .B1(n106062), .B2(n106064), 
        .ZN(n81471) );
  OAI21_X1 U66591 ( .B1(n81315), .B2(n106067), .A(n81473), .ZN(n104096) );
  AOI22_X1 U66592 ( .A1(n106066), .A2(n110271), .B1(n81474), .B2(n106064), 
        .ZN(n81473) );
  OAI21_X1 U66593 ( .B1(n105220), .B2(n106067), .A(n81475), .ZN(n104097) );
  AOI22_X1 U66594 ( .A1(n106066), .A2(n108792), .B1(n106063), .B2(n80188), 
        .ZN(n81475) );
  OAI21_X1 U66595 ( .B1(n106260), .B2(n106059), .A(n81477), .ZN(n104098) );
  AOI22_X1 U66596 ( .A1(n104766), .A2(n81269), .B1(n72276), .B2(n81479), .ZN(
        n81477) );
  OAI21_X1 U66597 ( .B1(n81340), .B2(n106059), .A(n81480), .ZN(n104099) );
  AOI22_X1 U66598 ( .A1(n104764), .A2(n106167), .B1(n70940), .B2(n104827), 
        .ZN(n81480) );
  OAI21_X1 U66599 ( .B1(n81340), .B2(n81439), .A(n81481), .ZN(n104100) );
  AOI22_X1 U66600 ( .A1(n106083), .A2(n106167), .B1(n106080), .B2(n108318), 
        .ZN(n81481) );
  OAI21_X1 U66601 ( .B1(n81278), .B2(n81439), .A(n81482), .ZN(n104101) );
  AOI22_X1 U66602 ( .A1(n106083), .A2(n106240), .B1(n106082), .B2(n108546), 
        .ZN(n81482) );
  OAI21_X1 U66603 ( .B1(n81315), .B2(n81439), .A(n81483), .ZN(n104102) );
  AOI22_X1 U66604 ( .A1(n81474), .A2(n106085), .B1(n106082), .B2(n110262), 
        .ZN(n81483) );
  OAI21_X1 U66605 ( .B1(n81318), .B2(n81439), .A(n81484), .ZN(n104103) );
  AOI22_X1 U66606 ( .A1(n106060), .A2(n106083), .B1(n106080), .B2(n110371), 
        .ZN(n81484) );
  OAI21_X1 U66607 ( .B1(n106246), .B2(n106059), .A(n81485), .ZN(n104104) );
  AOI22_X1 U66608 ( .A1(n104764), .A2(n106240), .B1(n71234), .B2(n104827), 
        .ZN(n81485) );
  OAI21_X1 U66609 ( .B1(n106149), .B2(n106059), .A(n81486), .ZN(n104105) );
  AOI22_X1 U66610 ( .A1(n104764), .A2(n81360), .B1(n70343), .B2(n104827), .ZN(
        n81486) );
  OAI21_X1 U66611 ( .B1(n106235), .B2(n106059), .A(n81487), .ZN(n104106) );
  AOI22_X1 U66612 ( .A1(n104765), .A2(n81283), .B1(n71085), .B2(n104828), .ZN(
        n81487) );
  OAI21_X1 U66613 ( .B1(n105220), .B2(n106059), .A(n81488), .ZN(n104107) );
  AOI22_X1 U66614 ( .A1(n104766), .A2(n80188), .B1(n71534), .B2(n104828), .ZN(
        n81488) );
  OAI21_X1 U66615 ( .B1(n106232), .B2(n106059), .A(n81489), .ZN(n104108) );
  AOI22_X1 U66616 ( .A1(n104764), .A2(n81286), .B1(n70781), .B2(n104827), .ZN(
        n81489) );
  OAI21_X1 U66617 ( .B1(n105220), .B2(n106086), .A(n81490), .ZN(n104109) );
  AOI22_X1 U66618 ( .A1(n106084), .A2(n80188), .B1(n106080), .B2(n108783), 
        .ZN(n81490) );
  OAI21_X1 U66619 ( .B1(n81267), .B2(n106086), .A(n81491), .ZN(n104110) );
  AOI22_X1 U66620 ( .A1(n106083), .A2(n81269), .B1(n106082), .B2(n109359), 
        .ZN(n81491) );
  OAI21_X1 U66621 ( .B1(n106236), .B2(n106086), .A(n81492), .ZN(n104111) );
  AOI22_X1 U66622 ( .A1(n106084), .A2(n81283), .B1(n106080), .B2(n108429), 
        .ZN(n81492) );
  OAI21_X1 U66623 ( .B1(n81284), .B2(n106058), .A(n81494), .ZN(n104112) );
  AOI22_X1 U66624 ( .A1(n81495), .A2(n108200), .B1(n104777), .B2(n81332), .ZN(
        n81494) );
  OAI21_X1 U66625 ( .B1(n106237), .B2(n106058), .A(n81497), .ZN(n104113) );
  AOI22_X1 U66626 ( .A1(n81495), .A2(n108434), .B1(n81496), .B2(n81322), .ZN(
        n81497) );
  OAI21_X1 U66627 ( .B1(n106058), .B2(n81498), .A(n81499), .ZN(n104114) );
  AOI22_X1 U66628 ( .A1(n81495), .A2(n108900), .B1(n81500), .B2(n81496), .ZN(
        n81499) );
  OAI21_X1 U66629 ( .B1(n81493), .B2(n106048), .A(n81502), .ZN(n104115) );
  AOI22_X1 U66630 ( .A1(n81495), .A2(n109138), .B1(n81503), .B2(n81496), .ZN(
        n81502) );
  OAI21_X1 U66631 ( .B1(n81267), .B2(n106058), .A(n81504), .ZN(n104116) );
  AOI22_X1 U66632 ( .A1(n81495), .A2(n109364), .B1(n81496), .B2(n81423), .ZN(
        n81504) );
  OAI21_X1 U66633 ( .B1(n106072), .B2(n81493), .A(n81505), .ZN(n104117) );
  AOI22_X1 U66634 ( .A1(n81495), .A2(n107672), .B1(n81506), .B2(n81496), .ZN(
        n81505) );
  OAI21_X1 U66635 ( .B1(n105220), .B2(n106058), .A(n81507), .ZN(n104118) );
  AOI22_X1 U66636 ( .A1(n81495), .A2(n108788), .B1(n81496), .B2(n81335), .ZN(
        n81507) );
  OAI21_X1 U66637 ( .B1(n81278), .B2(n106058), .A(n81508), .ZN(n104119) );
  AOI22_X1 U66638 ( .A1(n81495), .A2(n108551), .B1(n81496), .B2(n81330), .ZN(
        n81508) );
  OAI21_X1 U66639 ( .B1(n81493), .B2(n106046), .A(n81510), .ZN(n104120) );
  AOI22_X1 U66640 ( .A1(n81495), .A2(n109246), .B1(n81511), .B2(n104777), .ZN(
        n81510) );
  OAI21_X1 U66641 ( .B1(n81340), .B2(n106058), .A(n81512), .ZN(n104121) );
  AOI22_X1 U66642 ( .A1(n81495), .A2(n108323), .B1(n104777), .B2(n81373), .ZN(
        n81512) );
  OAI21_X1 U66643 ( .B1(n81501), .B2(n106041), .A(n81514), .ZN(n104122) );
  AOI22_X1 U66644 ( .A1(n104852), .A2(n81503), .B1(n106040), .B2(n109144), 
        .ZN(n81514) );
  OAI21_X1 U66645 ( .B1(n81498), .B2(n106042), .A(n81517), .ZN(n104123) );
  AOI22_X1 U66646 ( .A1(n104852), .A2(n81500), .B1(n106039), .B2(n108906), 
        .ZN(n81517) );
  OAI21_X1 U66647 ( .B1(n81267), .B2(n106041), .A(n81518), .ZN(n104124) );
  AOI22_X1 U66648 ( .A1(n104853), .A2(n81423), .B1(n106040), .B2(n109370), 
        .ZN(n81518) );
  OAI21_X1 U66649 ( .B1(n106243), .B2(n106042), .A(n81519), .ZN(n104125) );
  AOI22_X1 U66650 ( .A1(n81515), .A2(n81330), .B1(n106040), .B2(n108557), .ZN(
        n81519) );
  OAI21_X1 U66651 ( .B1(n106148), .B2(n106041), .A(n81520), .ZN(n104126) );
  AOI22_X1 U66652 ( .A1(n81521), .A2(n104852), .B1(n106039), .B2(n107895), 
        .ZN(n81520) );
  OAI21_X1 U66653 ( .B1(n106231), .B2(n106041), .A(n81522), .ZN(n104127) );
  AOI22_X1 U66654 ( .A1(n104853), .A2(n81332), .B1(n106039), .B2(n108206), 
        .ZN(n81522) );
  OAI21_X1 U66655 ( .B1(n106238), .B2(n106042), .A(n81523), .ZN(n104128) );
  AOI22_X1 U66656 ( .A1(n104852), .A2(n81322), .B1(n106040), .B2(n108440), 
        .ZN(n81523) );
  OAI21_X1 U66657 ( .B1(n81451), .B2(n106042), .A(n81524), .ZN(n104129) );
  AOI22_X1 U66658 ( .A1(n104852), .A2(n81506), .B1(n106040), .B2(n107678), 
        .ZN(n81524) );
  OAI21_X1 U66659 ( .B1(n105220), .B2(n106041), .A(n81525), .ZN(n104130) );
  AOI22_X1 U66660 ( .A1(n104853), .A2(n81335), .B1(n106040), .B2(n108794), 
        .ZN(n81525) );
  OAI21_X1 U66661 ( .B1(n81267), .B2(n106038), .A(n81527), .ZN(n104131) );
  AOI22_X1 U66662 ( .A1(n106036), .A2(n81269), .B1(n72264), .B2(n106034), .ZN(
        n81527) );
  OAI21_X1 U66663 ( .B1(n106243), .B2(n106037), .A(n81530), .ZN(n104132) );
  AOI22_X1 U66664 ( .A1(n106035), .A2(n106240), .B1(n71222), .B2(n106034), 
        .ZN(n81530) );
  OAI21_X1 U66665 ( .B1(n106235), .B2(n106037), .A(n81531), .ZN(n104133) );
  AOI22_X1 U66666 ( .A1(n106036), .A2(n81283), .B1(n71073), .B2(n106033), .ZN(
        n81531) );
  OAI21_X1 U66667 ( .B1(n81284), .B2(n106037), .A(n81532), .ZN(n104134) );
  AOI22_X1 U66668 ( .A1(n106035), .A2(n81286), .B1(n70769), .B2(n106034), .ZN(
        n81532) );
  OAI21_X1 U66669 ( .B1(n106165), .B2(n106037), .A(n81533), .ZN(n104135) );
  AOI22_X1 U66670 ( .A1(n106035), .A2(n81347), .B1(n73165), .B2(n106033), .ZN(
        n81533) );
  OAI21_X1 U66671 ( .B1(n81318), .B2(n106037), .A(n81534), .ZN(n104136) );
  AOI22_X1 U66672 ( .A1(n106035), .A2(n106060), .B1(n73603), .B2(n106034), 
        .ZN(n81534) );
  OAI21_X1 U66673 ( .B1(n81315), .B2(n106037), .A(n81535), .ZN(n104137) );
  AOI22_X1 U66674 ( .A1(n106036), .A2(n81474), .B1(n73454), .B2(n106033), .ZN(
        n81535) );
  OAI21_X1 U66675 ( .B1(n105220), .B2(n106037), .A(n81536), .ZN(n104138) );
  AOI22_X1 U66676 ( .A1(n106036), .A2(n80188), .B1(n71522), .B2(n106033), .ZN(
        n81536) );
  OAI21_X1 U66677 ( .B1(n81306), .B2(n106038), .A(n81537), .ZN(n104139) );
  AOI22_X1 U66678 ( .A1(n106035), .A2(n81308), .B1(n74033), .B2(n81529), .ZN(
        n81537) );
  OAI21_X1 U66679 ( .B1(n106137), .B2(n106037), .A(n81538), .ZN(n104140) );
  AOI22_X1 U66680 ( .A1(n81539), .A2(n81528), .B1(n69526), .B2(n106033), .ZN(
        n81538) );
  OAI21_X1 U66681 ( .B1(n81318), .B2(n106032), .A(n81541), .ZN(n104141) );
  AOI22_X1 U66682 ( .A1(n104876), .A2(n106060), .B1(n106031), .B2(n110367), 
        .ZN(n81541) );
  OAI21_X1 U66683 ( .B1(n105220), .B2(n106032), .A(n81544), .ZN(n104142) );
  AOI22_X1 U66684 ( .A1(n104875), .A2(n80188), .B1(n106031), .B2(n108779), 
        .ZN(n81544) );
  OAI21_X1 U66685 ( .B1(n106243), .B2(n81540), .A(n81545), .ZN(n104143) );
  AOI22_X1 U66686 ( .A1(n104875), .A2(n106240), .B1(n106031), .B2(n108542), 
        .ZN(n81545) );
  OAI21_X1 U66687 ( .B1(n106230), .B2(n106032), .A(n81546), .ZN(n104144) );
  AOI22_X1 U66688 ( .A1(n104876), .A2(n81286), .B1(n106031), .B2(n108191), 
        .ZN(n81546) );
  OAI21_X1 U66689 ( .B1(n106254), .B2(n106032), .A(n81547), .ZN(n104145) );
  AOI22_X1 U66690 ( .A1(n104877), .A2(n81272), .B1(n106031), .B2(n110782), 
        .ZN(n81547) );
  OAI21_X1 U66691 ( .B1(n106146), .B2(n106032), .A(n81548), .ZN(n104146) );
  AOI22_X1 U66692 ( .A1(n104876), .A2(n81360), .B1(n106031), .B2(n107882), 
        .ZN(n81548) );
  OAI21_X1 U66693 ( .B1(n106259), .B2(n106032), .A(n81549), .ZN(n104147) );
  AOI22_X1 U66694 ( .A1(n104876), .A2(n81269), .B1(n106031), .B2(n109355), 
        .ZN(n81549) );
  OAI21_X1 U66695 ( .B1(n106235), .B2(n106032), .A(n81550), .ZN(n104148) );
  AOI22_X1 U66696 ( .A1(n104875), .A2(n81283), .B1(n106031), .B2(n108425), 
        .ZN(n81550) );
  OAI21_X1 U66697 ( .B1(n81345), .B2(n106032), .A(n81551), .ZN(n104149) );
  AOI22_X1 U66698 ( .A1(n104877), .A2(n81347), .B1(n106030), .B2(n110043), 
        .ZN(n81551) );
  OAI21_X1 U66699 ( .B1(n81315), .B2(n106032), .A(n81552), .ZN(n104150) );
  AOI22_X1 U66700 ( .A1(n104877), .A2(n81474), .B1(n106030), .B2(n110259), 
        .ZN(n81552) );
  OAI21_X1 U66701 ( .B1(n81306), .B2(n106032), .A(n81553), .ZN(n104151) );
  AOI22_X1 U66702 ( .A1(n104877), .A2(n81308), .B1(n106030), .B2(n110684), 
        .ZN(n81553) );
  OAI21_X1 U66703 ( .B1(n106259), .B2(n106028), .A(n81555), .ZN(n104152) );
  AOI22_X1 U66704 ( .A1(n106027), .A2(n109348), .B1(n81557), .B2(n81269), .ZN(
        n81555) );
  OAI21_X1 U66705 ( .B1(n106243), .B2(n106028), .A(n81558), .ZN(n104153) );
  AOI22_X1 U66706 ( .A1(n106027), .A2(n108535), .B1(n104789), .B2(n106242), 
        .ZN(n81558) );
  OAI21_X1 U66707 ( .B1(n81299), .B2(n106028), .A(n81559), .ZN(n104154) );
  AOI22_X1 U66708 ( .A1(n106027), .A2(n107776), .B1(n104790), .B2(n81301), 
        .ZN(n81559) );
  OAI21_X1 U66709 ( .B1(n106235), .B2(n106028), .A(n81560), .ZN(n104155) );
  AOI22_X1 U66710 ( .A1(n106027), .A2(n108418), .B1(n104790), .B2(n81283), 
        .ZN(n81560) );
  OAI21_X1 U66711 ( .B1(n106233), .B2(n106028), .A(n81561), .ZN(n104156) );
  AOI22_X1 U66712 ( .A1(n106027), .A2(n108184), .B1(n104790), .B2(n81286), 
        .ZN(n81561) );
  OAI21_X1 U66713 ( .B1(n106163), .B2(n106028), .A(n81562), .ZN(n104157) );
  AOI22_X1 U66714 ( .A1(n106027), .A2(n110037), .B1(n104789), .B2(n81347), 
        .ZN(n81562) );
  OAI21_X1 U66715 ( .B1(n81318), .B2(n106028), .A(n81563), .ZN(n104158) );
  AOI22_X1 U66716 ( .A1(n106027), .A2(n110361), .B1(n104790), .B2(n106062), 
        .ZN(n81563) );
  OAI21_X1 U66717 ( .B1(n81394), .B2(n106025), .A(n81565), .ZN(n104159) );
  AOI22_X1 U66718 ( .A1(n106022), .A2(n109465), .B1(n106021), .B2(n106018), 
        .ZN(n81565) );
  OAI21_X1 U66719 ( .B1(n106243), .B2(n106025), .A(n81569), .ZN(n104160) );
  AOI22_X1 U66720 ( .A1(n106022), .A2(n108537), .B1(n106018), .B2(n106242), 
        .ZN(n81569) );
  OAI21_X1 U66721 ( .B1(n81299), .B2(n106025), .A(n81570), .ZN(n104161) );
  AOI22_X1 U66722 ( .A1(n106024), .A2(n107778), .B1(n106018), .B2(n81301), 
        .ZN(n81570) );
  OAI21_X1 U66723 ( .B1(n106231), .B2(n106025), .A(n81571), .ZN(n104162) );
  AOI22_X1 U66724 ( .A1(n106024), .A2(n108186), .B1(n106018), .B2(n81286), 
        .ZN(n81571) );
  OAI21_X1 U66725 ( .B1(n81345), .B2(n106025), .A(n81572), .ZN(n104163) );
  AOI22_X1 U66726 ( .A1(n106022), .A2(n110038), .B1(n106018), .B2(n81347), 
        .ZN(n81572) );
  OAI21_X1 U66727 ( .B1(n81318), .B2(n106025), .A(n81573), .ZN(n104164) );
  AOI22_X1 U66728 ( .A1(n106024), .A2(n110362), .B1(n106018), .B2(n106062), 
        .ZN(n81573) );
  OAI21_X1 U66729 ( .B1(n81315), .B2(n106025), .A(n81574), .ZN(n104165) );
  AOI22_X1 U66730 ( .A1(n106022), .A2(n110254), .B1(n106018), .B2(n81474), 
        .ZN(n81574) );
  OAI21_X1 U66731 ( .B1(n105220), .B2(n106025), .A(n81575), .ZN(n104166) );
  AOI22_X1 U66732 ( .A1(n106024), .A2(n108774), .B1(n106018), .B2(n80188), 
        .ZN(n81575) );
  OAI21_X1 U66733 ( .B1(n81349), .B2(n106025), .A(n81576), .ZN(n104167) );
  AOI22_X1 U66734 ( .A1(n106023), .A2(n109681), .B1(n106018), .B2(n81351), 
        .ZN(n81576) );
  OAI21_X1 U66735 ( .B1(n106254), .B2(n106025), .A(n81577), .ZN(n104168) );
  AOI22_X1 U66736 ( .A1(n106023), .A2(n110777), .B1(n106018), .B2(n81272), 
        .ZN(n81577) );
  OAI21_X1 U66737 ( .B1(n81306), .B2(n106025), .A(n81578), .ZN(n104169) );
  AOI22_X1 U66738 ( .A1(n106022), .A2(n110680), .B1(n106018), .B2(n81308), 
        .ZN(n81578) );
  OAI21_X1 U66739 ( .B1(n106149), .B2(n106025), .A(n81579), .ZN(n104170) );
  AOI22_X1 U66740 ( .A1(n106023), .A2(n107878), .B1(n106017), .B2(n81360), 
        .ZN(n81579) );
  OAI21_X1 U66741 ( .B1(n106054), .B2(n106015), .A(n81581), .ZN(n104171) );
  AOI22_X1 U66742 ( .A1(n104854), .A2(n81500), .B1(n71664), .B2(n106014), .ZN(
        n81581) );
  OAI21_X1 U66743 ( .B1(n106232), .B2(n106016), .A(n81584), .ZN(n104172) );
  AOI22_X1 U66744 ( .A1(n81582), .A2(n81332), .B1(n70767), .B2(n106013), .ZN(
        n81584) );
  OAI21_X1 U66745 ( .B1(n81501), .B2(n106015), .A(n81585), .ZN(n104173) );
  AOI22_X1 U66746 ( .A1(n104855), .A2(n81503), .B1(n71967), .B2(n106014), .ZN(
        n81585) );
  OAI21_X1 U66747 ( .B1(n81340), .B2(n106016), .A(n81586), .ZN(n104174) );
  AOI22_X1 U66748 ( .A1(n104854), .A2(n81373), .B1(n70926), .B2(n106013), .ZN(
        n81586) );
  OAI21_X1 U66749 ( .B1(n106243), .B2(n106015), .A(n81587), .ZN(n104175) );
  AOI22_X1 U66750 ( .A1(n104854), .A2(n81330), .B1(n71220), .B2(n106014), .ZN(
        n81587) );
  OAI21_X1 U66751 ( .B1(n106010), .B2(n106016), .A(n81589), .ZN(n104176) );
  AOI22_X1 U66752 ( .A1(n81590), .A2(n104854), .B1(n71813), .B2(n106014), .ZN(
        n81589) );
  OAI21_X1 U66753 ( .B1(n81394), .B2(n106016), .A(n81591), .ZN(n104177) );
  AOI22_X1 U66754 ( .A1(n104855), .A2(n81396), .B1(n72413), .B2(n106014), .ZN(
        n81591) );
  OAI21_X1 U66755 ( .B1(n106095), .B2(n106016), .A(n81592), .ZN(n104178) );
  AOI22_X1 U66756 ( .A1(n81582), .A2(n81417), .B1(n71369), .B2(n81583), .ZN(
        n81592) );
  OAI21_X1 U66757 ( .B1(n105218), .B2(n106015), .A(n81593), .ZN(n104179) );
  AOI22_X1 U66758 ( .A1(n104854), .A2(n81335), .B1(n71520), .B2(n106013), .ZN(
        n81593) );
  OAI21_X1 U66759 ( .B1(n81394), .B2(n106006), .A(n81595), .ZN(n104180) );
  AOI22_X1 U66760 ( .A1(n106003), .A2(n81396), .B1(n104941), .B2(n109464), 
        .ZN(n81595) );
  OAI21_X1 U66761 ( .B1(n81284), .B2(n81594), .A(n81598), .ZN(n104181) );
  AOI22_X1 U66762 ( .A1(n106005), .A2(n81332), .B1(n104942), .B2(n108185), 
        .ZN(n81598) );
  OAI21_X1 U66763 ( .B1(n106237), .B2(n81594), .A(n81599), .ZN(n104182) );
  AOI22_X1 U66764 ( .A1(n106004), .A2(n81322), .B1(n104942), .B2(n108419), 
        .ZN(n81599) );
  OAI21_X1 U66765 ( .B1(n106160), .B2(n81594), .A(n81600), .ZN(n104183) );
  AOI22_X1 U66766 ( .A1(n106005), .A2(n81425), .B1(n104943), .B2(n109680), 
        .ZN(n81600) );
  OAI21_X1 U66767 ( .B1(n81340), .B2(n106006), .A(n81601), .ZN(n104184) );
  AOI22_X1 U66768 ( .A1(n106004), .A2(n81373), .B1(n104941), .B2(n108308), 
        .ZN(n81601) );
  OAI21_X1 U66769 ( .B1(n106243), .B2(n81594), .A(n81602), .ZN(n104185) );
  AOI22_X1 U66770 ( .A1(n106005), .A2(n81330), .B1(n104944), .B2(n108536), 
        .ZN(n81602) );
  OAI21_X1 U66771 ( .B1(n106162), .B2(n81594), .A(n81603), .ZN(n104186) );
  AOI22_X1 U66772 ( .A1(n81604), .A2(n106003), .B1(n73159), .B2(n104941), .ZN(
        n81603) );
  OAI21_X1 U66773 ( .B1(n105219), .B2(n106006), .A(n81605), .ZN(n104187) );
  AOI22_X1 U66774 ( .A1(n106004), .A2(n81335), .B1(n104945), .B2(n108773), 
        .ZN(n81605) );
  OAI21_X1 U66775 ( .B1(n81299), .B2(n81594), .A(n81606), .ZN(n104188) );
  AOI22_X1 U66776 ( .A1(n106004), .A2(n81377), .B1(n104941), .B2(n107777), 
        .ZN(n81606) );
  OAI21_X1 U66777 ( .B1(n106094), .B2(n81594), .A(n81607), .ZN(n104189) );
  AOI22_X1 U66778 ( .A1(n106005), .A2(n81417), .B1(n104946), .B2(n108658), 
        .ZN(n81607) );
  OAI21_X1 U66779 ( .B1(n106147), .B2(n106002), .A(n81609), .ZN(n104190) );
  AOI22_X1 U66780 ( .A1(n104850), .A2(n81521), .B1(n104865), .B2(n107884), 
        .ZN(n81609) );
  OAI21_X1 U66781 ( .B1(n105218), .B2(n106002), .A(n81612), .ZN(n104191) );
  AOI22_X1 U66782 ( .A1(n104851), .A2(n81335), .B1(n104866), .B2(n108781), 
        .ZN(n81612) );
  OAI21_X1 U66783 ( .B1(n106232), .B2(n106002), .A(n81613), .ZN(n104192) );
  AOI22_X1 U66784 ( .A1(n104849), .A2(n81332), .B1(n104867), .B2(n108193), 
        .ZN(n81613) );
  OAI21_X1 U66785 ( .B1(n106096), .B2(n106002), .A(n81614), .ZN(n104193) );
  AOI22_X1 U66786 ( .A1(n104851), .A2(n81417), .B1(n104866), .B2(n108666), 
        .ZN(n81614) );
  OAI21_X1 U66787 ( .B1(n81501), .B2(n106002), .A(n81615), .ZN(n104194) );
  AOI22_X1 U66788 ( .A1(n104850), .A2(n81503), .B1(n104867), .B2(n109131), 
        .ZN(n81615) );
  OAI21_X1 U66789 ( .B1(n106259), .B2(n106002), .A(n81616), .ZN(n104195) );
  AOI22_X1 U66790 ( .A1(n104849), .A2(n81423), .B1(n104865), .B2(n109357), 
        .ZN(n81616) );
  OAI21_X1 U66791 ( .B1(n106243), .B2(n106002), .A(n81617), .ZN(n104196) );
  AOI22_X1 U66792 ( .A1(n104850), .A2(n81330), .B1(n104865), .B2(n108544), 
        .ZN(n81617) );
  OAI21_X1 U66793 ( .B1(n106237), .B2(n106002), .A(n81618), .ZN(n104197) );
  AOI22_X1 U66794 ( .A1(n104849), .A2(n81322), .B1(n104866), .B2(n108427), 
        .ZN(n81618) );
  OAI21_X1 U66795 ( .B1(n81284), .B2(n106001), .A(n81620), .ZN(n104198) );
  AOI22_X1 U66796 ( .A1(n106000), .A2(n108177), .B1(n105996), .B2(n81332), 
        .ZN(n81620) );
  OAI21_X1 U66797 ( .B1(n106158), .B2(n81619), .A(n81623), .ZN(n104199) );
  AOI22_X1 U66798 ( .A1(n105999), .A2(n109672), .B1(n105996), .B2(n81425), 
        .ZN(n81623) );
  OAI21_X1 U66799 ( .B1(n81340), .B2(n106001), .A(n81624), .ZN(n104200) );
  AOI22_X1 U66800 ( .A1(n106000), .A2(n108300), .B1(n105996), .B2(n81373), 
        .ZN(n81624) );
  OAI21_X1 U66801 ( .B1(n106163), .B2(n81619), .A(n81625), .ZN(n104201) );
  AOI22_X1 U66802 ( .A1(n105999), .A2(n110030), .B1(n105997), .B2(n81604), 
        .ZN(n81625) );
  OAI21_X1 U66803 ( .B1(n106105), .B2(n81619), .A(n81626), .ZN(n104202) );
  AOI22_X1 U66804 ( .A1(n106000), .A2(n110137), .B1(n105997), .B2(n81405), 
        .ZN(n81626) );
  OAI21_X1 U66805 ( .B1(n106243), .B2(n106001), .A(n81627), .ZN(n104203) );
  AOI22_X1 U66806 ( .A1(n106000), .A2(n108528), .B1(n105997), .B2(n81330), 
        .ZN(n81627) );
  OAI21_X1 U66807 ( .B1(n81628), .B2(n105992), .A(n81630), .ZN(n104204) );
  AOI22_X1 U66808 ( .A1(n105987), .A2(n81632), .B1(n105985), .B2(n110874), 
        .ZN(n81630) );
  OAI21_X1 U66809 ( .B1(n81498), .B2(n105983), .A(n81635), .ZN(n104205) );
  AOI22_X1 U66810 ( .A1(n105980), .A2(n108879), .B1(n105979), .B2(n81500), 
        .ZN(n81635) );
  OAI21_X1 U66811 ( .B1(n81378), .B2(n105983), .A(n81638), .ZN(n104206) );
  AOI22_X1 U66812 ( .A1(n105981), .A2(n107233), .B1(n105979), .B2(n81380), 
        .ZN(n81638) );
  OAI21_X1 U66813 ( .B1(n106172), .B2(n81634), .A(n81639), .ZN(n104207) );
  AOI22_X1 U66814 ( .A1(n105982), .A2(n108302), .B1(n105978), .B2(n81373), 
        .ZN(n81639) );
  OAI21_X1 U66815 ( .B1(n81284), .B2(n105983), .A(n81640), .ZN(n104208) );
  AOI22_X1 U66816 ( .A1(n105981), .A2(n108179), .B1(n105979), .B2(n81332), 
        .ZN(n81640) );
  OAI21_X1 U66817 ( .B1(n106236), .B2(n81634), .A(n81641), .ZN(n104209) );
  AOI22_X1 U66818 ( .A1(n105982), .A2(n108413), .B1(n105978), .B2(n81322), 
        .ZN(n81641) );
  OAI21_X1 U66819 ( .B1(n81299), .B2(n105983), .A(n81642), .ZN(n104210) );
  AOI22_X1 U66820 ( .A1(n105981), .A2(n107771), .B1(n105979), .B2(n81377), 
        .ZN(n81642) );
  OAI21_X1 U66821 ( .B1(n106243), .B2(n81634), .A(n81643), .ZN(n104211) );
  AOI22_X1 U66822 ( .A1(n105982), .A2(n108530), .B1(n105978), .B2(n81330), 
        .ZN(n81643) );
  OAI21_X1 U66823 ( .B1(n106093), .B2(n81634), .A(n81644), .ZN(n104212) );
  AOI22_X1 U66824 ( .A1(n105981), .A2(n108652), .B1(n105978), .B2(n81417), 
        .ZN(n81644) );
  OAI21_X1 U66825 ( .B1(n106149), .B2(n81634), .A(n81645), .ZN(n104213) );
  AOI22_X1 U66826 ( .A1(n70317), .A2(n105980), .B1(n105977), .B2(n81521), .ZN(
        n81645) );
  OAI21_X1 U66827 ( .B1(n105220), .B2(n81634), .A(n81646), .ZN(n104214) );
  AOI22_X1 U66828 ( .A1(n105982), .A2(n108767), .B1(n105979), .B2(n81335), 
        .ZN(n81646) );
  OAI21_X1 U66829 ( .B1(n106243), .B2(n105976), .A(n81648), .ZN(n104215) );
  AOI22_X1 U66830 ( .A1(n104929), .A2(n108512), .B1(n105975), .B2(n81330), 
        .ZN(n81648) );
  OAI21_X1 U66831 ( .B1(n81647), .B2(n81651), .A(n81652), .ZN(n104216) );
  AOI22_X1 U66832 ( .A1(n104930), .A2(n107953), .B1(n81653), .B2(n105973), 
        .ZN(n81652) );
  OAI21_X1 U66833 ( .B1(n81284), .B2(n105976), .A(n81654), .ZN(n104217) );
  AOI22_X1 U66834 ( .A1(n104931), .A2(n108161), .B1(n105974), .B2(n81332), 
        .ZN(n81654) );
  OAI21_X1 U66835 ( .B1(n105218), .B2(n81647), .A(n81655), .ZN(n104218) );
  AOI22_X1 U66836 ( .A1(n104930), .A2(n108749), .B1(n105974), .B2(n81335), 
        .ZN(n81655) );
  OAI21_X1 U66837 ( .B1(n106095), .B2(n81647), .A(n81656), .ZN(n104219) );
  AOI22_X1 U66838 ( .A1(n104929), .A2(n108634), .B1(n105974), .B2(n81417), 
        .ZN(n81656) );
  OAI21_X1 U66839 ( .B1(n81498), .B2(n81647), .A(n81657), .ZN(n104220) );
  AOI22_X1 U66840 ( .A1(n104929), .A2(n108861), .B1(n105975), .B2(n81500), 
        .ZN(n81657) );
  OAI21_X1 U66841 ( .B1(n106055), .B2(n105966), .A(n81659), .ZN(n104221) );
  AOI22_X1 U66842 ( .A1(n81660), .A2(n81500), .B1(n71632), .B2(n104990), .ZN(
        n81659) );
  OAI21_X1 U66843 ( .B1(n106231), .B2(n105967), .A(n81662), .ZN(n104222) );
  AOI22_X1 U66844 ( .A1(n105964), .A2(n81332), .B1(n70735), .B2(n104991), .ZN(
        n81662) );
  OAI21_X1 U66845 ( .B1(n106147), .B2(n105967), .A(n81663), .ZN(n104223) );
  AOI22_X1 U66846 ( .A1(n81660), .A2(n81521), .B1(n70297), .B2(n104990), .ZN(
        n81663) );
  OAI21_X1 U66847 ( .B1(n105971), .B2(n105967), .A(n81664), .ZN(n104224) );
  AOI22_X1 U66848 ( .A1(n105964), .A2(n81653), .B1(n70439), .B2(n81661), .ZN(
        n81664) );
  OAI21_X1 U66849 ( .B1(n106137), .B2(n105966), .A(n81665), .ZN(n104225) );
  AOI22_X1 U66850 ( .A1(n105964), .A2(n81380), .B1(n69492), .B2(n81661), .ZN(
        n81665) );
  OAI21_X1 U66851 ( .B1(n107369), .B2(n105961), .A(n81667), .ZN(n104226) );
  AOI22_X1 U66852 ( .A1(n105959), .A2(n81396), .B1(n105957), .B2(n109522), 
        .ZN(n81667) );
  OAI21_X1 U66853 ( .B1(n107412), .B2(n105962), .A(n81670), .ZN(n104227) );
  AOI22_X1 U66854 ( .A1(n105958), .A2(n81330), .B1(n105957), .B2(n108592), 
        .ZN(n81670) );
  OAI21_X1 U66855 ( .B1(n107408), .B2(n105961), .A(n81671), .ZN(n104228) );
  AOI22_X1 U66856 ( .A1(n105958), .A2(n81506), .B1(n105957), .B2(n107715), 
        .ZN(n81671) );
  OAI21_X1 U66857 ( .B1(n107406), .B2(n105961), .A(n81672), .ZN(n104229) );
  AOI22_X1 U66858 ( .A1(n105958), .A2(n81322), .B1(n105957), .B2(n108478), 
        .ZN(n81672) );
  OAI21_X1 U66859 ( .B1(n107404), .B2(n105962), .A(n81673), .ZN(n104230) );
  AOI22_X1 U66860 ( .A1(n105958), .A2(n81373), .B1(n105957), .B2(n108367), 
        .ZN(n81673) );
  OAI21_X1 U66861 ( .B1(n107402), .B2(n105961), .A(n81674), .ZN(n104231) );
  AOI22_X1 U66862 ( .A1(n105958), .A2(n81332), .B1(n105957), .B2(n108244), 
        .ZN(n81674) );
  OAI21_X1 U66863 ( .B1(n111057), .B2(n105962), .A(n81675), .ZN(n104232) );
  AOI22_X1 U66864 ( .A1(n105958), .A2(n81327), .B1(n105957), .B2(n107205), 
        .ZN(n81675) );
  OAI21_X1 U66865 ( .B1(n111058), .B2(n105962), .A(n81676), .ZN(n104233) );
  AOI22_X1 U66866 ( .A1(n105958), .A2(n81335), .B1(n105957), .B2(n108831), 
        .ZN(n81676) );
  OAI21_X1 U66867 ( .B1(n111059), .B2(n105962), .A(n81677), .ZN(n104234) );
  AOI22_X1 U66868 ( .A1(n105958), .A2(n81500), .B1(n105956), .B2(n108943), 
        .ZN(n81677) );
  OAI21_X1 U66869 ( .B1(n111060), .B2(n105962), .A(n81678), .ZN(n104235) );
  AOI22_X1 U66870 ( .A1(n105958), .A2(n81417), .B1(n105956), .B2(n108715), 
        .ZN(n81678) );
  OAI21_X1 U66871 ( .B1(n111062), .B2(n105962), .A(n81679), .ZN(n104236) );
  AOI22_X1 U66872 ( .A1(n105958), .A2(n81511), .B1(n105956), .B2(n109288), 
        .ZN(n81679) );
  OAI21_X1 U66873 ( .B1(n107412), .B2(n105953), .A(n81681), .ZN(n104237) );
  AOI22_X1 U66874 ( .A1(n104688), .A2(n108596), .B1(n104962), .B2(n81330), 
        .ZN(n81681) );
  OAI21_X1 U66875 ( .B1(n107408), .B2(n105952), .A(n81684), .ZN(n104238) );
  AOI22_X1 U66876 ( .A1(n81682), .A2(n107719), .B1(n104964), .B2(n81506), .ZN(
        n81684) );
  OAI21_X1 U66877 ( .B1(n107406), .B2(n105952), .A(n81685), .ZN(n104239) );
  AOI22_X1 U66878 ( .A1(n81682), .A2(n108482), .B1(n104964), .B2(n81322), .ZN(
        n81685) );
  OAI21_X1 U66879 ( .B1(n107404), .B2(n105953), .A(n81686), .ZN(n104240) );
  AOI22_X1 U66880 ( .A1(n104689), .A2(n108371), .B1(n104962), .B2(n81373), 
        .ZN(n81686) );
  OAI21_X1 U66881 ( .B1(n107402), .B2(n105952), .A(n81687), .ZN(n104241) );
  AOI22_X1 U66882 ( .A1(n81682), .A2(n108248), .B1(n104963), .B2(n81332), .ZN(
        n81687) );
  OAI21_X1 U66883 ( .B1(n107376), .B2(n105950), .A(n81689), .ZN(n104242) );
  AOI22_X1 U66884 ( .A1(n70260), .A2(n105946), .B1(n104955), .B2(n81377), .ZN(
        n81689) );
  OAI21_X1 U66885 ( .B1(n107371), .B2(n105949), .A(n81692), .ZN(n104243) );
  AOI22_X1 U66886 ( .A1(n70404), .A2(n105946), .B1(n104954), .B2(n81521), .ZN(
        n81692) );
  OAI21_X1 U66887 ( .B1(n106832), .B2(n105950), .A(n81693), .ZN(n104244) );
  AOI22_X1 U66888 ( .A1(n69465), .A2(n105947), .B1(n104953), .B2(n81380), .ZN(
        n81693) );
  OAI21_X1 U66889 ( .B1(n107380), .B2(n105949), .A(n81694), .ZN(n104245) );
  AOI22_X1 U66890 ( .A1(n70693), .A2(n105947), .B1(n104953), .B2(n81410), .ZN(
        n81694) );
  OAI21_X1 U66891 ( .B1(n107388), .B2(n105949), .A(n81695), .ZN(n104246) );
  AOI22_X1 U66892 ( .A1(n73527), .A2(n105946), .B1(n104953), .B2(n81317), .ZN(
        n81695) );
  OAI21_X1 U66893 ( .B1(n107394), .B2(n105950), .A(n81696), .ZN(n104247) );
  AOI22_X1 U66894 ( .A1(n73238), .A2(n105947), .B1(n104954), .B2(n81604), .ZN(
        n81696) );
  OAI21_X1 U66895 ( .B1(n107392), .B2(n105949), .A(n81697), .ZN(n104248) );
  AOI22_X1 U66896 ( .A1(n73676), .A2(n105946), .B1(n104955), .B2(n81320), .ZN(
        n81697) );
  OAI21_X1 U66897 ( .B1(n107378), .B2(n105950), .A(n81698), .ZN(n104249) );
  AOI22_X1 U66898 ( .A1(n74106), .A2(n105947), .B1(n104955), .B2(n81428), .ZN(
        n81698) );
  OAI21_X1 U66899 ( .B1(n107382), .B2(n105950), .A(n81699), .ZN(n104250) );
  AOI22_X1 U66900 ( .A1(n74247), .A2(n105948), .B1(n81700), .B2(n104955), .ZN(
        n81699) );
  OAI21_X1 U66901 ( .B1(n107373), .B2(n105950), .A(n81701), .ZN(n104251) );
  AOI22_X1 U66902 ( .A1(n70546), .A2(n105948), .B1(n104954), .B2(n81653), .ZN(
        n81701) );
  OAI21_X1 U66903 ( .B1(n107396), .B2(n105950), .A(n81702), .ZN(n104252) );
  AOI22_X1 U66904 ( .A1(n73380), .A2(n105948), .B1(n104954), .B2(n81405), .ZN(
        n81702) );
  OAI21_X1 U66905 ( .B1(n111060), .B2(n105944), .A(n81704), .ZN(n104253) );
  AOI22_X1 U66906 ( .A1(n105942), .A2(n81417), .B1(n105939), .B2(n108711), 
        .ZN(n81704) );
  OAI21_X1 U66907 ( .B1(n111059), .B2(n105943), .A(n81707), .ZN(n104254) );
  AOI22_X1 U66908 ( .A1(n105942), .A2(n81500), .B1(n105939), .B2(n108939), 
        .ZN(n81707) );
  OAI21_X1 U66909 ( .B1(n108974), .B2(n105943), .A(n81708), .ZN(n104255) );
  AOI22_X1 U66910 ( .A1(n105942), .A2(n81590), .B1(n105939), .B2(n109056), 
        .ZN(n81708) );
  OAI21_X1 U66911 ( .B1(n111058), .B2(n105944), .A(n81709), .ZN(n104256) );
  AOI22_X1 U66912 ( .A1(n105942), .A2(n81335), .B1(n105939), .B2(n108827), 
        .ZN(n81709) );
  OAI21_X1 U66913 ( .B1(n111061), .B2(n105944), .A(n81710), .ZN(n104257) );
  AOI22_X1 U66914 ( .A1(n105942), .A2(n81503), .B1(n105939), .B2(n109176), 
        .ZN(n81710) );
  OAI21_X1 U66915 ( .B1(n111062), .B2(n105943), .A(n81711), .ZN(n104258) );
  AOI22_X1 U66916 ( .A1(n105942), .A2(n81511), .B1(n105939), .B2(n109284), 
        .ZN(n81711) );
  OAI21_X1 U66917 ( .B1(n111057), .B2(n105944), .A(n81712), .ZN(n104259) );
  AOI22_X1 U66918 ( .A1(n105942), .A2(n81327), .B1(n105939), .B2(n107213), 
        .ZN(n81712) );
  OAI21_X1 U66919 ( .B1(n111063), .B2(n105943), .A(n81713), .ZN(n104260) );
  AOI22_X1 U66920 ( .A1(n105942), .A2(n81423), .B1(n105939), .B2(n109403), 
        .ZN(n81713) );
  OAI21_X1 U66921 ( .B1(n107371), .B2(n105944), .A(n81714), .ZN(n104261) );
  AOI22_X1 U66922 ( .A1(n105941), .A2(n81521), .B1(n105938), .B2(n107922), 
        .ZN(n81714) );
  OAI21_X1 U66923 ( .B1(n107380), .B2(n105944), .A(n81715), .ZN(n104262) );
  AOI22_X1 U66924 ( .A1(n105941), .A2(n81410), .B1(n105938), .B2(n108126), 
        .ZN(n81715) );
  OAI21_X1 U66925 ( .B1(n107373), .B2(n105944), .A(n81716), .ZN(n104263) );
  AOI22_X1 U66926 ( .A1(n105941), .A2(n81653), .B1(n105938), .B2(n108018), 
        .ZN(n81716) );
  OAI21_X1 U66927 ( .B1(n107376), .B2(n105944), .A(n81717), .ZN(n104264) );
  AOI22_X1 U66928 ( .A1(n105941), .A2(n81377), .B1(n105938), .B2(n107826), 
        .ZN(n81717) );
  OAI21_X1 U66929 ( .B1(n106832), .B2(n105944), .A(n81718), .ZN(n104265) );
  AOI22_X1 U66930 ( .A1(n105941), .A2(n81380), .B1(n105938), .B2(n107212), 
        .ZN(n81718) );
  OAI21_X1 U66931 ( .B1(n107384), .B2(n105944), .A(n81719), .ZN(n104266) );
  AOI22_X1 U66932 ( .A1(n105941), .A2(n81632), .B1(n105938), .B2(n110926), 
        .ZN(n81719) );
  OAI21_X1 U66933 ( .B1(n107388), .B2(n105944), .A(n81720), .ZN(n104267) );
  AOI22_X1 U66934 ( .A1(n105941), .A2(n81317), .B1(n105938), .B2(n110304), 
        .ZN(n81720) );
  OAI21_X1 U66935 ( .B1(n107412), .B2(n105944), .A(n81721), .ZN(n104268) );
  AOI22_X1 U66936 ( .A1(n105941), .A2(n81330), .B1(n105938), .B2(n108588), 
        .ZN(n81721) );
  OAI21_X1 U66937 ( .B1(n107404), .B2(n105944), .A(n81722), .ZN(n104269) );
  AOI22_X1 U66938 ( .A1(n105941), .A2(n81373), .B1(n105938), .B2(n108363), 
        .ZN(n81722) );
  OAI21_X1 U66939 ( .B1(n107408), .B2(n105944), .A(n81723), .ZN(n104270) );
  AOI22_X1 U66940 ( .A1(n105941), .A2(n81506), .B1(n105938), .B2(n107711), 
        .ZN(n81723) );
  OAI21_X1 U66941 ( .B1(n107367), .B2(n105944), .A(n81724), .ZN(n104271) );
  AOI22_X1 U66942 ( .A1(n105941), .A2(n81425), .B1(n105938), .B2(n109733), 
        .ZN(n81724) );
  OAI21_X1 U66943 ( .B1(n107394), .B2(n105944), .A(n81725), .ZN(n104272) );
  AOI22_X1 U66944 ( .A1(n105941), .A2(n81604), .B1(n105938), .B2(n110091), 
        .ZN(n81725) );
  OAI21_X1 U66945 ( .B1(n107369), .B2(n105943), .A(n81726), .ZN(n104273) );
  AOI22_X1 U66946 ( .A1(n105940), .A2(n81396), .B1(n105937), .B2(n109518), 
        .ZN(n81726) );
  OAI21_X1 U66947 ( .B1(n107400), .B2(n105943), .A(n81727), .ZN(n104274) );
  AOI22_X1 U66948 ( .A1(n105940), .A2(n81400), .B1(n105937), .B2(n109866), 
        .ZN(n81727) );
  OAI21_X1 U66949 ( .B1(n107406), .B2(n105943), .A(n81728), .ZN(n104275) );
  AOI22_X1 U66950 ( .A1(n105940), .A2(n81322), .B1(n105937), .B2(n108474), 
        .ZN(n81728) );
  OAI21_X1 U66951 ( .B1(n107410), .B2(n105943), .A(n81729), .ZN(n104276) );
  AOI22_X1 U66952 ( .A1(n105940), .A2(n81313), .B1(n105937), .B2(n109626), 
        .ZN(n81729) );
  OAI21_X1 U66953 ( .B1(n107402), .B2(n105943), .A(n81730), .ZN(n104277) );
  AOI22_X1 U66954 ( .A1(n105940), .A2(n81332), .B1(n105937), .B2(n108240), 
        .ZN(n81730) );
  OAI21_X1 U66955 ( .B1(n107396), .B2(n105943), .A(n81731), .ZN(n104278) );
  AOI22_X1 U66956 ( .A1(n105940), .A2(n81405), .B1(n105937), .B2(n110198), 
        .ZN(n81731) );
  OAI21_X1 U66957 ( .B1(n107398), .B2(n105943), .A(n81732), .ZN(n104279) );
  AOI22_X1 U66958 ( .A1(n105940), .A2(n81402), .B1(n105937), .B2(n109983), 
        .ZN(n81732) );
  OAI21_X1 U66959 ( .B1(n105219), .B2(n105936), .A(n81734), .ZN(n104280) );
  AOI22_X1 U66960 ( .A1(n105935), .A2(n108766), .B1(n105932), .B2(n80188), 
        .ZN(n81734) );
  OAI21_X1 U66961 ( .B1(n106243), .B2(n105936), .A(n81737), .ZN(n104281) );
  AOI22_X1 U66962 ( .A1(n105933), .A2(n108529), .B1(n105930), .B2(n106242), 
        .ZN(n81737) );
  OAI21_X1 U66963 ( .B1(n81299), .B2(n105936), .A(n81738), .ZN(n104282) );
  AOI22_X1 U66964 ( .A1(n105935), .A2(n107770), .B1(n105932), .B2(n81301), 
        .ZN(n81738) );
  OAI21_X1 U66965 ( .B1(n106138), .B2(n105936), .A(n81739), .ZN(n104283) );
  AOI22_X1 U66966 ( .A1(n105933), .A2(n107232), .B1(n105930), .B2(n81539), 
        .ZN(n81739) );
  OAI21_X1 U66967 ( .B1(n106259), .B2(n105936), .A(n81740), .ZN(n104284) );
  AOI22_X1 U66968 ( .A1(n105935), .A2(n109342), .B1(n105932), .B2(n81269), 
        .ZN(n81740) );
  OAI21_X1 U66969 ( .B1(n106116), .B2(n105936), .A(n81741), .ZN(n104285) );
  AOI22_X1 U66970 ( .A1(n105933), .A2(n109457), .B1(n105930), .B2(n106020), 
        .ZN(n81741) );
  OAI21_X1 U66971 ( .B1(n106238), .B2(n105936), .A(n81742), .ZN(n104286) );
  AOI22_X1 U66972 ( .A1(n105935), .A2(n108412), .B1(n105932), .B2(n81283), 
        .ZN(n81742) );
  OAI21_X1 U66973 ( .B1(n106230), .B2(n105936), .A(n81743), .ZN(n104287) );
  AOI22_X1 U66974 ( .A1(n105933), .A2(n108178), .B1(n105930), .B2(n81286), 
        .ZN(n81743) );
  OAI21_X1 U66975 ( .B1(n106148), .B2(n105936), .A(n81744), .ZN(n104288) );
  AOI22_X1 U66976 ( .A1(n105935), .A2(n107872), .B1(n105932), .B2(n81360), 
        .ZN(n81744) );
  OAI21_X1 U66977 ( .B1(n105220), .B2(n105929), .A(n81746), .ZN(n104289) );
  AOI22_X1 U66978 ( .A1(n105926), .A2(n108769), .B1(n105925), .B2(n80188), 
        .ZN(n81746) );
  OAI21_X1 U66979 ( .B1(n106259), .B2(n105929), .A(n81749), .ZN(n104290) );
  AOI22_X1 U66980 ( .A1(n105926), .A2(n109345), .B1(n105923), .B2(n81269), 
        .ZN(n81749) );
  OAI21_X1 U66981 ( .B1(n106113), .B2(n105929), .A(n81750), .ZN(n104291) );
  AOI22_X1 U66982 ( .A1(n105928), .A2(n109460), .B1(n105923), .B2(n106020), 
        .ZN(n81750) );
  OAI21_X1 U66983 ( .B1(n81278), .B2(n105929), .A(n81751), .ZN(n104292) );
  AOI22_X1 U66984 ( .A1(n105926), .A2(n108532), .B1(n105923), .B2(n106242), 
        .ZN(n81751) );
  OAI21_X1 U66985 ( .B1(n81299), .B2(n105929), .A(n81752), .ZN(n104293) );
  AOI22_X1 U66986 ( .A1(n105928), .A2(n107773), .B1(n105925), .B2(n81301), 
        .ZN(n81752) );
  OAI21_X1 U66987 ( .B1(n106146), .B2(n105929), .A(n81753), .ZN(n104294) );
  AOI22_X1 U66988 ( .A1(n105926), .A2(n107874), .B1(n105925), .B2(n81360), 
        .ZN(n81753) );
  OAI21_X1 U66989 ( .B1(n106254), .B2(n105929), .A(n81754), .ZN(n104295) );
  AOI22_X1 U66990 ( .A1(n74162), .A2(n105927), .B1(n105923), .B2(n81272), .ZN(
        n81754) );
  OAI21_X1 U66991 ( .B1(n106235), .B2(n105929), .A(n81755), .ZN(n104296) );
  AOI22_X1 U66992 ( .A1(n105926), .A2(n108415), .B1(n105925), .B2(n81283), 
        .ZN(n81755) );
  OAI21_X1 U66993 ( .B1(n106230), .B2(n105929), .A(n81756), .ZN(n104297) );
  AOI22_X1 U66994 ( .A1(n105928), .A2(n108181), .B1(n105923), .B2(n81286), 
        .ZN(n81756) );
  OAI21_X1 U66995 ( .B1(n106230), .B2(n105922), .A(n81758), .ZN(n104298) );
  AOI22_X1 U66996 ( .A1(n104819), .A2(n81286), .B1(n105920), .B2(n108172), 
        .ZN(n81758) );
  OAI21_X1 U66997 ( .B1(n106162), .B2(n105922), .A(n81761), .ZN(n104299) );
  AOI22_X1 U66998 ( .A1(n104819), .A2(n81347), .B1(n105920), .B2(n110025), 
        .ZN(n81761) );
  OAI21_X1 U66999 ( .B1(n106259), .B2(n105922), .A(n81762), .ZN(n104300) );
  AOI22_X1 U67000 ( .A1(n104819), .A2(n81269), .B1(n105920), .B2(n109336), 
        .ZN(n81762) );
  OAI21_X1 U67001 ( .B1(n106244), .B2(n105922), .A(n81763), .ZN(n104301) );
  AOI22_X1 U67002 ( .A1(n104820), .A2(n106240), .B1(n105920), .B2(n108523), 
        .ZN(n81763) );
  OAI21_X1 U67003 ( .B1(n106236), .B2(n105922), .A(n81764), .ZN(n104302) );
  AOI22_X1 U67004 ( .A1(n104719), .A2(n81283), .B1(n81760), .B2(n108406), .ZN(
        n81764) );
  OAI21_X1 U67005 ( .B1(n81394), .B2(n105922), .A(n81765), .ZN(n104303) );
  AOI22_X1 U67006 ( .A1(n104820), .A2(n106019), .B1(n105919), .B2(n109451), 
        .ZN(n81765) );
  OAI21_X1 U67007 ( .B1(n81349), .B2(n105922), .A(n81766), .ZN(n104304) );
  AOI22_X1 U67008 ( .A1(n104718), .A2(n81351), .B1(n105920), .B2(n109667), 
        .ZN(n81766) );
  OAI21_X1 U67009 ( .B1(n81318), .B2(n105922), .A(n81767), .ZN(n104305) );
  AOI22_X1 U67010 ( .A1(n81759), .A2(n106060), .B1(n105920), .B2(n110350), 
        .ZN(n81767) );
  OAI21_X1 U67011 ( .B1(n106146), .B2(n105922), .A(n81768), .ZN(n104306) );
  AOI22_X1 U67012 ( .A1(n104718), .A2(n81360), .B1(n105919), .B2(n107866), 
        .ZN(n81768) );
  OAI21_X1 U67013 ( .B1(n81315), .B2(n105921), .A(n81769), .ZN(n104307) );
  AOI22_X1 U67014 ( .A1(n104718), .A2(n81474), .B1(n105919), .B2(n110242), 
        .ZN(n81769) );
  OAI21_X1 U67015 ( .B1(n81299), .B2(n105921), .A(n81770), .ZN(n104308) );
  AOI22_X1 U67016 ( .A1(n104820), .A2(n81301), .B1(n105919), .B2(n107764), 
        .ZN(n81770) );
  OAI21_X1 U67017 ( .B1(n106135), .B2(n105921), .A(n81771), .ZN(n104309) );
  AOI22_X1 U67018 ( .A1(n104718), .A2(n81539), .B1(n105919), .B2(n107226), 
        .ZN(n81771) );
  OAI21_X1 U67019 ( .B1(n105219), .B2(n105921), .A(n81772), .ZN(n104310) );
  AOI22_X1 U67020 ( .A1(n104819), .A2(n80188), .B1(n105919), .B2(n108760), 
        .ZN(n81772) );
  OAI21_X1 U67021 ( .B1(n81306), .B2(n105921), .A(n81773), .ZN(n104311) );
  AOI22_X1 U67022 ( .A1(n104719), .A2(n81308), .B1(n105919), .B2(n110667), 
        .ZN(n81773) );
  OAI21_X1 U67023 ( .B1(n106259), .B2(n105917), .A(n81775), .ZN(n104312) );
  AOI22_X1 U67024 ( .A1(n72228), .A2(n105000), .B1(n105916), .B2(n81269), .ZN(
        n81775) );
  OAI21_X1 U67025 ( .B1(n106244), .B2(n105918), .A(n81778), .ZN(n104313) );
  AOI22_X1 U67026 ( .A1(n71186), .A2(n105001), .B1(n105915), .B2(n106241), 
        .ZN(n81778) );
  OAI21_X1 U67027 ( .B1(n106135), .B2(n105917), .A(n81779), .ZN(n104314) );
  AOI22_X1 U67028 ( .A1(n69490), .A2(n81776), .B1(n105915), .B2(n81539), .ZN(
        n81779) );
  OAI21_X1 U67029 ( .B1(n106254), .B2(n105917), .A(n81780), .ZN(n104315) );
  AOI22_X1 U67030 ( .A1(n74138), .A2(n105001), .B1(n105916), .B2(n81272), .ZN(
        n81780) );
  OAI21_X1 U67031 ( .B1(n111059), .B2(n105913), .A(n81782), .ZN(n104316) );
  AOI22_X1 U67032 ( .A1(n105911), .A2(n105908), .B1(n105907), .B2(n108941), 
        .ZN(n81782) );
  OAI21_X1 U67033 ( .B1(n111063), .B2(n105912), .A(n81786), .ZN(n104317) );
  AOI22_X1 U67034 ( .A1(n105909), .A2(n81269), .B1(n105907), .B2(n109405), 
        .ZN(n81786) );
  OAI21_X1 U67037 ( .B1(n105189), .B2(n104527), .A(n81788), .ZN(n104320) );
  NAND2_X1 U67038 ( .A1(n105904), .A2(n81790), .ZN(n81788) );
  OAI21_X1 U67039 ( .B1(n105188), .B2(n104526), .A(n81791), .ZN(n104321) );
  NAND2_X1 U67040 ( .A1(n105904), .A2(n81792), .ZN(n81791) );
  OAI21_X1 U67041 ( .B1(n105189), .B2(n104525), .A(n81793), .ZN(n104322) );
  NAND2_X1 U67042 ( .A1(n105904), .A2(n81794), .ZN(n81793) );
  OAI21_X1 U67043 ( .B1(n81498), .B2(n105902), .A(n81796), .ZN(n104323) );
  AOI22_X1 U67044 ( .A1(n81797), .A2(n81500), .B1(n105190), .B2(n108938), .ZN(
        n81796) );
  OAI21_X1 U67045 ( .B1(n102318), .B2(n81798), .A(n81799), .ZN(n104324) );
  AOI22_X1 U67046 ( .A1(n81797), .A2(n81590), .B1(n105903), .B2(n106012), .ZN(
        n81799) );
  OAI21_X1 U67047 ( .B1(n62189), .B2(n58728), .A(n81800), .ZN(n104325) );
  NAND2_X1 U67048 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [0]), .A2(n62189), 
        .ZN(n81800) );
  NOR2_X1 U67049 ( .A1(n105072), .A2(net67007), .ZN(n104326) );
  OAI21_X1 U67050 ( .B1(n62189), .B2(n58724), .A(n81801), .ZN(n104327) );
  NAND2_X1 U67051 ( .A1(\DLX_Datapath/next_ALUOut_EXMEM [29]), .A2(n106358), 
        .ZN(n81801) );
  AOI22_X1 U67052 ( .A1(n81803), .A2(n105097), .B1(
        \DLX_Datapath/MUX_HDU_ALUInA [29]), .B2(n81805), .ZN(n81802) );
  XNOR2_X1 U67053 ( .A(n81806), .B(n81807), .ZN(n81803) );
  AOI22_X1 U67055 ( .A1(n81810), .A2(n105097), .B1(
        \DLX_Datapath/MUX_HDU_ALUInA [30]), .B2(n81805), .ZN(n81809) );
  XNOR2_X1 U67056 ( .A(n81806), .B(n81811), .ZN(n81810) );
  AOI22_X1 U67058 ( .A1(n81814), .A2(n105096), .B1(
        \DLX_Datapath/MUX_HDU_ALUInA [31]), .B2(n81805), .ZN(n81813) );
  XNOR2_X1 U67059 ( .A(n81806), .B(n81815), .ZN(n81814) );
  OAI21_X1 U67061 ( .B1(n107556), .B2(n81817), .A(n81818), .ZN(n81816) );
  AOI21_X1 U67062 ( .B1(n81819), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[17] ), .A(n108267), .ZN(
        n81818) );
  NOR2_X1 U67063 ( .A1(n107027), .A2(n111023), .ZN(n104328) );
  OAI21_X1 U67064 ( .B1(n109771), .B2(n107951), .A(n81820), .ZN(n69975) );
  OAI21_X1 U67065 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [31]), .B2(
        \DLX_Datapath/ArithLogUnit/A_add [31]), .A(n81821), .ZN(n81820) );
  AOI21_X1 U67066 ( .B1(n81822), .B2(n110955), .A(n81823), .ZN(n81821) );
  AOI21_X1 U67067 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [30]), .B2(n107587), 
        .A(\DLX_Datapath/ArithLogUnit/B_add [30]), .ZN(n81823) );
  OAI21_X1 U67068 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [29]), .B2(n81824), 
        .A(n81825), .ZN(n81822) );
  NAND2_X1 U67069 ( .A1(n81826), .A2(n109772), .ZN(n81825) );
  NOR2_X1 U67070 ( .A1(n81826), .A2(n109772), .ZN(n81824) );
  AOI21_X1 U67071 ( .B1(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[1] ), .B2(n107591), .A(n104369), .ZN(n81826) );
  OAI21_X1 U67073 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [27]), .B2(
        \DLX_Datapath/ArithLogUnit/A_add [27]), .A(n81827), .ZN(n79720) );
  OAI21_X1 U67074 ( .B1(n110749), .B2(n108047), .A(n81828), .ZN(n81827) );
  AOI22_X1 U67075 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [26]), .A2(n81829), 
        .B1(\DLX_Datapath/ArithLogUnit/A_add [26]), .B2(n81830), .ZN(n81828)
         );
  OR2_X1 U67076 ( .A1(\DLX_Datapath/ArithLogUnit/A_add [26]), .A2(n81830), 
        .ZN(n81829) );
  AOI21_X1 U67077 ( .B1(n110953), .B2(n81831), .A(n81832), .ZN(n81830) );
  AOI21_X1 U67078 ( .B1(n107592), .B2(\DLX_Datapath/ArithLogUnit/A_add [25]), 
        .A(\DLX_Datapath/ArithLogUnit/B_add [25]), .ZN(n81832) );
  AOI21_X1 U67079 ( .B1(n107596), .B2(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[1] ), .A(n104376), .ZN(n81831) );
  AOI21_X1 U67081 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [23]), .B2(
        \DLX_Datapath/ArithLogUnit/B_add [23]), .A(n107597), .ZN(n79755) );
  OAI21_X1 U67082 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [23]), .B2(
        \DLX_Datapath/ArithLogUnit/A_add [23]), .A(n81834), .ZN(n81833) );
  AOI21_X1 U67083 ( .B1(n81835), .B2(n110331), .A(n81836), .ZN(n81834) );
  AOI21_X1 U67084 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [22]), .B2(n107598), 
        .A(\DLX_Datapath/ArithLogUnit/B_add [22]), .ZN(n81836) );
  OAI21_X1 U67085 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [21]), .B2(n81837), 
        .A(n81838), .ZN(n81835) );
  NAND2_X1 U67086 ( .A1(n81839), .A2(n110651), .ZN(n81838) );
  NOR2_X1 U67087 ( .A1(n81839), .A2(n110651), .ZN(n81837) );
  AOI21_X1 U67088 ( .B1(n79788), .B2(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[1] ), .A(n104375), .ZN(n81839) );
  OAI21_X1 U67090 ( .B1(n81840), .B2(n110118), .A(n81841), .ZN(n79788) );
  AOI21_X1 U67091 ( .B1(n81842), .B2(n81843), .A(n81844), .ZN(n81841) );
  AOI21_X1 U67092 ( .B1(n81840), .B2(n110118), .A(n109779), .ZN(n81844) );
  NOR3_X1 U67093 ( .A1(n81845), .A2(n79821), .A3(n81846), .ZN(n81843) );
  AOI21_X1 U67094 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [15]), .B2(
        \DLX_Datapath/ArithLogUnit/B_add [15]), .A(n107599), .ZN(n79821) );
  OAI21_X1 U67095 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [15]), .B2(
        \DLX_Datapath/ArithLogUnit/A_add [15]), .A(n81848), .ZN(n81847) );
  AOI21_X1 U67096 ( .B1(n81849), .B2(n109770), .A(n81850), .ZN(n81848) );
  AOI21_X1 U67097 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [14]), .B2(n107600), 
        .A(\DLX_Datapath/ArithLogUnit/B_add [14]), .ZN(n81850) );
  OAI21_X1 U67098 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [13]), .B2(n81851), 
        .A(n81852), .ZN(n81849) );
  NAND2_X1 U67099 ( .A1(n81853), .A2(n109769), .ZN(n81852) );
  NOR2_X1 U67100 ( .A1(n81853), .A2(n109769), .ZN(n81851) );
  AOI21_X1 U67101 ( .B1(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[1] ), .B2(n107604), .A(n104373), .ZN(n81853) );
  OAI21_X1 U67103 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [11]), .B2(
        \DLX_Datapath/ArithLogUnit/A_add [11]), .A(n81854), .ZN(n79854) );
  OAI21_X1 U67104 ( .B1(n108502), .B2(n108507), .A(n81855), .ZN(n81854) );
  AOI22_X1 U67105 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [10]), .A2(n81856), 
        .B1(\DLX_Datapath/ArithLogUnit/A_add [10]), .B2(n81857), .ZN(n81855)
         );
  OR2_X1 U67106 ( .A1(\DLX_Datapath/ArithLogUnit/A_add [10]), .A2(n81857), 
        .ZN(n81856) );
  AOI21_X1 U67107 ( .B1(n109764), .B2(n81858), .A(n81859), .ZN(n81857) );
  AOI21_X1 U67108 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [9]), .B2(n107605), 
        .A(\DLX_Datapath/ArithLogUnit/B_add [9]), .ZN(n81859) );
  AOI21_X1 U67109 ( .B1(n107609), .B2(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[1] ), .A(n104372), .ZN(n81858) );
  AOI21_X1 U67111 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [7]), .B2(
        \DLX_Datapath/ArithLogUnit/B_add [7]), .A(n107610), .ZN(n79887) );
  OAI21_X1 U67112 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [7]), .B2(
        \DLX_Datapath/ArithLogUnit/A_add [7]), .A(n81861), .ZN(n81860) );
  AOI21_X1 U67113 ( .B1(n81862), .B2(n109433), .A(n81863), .ZN(n81861) );
  AOI21_X1 U67114 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [6]), .B2(n107611), 
        .A(\DLX_Datapath/ArithLogUnit/B_add [6]), .ZN(n81863) );
  OAI21_X1 U67115 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [5]), .B2(n81864), 
        .A(n81865), .ZN(n81862) );
  NAND2_X1 U67116 ( .A1(n81866), .A2(n109315), .ZN(n81865) );
  NOR2_X1 U67117 ( .A1(n81866), .A2(n109315), .ZN(n81864) );
  AOI21_X1 U67118 ( .B1(n107615), .B2(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[1] ), .A(n104370), .ZN(n81866) );
  AOI21_X1 U67120 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [3]), .B2(
        \DLX_Datapath/ArithLogUnit/B_add [3]), .A(n107616), .ZN(n79920) );
  OAI21_X1 U67121 ( .B1(\DLX_Datapath/ArithLogUnit/B_add [3]), .B2(
        \DLX_Datapath/ArithLogUnit/A_add [3]), .A(n81868), .ZN(n81867) );
  AOI21_X1 U67122 ( .B1(n81869), .B2(n108969), .A(n81870), .ZN(n81868) );
  AOI21_X1 U67123 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [2]), .B2(n107617), 
        .A(\DLX_Datapath/ArithLogUnit/B_add [2]), .ZN(n81870) );
  OAI21_X1 U67124 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [1]), .B2(n107619), 
        .A(n107618), .ZN(n81869) );
  AOI21_X1 U67125 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [1]), .B2(n107619), 
        .A(\DLX_Datapath/ArithLogUnit/B_add [1]), .ZN(n81871) );
  OAI21_X1 U67126 ( .B1(\DLX_Datapath/ArithLogUnit/Cin_add ), .B2(n104367), 
        .A(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[1] ), .ZN(n81872) );
  NOR2_X1 U67127 ( .A1(n108858), .A2(n107620), .ZN(n104367) );
  NOR2_X1 U67128 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [17]), .A2(
        \DLX_Datapath/ArithLogUnit/A_add [17]), .ZN(n81845) );
  AOI22_X1 U67129 ( .A1(n110225), .A2(n109781), .B1(n110118), .B2(n109779), 
        .ZN(n81842) );
  AOI21_X1 U67130 ( .B1(n109892), .B2(\DLX_Datapath/ArithLogUnit/A_add [18]), 
        .A(n81873), .ZN(n81840) );
  AOI21_X1 U67131 ( .B1(n81874), .B2(n110225), .A(n109781), .ZN(n81873) );
  OAI21_X1 U67132 ( .B1(\DLX_Datapath/ArithLogUnit/A_add [17]), .B2(n104374), 
        .A(n109893), .ZN(n81874) );
  AOI21_X1 U67133 ( .B1(n104374), .B2(\DLX_Datapath/ArithLogUnit/A_add [17]), 
        .A(\DLX_Datapath/ArithLogUnit/B_add [17]), .ZN(n81875) );
  NOR2_X1 U67135 ( .A1(net113157), .A2(n104501), .ZN(n64127) );
  NOR2_X1 U67136 ( .A1(net113155), .A2(n107130), .ZN(n64126) );
  NOR2_X1 U67137 ( .A1(n105029), .A2(n100801), .ZN(n62664) );
  OAI21_X1 U67140 ( .B1(n107021), .B2(n81879), .A(n81880), .ZN(n60377) );
  NAND2_X1 U67141 ( .A1(n81881), .A2(n81882), .ZN(n81880) );
  OAI21_X1 U67143 ( .B1(net113091), .B2(n106957), .A(n81884), .ZN(n60376) );
  NAND2_X1 U67144 ( .A1(n81885), .A2(n81886), .ZN(n81884) );
  NOR4_X1 U67145 ( .A1(IR_in[24]), .A2(n105152), .A3(n111150), .A4(n111153), 
        .ZN(n81886) );
  NOR3_X1 U67146 ( .A1(n81887), .A2(n111152), .A3(n111151), .ZN(n81885) );
  OAI21_X1 U67147 ( .B1(n107023), .B2(n81879), .A(n81888), .ZN(n60375) );
  XOR2_X1 U67149 ( .A(n107096), .B(n106696), .Z(n60374) );
  OAI21_X1 U67150 ( .B1(n69283), .B2(n81890), .A(n81891), .ZN(n60373) );
  AOI22_X1 U67151 ( .A1(n81892), .A2(n106696), .B1(n81893), .B2(n104898), .ZN(
        n81891) );
  NOR2_X1 U67152 ( .A1(n81894), .A2(n104898), .ZN(n81892) );
  XOR2_X1 U67153 ( .A(n106695), .B(n59516), .Z(n81894) );
  OAI21_X1 U67154 ( .B1(n81895), .B2(n81896), .A(n81897), .ZN(n60372) );
  OAI21_X1 U67155 ( .B1(n81893), .B2(n81898), .A(\DLX_Datapath/CWP_IDEX[2] ), 
        .ZN(n81897) );
  OAI21_X1 U67156 ( .B1(n69283), .B2(n105012), .A(n107099), .ZN(n81898) );
  OAI21_X1 U67157 ( .B1(n107096), .B2(n106695), .A(n106696), .ZN(n81893) );
  OR2_X1 U67158 ( .A1(n81900), .A2(\DLX_Datapath/CWP_IDEX[2] ), .ZN(n81896) );
  AOI22_X1 U67159 ( .A1(n81901), .A2(n106695), .B1(n69283), .B2(n105052), .ZN(
        n81900) );
  XOR2_X1 U67160 ( .A(n81902), .B(
        \dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .Z(n60371) );
  OAI21_X1 U67161 ( .B1(n81882), .B2(n81903), .A(n106696), .ZN(n81902) );
  XOR2_X1 U67162 ( .A(n106764), .B(n81904), .Z(n60370) );
  AOI21_X1 U67163 ( .B1(n106517), .B2(n107027), .A(n81905), .ZN(n81904) );
  OAI21_X1 U67164 ( .B1(n59515), .B2(n81906), .A(n81907), .ZN(n60369) );
  NAND2_X1 U67165 ( .A1(n106696), .A2(n81908), .ZN(n81907) );
  OAI21_X1 U67166 ( .B1(n69283), .B2(n81909), .A(n81910), .ZN(n81908) );
  AOI22_X1 U67167 ( .A1(n81911), .A2(n107027), .B1(n81912), .B2(n81882), .ZN(
        n81910) );
  OAI21_X1 U67168 ( .B1(n106517), .B2(n81913), .A(n81914), .ZN(n81911) );
  NAND2_X1 U67169 ( .A1(n59515), .A2(n106764), .ZN(n81913) );
  AOI21_X1 U67170 ( .B1(n69283), .B2(n81915), .A(n81905), .ZN(n81906) );
  OAI21_X1 U67171 ( .B1(n81882), .B2(n107027), .A(n106696), .ZN(n81905) );
  NAND2_X1 U67172 ( .A1(n81889), .A2(n81883), .ZN(n81895) );
  NAND2_X1 U67173 ( .A1(n81916), .A2(n106958), .ZN(n81883) );
  NOR2_X1 U67174 ( .A1(n69340), .A2(n69283), .ZN(n81916) );
  OAI21_X1 U67175 ( .B1(net113081), .B2(n106942), .A(n81917), .ZN(n60368) );
  AOI21_X1 U67176 ( .B1(IR_in[26]), .B2(net113091), .A(n81918), .ZN(n81917) );
  OAI21_X1 U67177 ( .B1(n104753), .B2(n106936), .A(n81919), .ZN(n60367) );
  AOI21_X1 U67178 ( .B1(IR_in[28]), .B2(net113081), .A(n81918), .ZN(n81919) );
  OAI21_X1 U67179 ( .B1(net113091), .B2(n106847), .A(n81920), .ZN(n60366) );
  AOI21_X1 U67180 ( .B1(IR_in[30]), .B2(net113091), .A(n81918), .ZN(n81920) );
  NOR2_X1 U67181 ( .A1(net113156), .A2(n104788), .ZN(n81918) );
  OAI21_X1 U67182 ( .B1(net113081), .B2(n111032), .A(n106597), .ZN(n60365) );
  OAI21_X1 U67183 ( .B1(net113091), .B2(n111031), .A(n106597), .ZN(n60364) );
  OAI21_X1 U67184 ( .B1(n104753), .B2(n111030), .A(n106597), .ZN(n60362) );
  OAI21_X1 U67185 ( .B1(net113102), .B2(n111029), .A(n106597), .ZN(n60360) );
  OAI21_X1 U67186 ( .B1(net113091), .B2(n107151), .A(n106597), .ZN(n60358) );
  NOR2_X1 U67187 ( .A1(n105150), .A2(n81922), .ZN(n80097) );
  OAI21_X1 U67188 ( .B1(n104564), .B2(n81923), .A(n81924), .ZN(n60356) );
  OR2_X1 U67189 ( .A1(n105898), .A2(n100648), .ZN(n81924) );
  OAI21_X1 U67190 ( .B1(n104563), .B2(n81923), .A(n81926), .ZN(n60355) );
  OR2_X1 U67191 ( .A1(n105898), .A2(n100647), .ZN(n81926) );
  OAI21_X1 U67192 ( .B1(n107110), .B2(n81923), .A(n81927), .ZN(n60354) );
  OR2_X1 U67193 ( .A1(n105898), .A2(n100646), .ZN(n81927) );
  OAI21_X1 U67194 ( .B1(n104562), .B2(n81923), .A(n81928), .ZN(n60353) );
  OR2_X1 U67195 ( .A1(n105898), .A2(n100645), .ZN(n81928) );
  OAI21_X1 U67196 ( .B1(n104561), .B2(n81923), .A(n81929), .ZN(n60352) );
  OR2_X1 U67197 ( .A1(n105898), .A2(n100644), .ZN(n81929) );
  OAI21_X1 U67198 ( .B1(n104560), .B2(n81923), .A(n81930), .ZN(n60351) );
  OR2_X1 U67199 ( .A1(n105898), .A2(n100643), .ZN(n81930) );
  OAI21_X1 U67200 ( .B1(n107111), .B2(n81923), .A(n81931), .ZN(n60350) );
  OR2_X1 U67201 ( .A1(n105898), .A2(n100642), .ZN(n81931) );
  OAI21_X1 U67202 ( .B1(n104559), .B2(n81923), .A(n81932), .ZN(n60349) );
  OR2_X1 U67203 ( .A1(n105898), .A2(n100641), .ZN(n81932) );
  OAI21_X1 U67204 ( .B1(n107112), .B2(n81923), .A(n81933), .ZN(n60348) );
  OR2_X1 U67205 ( .A1(n81925), .A2(n100640), .ZN(n81933) );
  OAI21_X1 U67206 ( .B1(n104558), .B2(n81923), .A(n81934), .ZN(n60347) );
  OR2_X1 U67207 ( .A1(n105898), .A2(n100639), .ZN(n81934) );
  OAI21_X1 U67208 ( .B1(n104557), .B2(n81923), .A(n81935), .ZN(n60346) );
  OR2_X1 U67209 ( .A1(n105898), .A2(n100638), .ZN(n81935) );
  OAI21_X1 U67210 ( .B1(n104580), .B2(n105898), .A(n81936), .ZN(n60345) );
  AOI21_X1 U67211 ( .B1(n105154), .B2(n69349), .A(n81938), .ZN(n81936) );
  OAI21_X1 U67212 ( .B1(n104579), .B2(n105898), .A(n81939), .ZN(n60344) );
  AOI21_X1 U67213 ( .B1(n105154), .B2(n69350), .A(n81938), .ZN(n81939) );
  OAI21_X1 U67214 ( .B1(n104578), .B2(n105898), .A(n81940), .ZN(n60343) );
  AOI21_X1 U67215 ( .B1(n105154), .B2(n69351), .A(n81938), .ZN(n81940) );
  OAI21_X1 U67216 ( .B1(n104577), .B2(n105898), .A(n81941), .ZN(n60342) );
  AOI21_X1 U67217 ( .B1(n81937), .B2(n69352), .A(n81938), .ZN(n81941) );
  OAI21_X1 U67218 ( .B1(n104576), .B2(n105898), .A(n81942), .ZN(n60341) );
  AOI21_X1 U67219 ( .B1(n105154), .B2(n69353), .A(n81938), .ZN(n81942) );
  OAI21_X1 U67220 ( .B1(n104575), .B2(n81925), .A(n81943), .ZN(n60340) );
  AOI21_X1 U67221 ( .B1(n105154), .B2(n69354), .A(n81938), .ZN(n81943) );
  OAI21_X1 U67222 ( .B1(n104574), .B2(n81925), .A(n81944), .ZN(n60339) );
  AOI21_X1 U67223 ( .B1(n105154), .B2(n69355), .A(n81938), .ZN(n81944) );
  OAI21_X1 U67224 ( .B1(n104573), .B2(n81925), .A(n81945), .ZN(n60338) );
  AOI21_X1 U67225 ( .B1(n81937), .B2(n69356), .A(n81938), .ZN(n81945) );
  OAI21_X1 U67226 ( .B1(n104572), .B2(n81925), .A(n81946), .ZN(n60337) );
  AOI21_X1 U67227 ( .B1(n105154), .B2(n69357), .A(n81938), .ZN(n81946) );
  OAI21_X1 U67228 ( .B1(n104571), .B2(n81925), .A(n81947), .ZN(n60336) );
  AOI21_X1 U67229 ( .B1(n105154), .B2(n69358), .A(n81938), .ZN(n81947) );
  OAI21_X1 U67230 ( .B1(n104570), .B2(n81925), .A(n81948), .ZN(n60335) );
  AOI21_X1 U67231 ( .B1(n105154), .B2(n69359), .A(n81938), .ZN(n81948) );
  OAI21_X1 U67232 ( .B1(n104569), .B2(n81925), .A(n81949), .ZN(n60334) );
  AOI21_X1 U67233 ( .B1(n105154), .B2(\DLX_Datapath/IR_IFID[11] ), .A(n81938), 
        .ZN(n81949) );
  OAI21_X1 U67234 ( .B1(n104568), .B2(n81925), .A(n81950), .ZN(n60333) );
  AOI21_X1 U67235 ( .B1(n105154), .B2(\DLX_Datapath/IR_IFID[12] ), .A(n81938), 
        .ZN(n81950) );
  OAI21_X1 U67236 ( .B1(n104567), .B2(n81925), .A(n81951), .ZN(n60332) );
  AOI21_X1 U67237 ( .B1(n81937), .B2(\DLX_Datapath/IR_IFID[13] ), .A(n81938), 
        .ZN(n81951) );
  OAI21_X1 U67238 ( .B1(n104566), .B2(n81925), .A(n81952), .ZN(n60331) );
  AOI21_X1 U67239 ( .B1(n105154), .B2(n69362), .A(n81938), .ZN(n81952) );
  OAI21_X1 U67240 ( .B1(n104565), .B2(n81925), .A(n81953), .ZN(n60330) );
  AOI21_X1 U67241 ( .B1(n105154), .B2(n69369), .A(n81938), .ZN(n81953) );
  AND2_X2 U67242 ( .A1(n81954), .A2(n61670), .ZN(n81938) );
  NOR2_X1 U67243 ( .A1(n107130), .A2(n81923), .ZN(n81954) );
  NOR2_X1 U67244 ( .A1(n81955), .A2(n107421), .ZN(n81937) );
  NAND2_X1 U67245 ( .A1(n81925), .A2(net113102), .ZN(n81955) );
  NAND2_X1 U67246 ( .A1(n81956), .A2(n81957), .ZN(n60329) );
  AOI21_X1 U67247 ( .B1(n81958), .B2(net67007), .A(n81959), .ZN(n81957) );
  NOR3_X1 U67248 ( .A1(n81960), .A2(IR_in[3]), .A3(n81961), .ZN(n81959) );
  AOI21_X1 U67249 ( .B1(n81962), .B2(net112601), .A(n81963), .ZN(n81961) );
  OAI33_X1 U67250 ( .A1(net67007), .A2(n111157), .A3(n111160), .B1(n81964), 
        .B2(IR_in[0]), .B3(n81965), .ZN(n81963) );
  OR2_X1 U67251 ( .A1(IR_in[5]), .A2(IR_in[6]), .ZN(n81964) );
  AOI22_X1 U67252 ( .A1(n105165), .A2(n111120), .B1(net113157), .B2(n111034), 
        .ZN(n81956) );
  NOR4_X1 U67253 ( .A1(n81969), .A2(n81970), .A3(n111125), .A4(n81971), .ZN(
        n81968) );
  OAI21_X1 U67254 ( .B1(n81973), .B2(n81974), .A(n111145), .ZN(n81972) );
  AOI21_X1 U67255 ( .B1(n81975), .B2(n80064), .A(n81976), .ZN(n81970) );
  NOR3_X1 U67256 ( .A1(n81977), .A2(IR_in[0]), .A3(n81965), .ZN(n81969) );
  NAND2_X1 U67257 ( .A1(n81978), .A2(n81979), .ZN(n60328) );
  AOI22_X1 U67258 ( .A1(n81980), .A2(IR_in[0]), .B1(n104809), .B2(n81966), 
        .ZN(n81979) );
  OAI21_X1 U67259 ( .B1(IR_in[1]), .B2(n81967), .A(n81982), .ZN(n81966) );
  NAND2_X1 U67260 ( .A1(n81983), .A2(IR_in[1]), .ZN(n81982) );
  NOR2_X1 U67261 ( .A1(IR_in[6]), .A2(IR_in[5]), .ZN(n81983) );
  AOI22_X1 U67262 ( .A1(n105164), .A2(n81984), .B1(net113156), .B2(n111033), 
        .ZN(n81978) );
  NAND2_X1 U67263 ( .A1(n81985), .A2(n81986), .ZN(n81984) );
  AOI21_X1 U67264 ( .B1(n111148), .B2(n81974), .A(n81971), .ZN(n81986) );
  NAND2_X1 U67265 ( .A1(n81987), .A2(n81988), .ZN(n81971) );
  AOI22_X1 U67266 ( .A1(n81989), .A2(n111139), .B1(n81974), .B2(n111147), .ZN(
        n81988) );
  NOR2_X1 U67267 ( .A1(n111121), .A2(n81990), .ZN(n81987) );
  AOI22_X1 U67269 ( .A1(n81992), .A2(n111138), .B1(n80042), .B2(n81973), .ZN(
        n81991) );
  NAND2_X1 U67270 ( .A1(n81993), .A2(n111126), .ZN(n81973) );
  NOR2_X1 U67271 ( .A1(net67007), .A2(n81965), .ZN(n81992) );
  NAND2_X1 U67272 ( .A1(n81995), .A2(n81994), .ZN(n60327) );
  NOR3_X1 U67273 ( .A1(n81996), .A2(n81958), .A3(n81980), .ZN(n81995) );
  NAND2_X1 U67280 ( .A1(n82001), .A2(n111139), .ZN(n81960) );
  NOR2_X1 U67281 ( .A1(IR_in[4]), .A2(n105152), .ZN(n82001) );
  NAND2_X1 U67282 ( .A1(n111159), .A2(IR_in[2]), .ZN(n82000) );
  AOI22_X1 U67283 ( .A1(n105162), .A2(n82002), .B1(net113157), .B2(
        \DLX_ControlUnit/ALUop2 [3]), .ZN(n81994) );
  NAND2_X1 U67284 ( .A1(n82003), .A2(n82004), .ZN(n82002) );
  NOR3_X1 U67285 ( .A1(n82005), .A2(n82006), .A3(n111122), .ZN(n82004) );
  AOI21_X1 U67286 ( .B1(n111128), .B2(n111148), .A(n81990), .ZN(n82003) );
  OAI21_X1 U67287 ( .B1(n81975), .B2(n111126), .A(n82007), .ZN(n81990) );
  AOI22_X1 U67288 ( .A1(n105162), .A2(n82009), .B1(net113157), .B2(
        \DLX_ControlUnit/ALUop2 [4]), .ZN(n82008) );
  NAND2_X1 U67289 ( .A1(n82010), .A2(n82011), .ZN(n82009) );
  AOI22_X1 U67290 ( .A1(n82012), .A2(n111138), .B1(n81989), .B2(n111139), .ZN(
        n82011) );
  NOR4_X1 U67292 ( .A1(IR_in[5]), .A2(IR_in[4]), .A3(IR_in[3]), .A4(IR_in[2]), 
        .ZN(n82014) );
  AOI21_X1 U67295 ( .B1(n111128), .B2(n111147), .A(n82016), .ZN(n82010) );
  OR2_X1 U67296 ( .A1(n82017), .A2(n82018), .ZN(n60325) );
  OAI21_X1 U67297 ( .B1(n100462), .B2(n82019), .A(n82020), .ZN(n82018) );
  AOI22_X1 U67298 ( .A1(n104706), .A2(n106772), .B1(n82022), .B2(DataAddr[0]), 
        .ZN(n82020) );
  AOI22_X1 U67300 ( .A1(n82026), .A2(PC_out[0]), .B1(n105891), .B2(n108615), 
        .ZN(n82025) );
  OR2_X1 U67301 ( .A1(n82028), .A2(n82029), .ZN(n60324) );
  OAI21_X1 U67302 ( .B1(n100460), .B2(n82019), .A(n82030), .ZN(n82029) );
  AOI22_X1 U67303 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 [1]), 
        .A2(n104706), .B1(n82022), .B2(DataAddr[1]), .ZN(n82030) );
  AOI22_X1 U67305 ( .A1(n82026), .A2(PC_out[1]), .B1(n105893), .B2(n108616), 
        .ZN(n82031) );
  OR2_X1 U67307 ( .A1(n82034), .A2(n82033), .ZN(n60323) );
  OAI21_X1 U67308 ( .B1(n105078), .B2(net113091), .A(n82035), .ZN(n82034) );
  AOI22_X1 U67309 ( .A1(n105895), .A2(DataAddr[2]), .B1(n105156), .B2(n108621), 
        .ZN(n82035) );
  NAND2_X1 U67310 ( .A1(n82036), .A2(n82037), .ZN(n82033) );
  AOI22_X1 U67311 ( .A1(n105891), .A2(n108617), .B1(n105045), .B2(n105078), 
        .ZN(n82037) );
  AOI22_X1 U67312 ( .A1(n105158), .A2(\DLX_Datapath/next_A_IDEX[2] ), .B1(
        \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 [2]), .B2(n104706), .ZN(
        n82036) );
  OR2_X1 U67313 ( .A1(n82038), .A2(n82039), .ZN(n60322) );
  AOI22_X1 U67315 ( .A1(n105895), .A2(DataAddr[3]), .B1(n105156), .B2(n108631), 
        .ZN(n82040) );
  NAND2_X1 U67316 ( .A1(n82041), .A2(n82042), .ZN(n82038) );
  AOI22_X1 U67317 ( .A1(n105891), .A2(n108618), .B1(n105045), .B2(n82043), 
        .ZN(n82042) );
  AOI22_X1 U67318 ( .A1(n105158), .A2(\DLX_Datapath/next_A_IDEX[3] ), .B1(
        \DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 [3]), .B2(n104706), .ZN(
        n82041) );
  OR2_X1 U67319 ( .A1(n82045), .A2(n82044), .ZN(n60321) );
  OAI21_X1 U67320 ( .B1(net2465400), .B2(n104753), .A(n82046), .ZN(n82045) );
  AOI22_X1 U67321 ( .A1(n105895), .A2(DataAddr[4]), .B1(n105156), .B2(n109092), 
        .ZN(n82046) );
  NAND2_X1 U67322 ( .A1(n82047), .A2(n82048), .ZN(n82044) );
  AOI22_X1 U67323 ( .A1(n105897), .A2(n106799), .B1(n105893), .B2(n109316), 
        .ZN(n82048) );
  XOR2_X1 U67324 ( .A(n106800), .B(n82049), .Z(n80139) );
  XOR2_X1 U67325 ( .A(net2465400), .B(IR_in[4]), .Z(n82049) );
  AOI22_X1 U67326 ( .A1(n82050), .A2(n105890), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[4] ), .ZN(n82047) );
  OR2_X1 U67327 ( .A1(n82051), .A2(n82052), .ZN(n60320) );
  OAI21_X1 U67328 ( .B1(n62201), .B2(net113091), .A(n82053), .ZN(n82052) );
  AOI22_X1 U67329 ( .A1(n105894), .A2(DataAddr[5]), .B1(n105157), .B2(n109094), 
        .ZN(n82053) );
  NAND2_X1 U67330 ( .A1(n82054), .A2(n82055), .ZN(n82051) );
  AOI22_X1 U67331 ( .A1(n105896), .A2(n106798), .B1(n105893), .B2(n109321), 
        .ZN(n82055) );
  AOI22_X1 U67332 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_0 [1]), 
        .A2(n82056), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_1 [1]), 
        .B2(n106800), .ZN(n80107) );
  AOI22_X1 U67333 ( .A1(n82057), .A2(n105050), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[5] ), .ZN(n82054) );
  OR2_X1 U67334 ( .A1(n82058), .A2(n82059), .ZN(n60319) );
  OAI21_X1 U67335 ( .B1(n62200), .B2(net113091), .A(n82060), .ZN(n82059) );
  AOI22_X1 U67336 ( .A1(n105894), .A2(DataAddr[6]), .B1(n105157), .B2(n109096), 
        .ZN(n82060) );
  NAND2_X1 U67337 ( .A1(n82061), .A2(n82062), .ZN(n82058) );
  AOI22_X1 U67338 ( .A1(n104706), .A2(n106797), .B1(n105893), .B2(n109322), 
        .ZN(n82062) );
  AOI22_X1 U67339 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_0 [2]), 
        .A2(n82056), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_1 [2]), 
        .B2(n106800), .ZN(n80109) );
  AOI22_X1 U67340 ( .A1(n82063), .A2(n105050), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[6] ), .ZN(n82061) );
  OR2_X1 U67341 ( .A1(n82064), .A2(n82065), .ZN(n60318) );
  OAI21_X1 U67342 ( .B1(n62183), .B2(net113091), .A(n82066), .ZN(n82065) );
  AOI22_X1 U67343 ( .A1(n105894), .A2(DataAddr[7]), .B1(n105157), .B2(n108972), 
        .ZN(n82066) );
  NAND2_X1 U67344 ( .A1(n82067), .A2(n82068), .ZN(n82064) );
  AOI22_X1 U67345 ( .A1(n105896), .A2(n106796), .B1(n105893), .B2(n109323), 
        .ZN(n82068) );
  AOI22_X1 U67346 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_0 [3]), 
        .A2(n82056), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/S_1 [3]), 
        .B2(n106800), .ZN(n80111) );
  AOI21_X1 U67347 ( .B1(IR_in[2]), .B2(n105076), .A(n82070), .ZN(n82056) );
  OR2_X1 U67348 ( .A1(n82071), .A2(n82072), .ZN(n82070) );
  AOI21_X1 U67349 ( .B1(n82073), .B2(n104912), .A(n111159), .ZN(n82072) );
  AOI22_X1 U67350 ( .A1(n82074), .A2(n106813), .B1(IR_in[2]), .B2(PC_out[2]), 
        .ZN(n82073) );
  NOR2_X1 U67351 ( .A1(n82076), .A2(n104835), .ZN(n82074) );
  NOR4_X1 U67352 ( .A1(n104912), .A2(n82076), .A3(n104835), .A4(n104857), .ZN(
        n82071) );
  AOI22_X1 U67353 ( .A1(n82078), .A2(n105050), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[7] ), .ZN(n82067) );
  OR2_X1 U67354 ( .A1(n82079), .A2(n82080), .ZN(n60317) );
  OAI21_X1 U67355 ( .B1(n62202), .B2(net113102), .A(n82081), .ZN(n82080) );
  AOI22_X1 U67356 ( .A1(n105894), .A2(DataAddr[8]), .B1(n105157), .B2(n109435), 
        .ZN(n82081) );
  NAND2_X1 U67357 ( .A1(n82082), .A2(n82083), .ZN(n82079) );
  AOI22_X1 U67358 ( .A1(n105897), .A2(n106795), .B1(n105893), .B2(n109547), 
        .ZN(n82083) );
  XOR2_X1 U67359 ( .A(n82084), .B(n104738), .Z(n80131) );
  XOR2_X1 U67360 ( .A(IR_in[8]), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [0]), .Z(n82084) );
  AOI22_X1 U67361 ( .A1(n82085), .A2(n105050), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[8] ), .ZN(n82082) );
  OR2_X1 U67362 ( .A1(n82087), .A2(n82086), .ZN(n60316) );
  OAI21_X1 U67363 ( .B1(n104502), .B2(net113091), .A(n82088), .ZN(n82087) );
  AOI22_X1 U67364 ( .A1(n105895), .A2(DataAddr[9]), .B1(n105157), .B2(n109437), 
        .ZN(n82088) );
  NAND2_X1 U67365 ( .A1(n82089), .A2(n82090), .ZN(n82086) );
  AOI22_X1 U67366 ( .A1(n105896), .A2(n106794), .B1(n105893), .B2(n109548), 
        .ZN(n82090) );
  AOI22_X1 U67367 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_0 [1]), 
        .A2(n104738), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_1 [1]), 
        .B2(n82091), .ZN(n80141) );
  AOI22_X1 U67368 ( .A1(n82092), .A2(n105889), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[9] ), .ZN(n82089) );
  OR2_X1 U67369 ( .A1(n82094), .A2(n82093), .ZN(n60315) );
  AOI22_X1 U67371 ( .A1(n105895), .A2(DataAddr[10]), .B1(n105156), .B2(n108508), .ZN(n82095) );
  NAND2_X1 U67372 ( .A1(n82096), .A2(n82097), .ZN(n82093) );
  AOI22_X1 U67373 ( .A1(n105897), .A2(n106793), .B1(n105893), .B2(n109549), 
        .ZN(n82097) );
  AOI22_X1 U67374 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_0 [2]), 
        .A2(n104738), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_1 [2]), 
        .B2(n82091), .ZN(n80113) );
  AOI22_X1 U67375 ( .A1(n104507), .A2(n105890), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[10] ), .ZN(n82096) );
  OR2_X1 U67376 ( .A1(n82100), .A2(n82099), .ZN(n60314) );
  OAI21_X1 U67377 ( .B1(n104499), .B2(n104753), .A(n82101), .ZN(n82100) );
  AOI22_X1 U67378 ( .A1(n105895), .A2(DataAddr[11]), .B1(n105157), .B2(n107621), .ZN(n82101) );
  NAND2_X1 U67379 ( .A1(n82102), .A2(n82103), .ZN(n82099) );
  AOI22_X1 U67380 ( .A1(n105897), .A2(n106792), .B1(n105892), .B2(n106842), 
        .ZN(n82103) );
  AOI22_X1 U67381 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_0 [3]), 
        .A2(n104738), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_2/S_1 [3]), 
        .B2(n82091), .ZN(n80101) );
  AOI22_X1 U67382 ( .A1(n82104), .A2(n105889), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[11] ), .ZN(n82102) );
  OR2_X1 U67383 ( .A1(n82105), .A2(n82106), .ZN(n60313) );
  AOI22_X1 U67385 ( .A1(n105895), .A2(DataAddr[12]), .B1(n105156), .B2(n108276), .ZN(n82107) );
  NAND2_X1 U67386 ( .A1(n82108), .A2(n82109), .ZN(n82105) );
  AOI22_X1 U67387 ( .A1(n105896), .A2(n80134), .B1(n105892), .B2(n109774), 
        .ZN(n82109) );
  XOR2_X1 U67388 ( .A(net112354), .B(n82111), .Z(n80134) );
  XOR2_X1 U67389 ( .A(n104494), .B(IR_in[12]), .Z(n82111) );
  AOI22_X1 U67390 ( .A1(n82112), .A2(n105050), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[12] ), .ZN(n82108) );
  OR2_X1 U67391 ( .A1(n82114), .A2(n82113), .ZN(n60312) );
  OAI21_X1 U67392 ( .B1(n62194), .B2(n104753), .A(n82115), .ZN(n82114) );
  AOI22_X1 U67393 ( .A1(n105895), .A2(DataAddr[13]), .B1(n105156), .B2(n108278), .ZN(n82115) );
  NAND2_X1 U67394 ( .A1(n82116), .A2(n82117), .ZN(n82113) );
  AOI22_X1 U67395 ( .A1(n105897), .A2(n106790), .B1(n105892), .B2(n109775), 
        .ZN(n82117) );
  AOI22_X1 U67396 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_1 [1]), 
        .A2(net112358), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_0 [1]), 
        .B2(net112354), .ZN(n80143) );
  AOI22_X1 U67397 ( .A1(n106821), .A2(n105890), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[13] ), .ZN(n82116) );
  OR2_X1 U67398 ( .A1(n82119), .A2(n82118), .ZN(n60311) );
  OAI21_X1 U67399 ( .B1(n62199), .B2(n104753), .A(n82120), .ZN(n82119) );
  AOI22_X1 U67400 ( .A1(n105895), .A2(DataAddr[14]), .B1(n105156), .B2(n108280), .ZN(n82120) );
  NAND2_X1 U67401 ( .A1(n82121), .A2(n82122), .ZN(n82118) );
  AOI22_X1 U67402 ( .A1(n105897), .A2(n106789), .B1(n105892), .B2(n109776), 
        .ZN(n82122) );
  AOI22_X1 U67403 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_1 [2]), 
        .A2(net112358), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_0 [2]), 
        .B2(net112354), .ZN(n80115) );
  AOI22_X1 U67404 ( .A1(n82123), .A2(n105051), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[14] ), .ZN(n82121) );
  OR2_X1 U67405 ( .A1(n82124), .A2(n82125), .ZN(n60310) );
  OAI21_X1 U67406 ( .B1(n62182), .B2(n104753), .A(n82126), .ZN(n82125) );
  AOI22_X1 U67407 ( .A1(n105894), .A2(DataAddr[15]), .B1(n105156), .B2(n108158), .ZN(n82126) );
  NAND2_X1 U67408 ( .A1(n82127), .A2(n82128), .ZN(n82124) );
  AOI22_X1 U67409 ( .A1(n105896), .A2(n106788), .B1(n105892), .B2(n109777), 
        .ZN(n82128) );
  AOI22_X1 U67410 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_1 [3]), 
        .A2(net112358), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/S_0 [3]), 
        .B2(net112354), .ZN(n80117) );
  AOI22_X1 U67411 ( .A1(n106820), .A2(n105890), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[15] ), .ZN(n82127) );
  OR2_X1 U67412 ( .A1(n82130), .A2(n82129), .ZN(n60309) );
  OAI21_X1 U67413 ( .B1(n59471), .B2(net113081), .A(n82131), .ZN(n82130) );
  AOI22_X1 U67414 ( .A1(n105895), .A2(DataAddr[16]), .B1(n105157), .B2(n109899), .ZN(n82131) );
  NAND2_X1 U67415 ( .A1(n82132), .A2(n82133), .ZN(n82129) );
  AOI22_X1 U67416 ( .A1(n104706), .A2(n80146), .B1(n105892), .B2(n109897), 
        .ZN(n82133) );
  XOR2_X1 U67417 ( .A(n82134), .B(n106777), .Z(n80146) );
  XNOR2_X1 U67418 ( .A(n82135), .B(n59471), .ZN(n82134) );
  AOI22_X1 U67419 ( .A1(n82136), .A2(n105889), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[16] ), .ZN(n82132) );
  OR2_X1 U67420 ( .A1(n82137), .A2(n82138), .ZN(n60308) );
  OAI21_X1 U67421 ( .B1(n59472), .B2(net113091), .A(n82139), .ZN(n82138) );
  AOI22_X1 U67422 ( .A1(n105894), .A2(DataAddr[17]), .B1(n105157), .B2(n109901), .ZN(n82139) );
  NAND2_X1 U67423 ( .A1(n82140), .A2(n82141), .ZN(n82137) );
  AOI22_X1 U67424 ( .A1(n105897), .A2(n106775), .B1(n105892), .B2(n109898), 
        .ZN(n82141) );
  AOI22_X1 U67425 ( .A1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/S_0[1] ), 
        .A2(n106777), .B1(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/S_1[1] ), 
        .B2(n104893), .ZN(n80119) );
  AOI22_X1 U67426 ( .A1(n106819), .A2(n105050), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[17] ), .ZN(n82140) );
  OR2_X1 U67427 ( .A1(n82144), .A2(n82143), .ZN(n60307) );
  AOI22_X1 U67429 ( .A1(n105895), .A2(DataAddr[18]), .B1(n105156), .B2(n109783), .ZN(n82145) );
  NAND2_X1 U67430 ( .A1(n82147), .A2(n82146), .ZN(n82143) );
  AOI22_X1 U67431 ( .A1(n105897), .A2(n106774), .B1(n105892), .B2(n107744), 
        .ZN(n82147) );
  OAI21_X1 U67432 ( .B1(n82148), .B2(n107746), .A(n82149), .ZN(n80129) );
  NAND2_X1 U67433 ( .A1(n82150), .A2(n82148), .ZN(n82149) );
  OAI21_X1 U67435 ( .B1(n106777), .B2(n109782), .A(n82152), .ZN(n82148) );
  NAND2_X1 U67436 ( .A1(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[2] ), .A2(n106777), .ZN(n82152) );
  AOI22_X1 U67437 ( .A1(n82153), .A2(n105890), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[18] ), .ZN(n82146) );
  OR2_X1 U67438 ( .A1(n82155), .A2(n82154), .ZN(n60306) );
  OAI21_X1 U67439 ( .B1(n57424), .B2(net113091), .A(n82156), .ZN(n82155) );
  AOI22_X1 U67440 ( .A1(n105895), .A2(DataAddr[19]), .B1(n105157), .B2(n106822), .ZN(n82156) );
  NAND2_X1 U67441 ( .A1(n82157), .A2(n82158), .ZN(n82154) );
  AOI22_X1 U67442 ( .A1(n104706), .A2(n80122), .B1(n105892), .B2(n110958), 
        .ZN(n82158) );
  OAI21_X1 U67443 ( .B1(n106777), .B2(n82159), .A(n82160), .ZN(n80122) );
  NAND2_X1 U67444 ( .A1(n82161), .A2(n106777), .ZN(n82160) );
  XNOR2_X1 U67445 ( .A(n82162), .B(n82163), .ZN(n82161) );
  AOI21_X1 U67446 ( .B1(n82151), .B2(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[2] ), .A(n82164), .ZN(n82162) );
  XOR2_X1 U67447 ( .A(n82165), .B(n82163), .Z(n82159) );
  XNOR2_X1 U67448 ( .A(n82166), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [3]), .ZN(n82163) );
  AOI21_X1 U67449 ( .B1(n82151), .B2(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[2] ), .A(n82164), .ZN(n82165) );
  NAND2_X1 U67450 ( .A1(n82167), .A2(n57425), .ZN(n82151) );
  AOI22_X1 U67451 ( .A1(n106818), .A2(n105051), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[19] ), .ZN(n82157) );
  OR2_X1 U67452 ( .A1(n82168), .A2(n82169), .ZN(n60305) );
  AOI22_X1 U67454 ( .A1(n105895), .A2(DataAddr[20]), .B1(n105156), .B2(n110334), .ZN(n82170) );
  NAND2_X1 U67455 ( .A1(n82171), .A2(n82172), .ZN(n82168) );
  AOI22_X1 U67456 ( .A1(n105891), .A2(n110443), .B1(n82173), .B2(n105045), 
        .ZN(n82172) );
  AOI22_X1 U67457 ( .A1(n105158), .A2(\DLX_Datapath/next_A_IDEX[20] ), .B1(
        n82174), .B2(n104706), .ZN(n82171) );
  OR2_X1 U67458 ( .A1(n82175), .A2(n82176), .ZN(n60304) );
  OAI21_X1 U67459 ( .B1(n62204), .B2(n104753), .A(n82177), .ZN(n82176) );
  AOI22_X1 U67460 ( .A1(n105894), .A2(DataAddr[21]), .B1(n105156), .B2(n110336), .ZN(n82177) );
  NAND2_X1 U67461 ( .A1(n82178), .A2(n82179), .ZN(n82175) );
  AOI22_X1 U67462 ( .A1(n105896), .A2(n82180), .B1(n105892), .B2(n110444), 
        .ZN(n82179) );
  AOI22_X1 U67463 ( .A1(n106817), .A2(n105051), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[21] ), .ZN(n82178) );
  AOI22_X1 U67466 ( .A1(n105894), .A2(DataAddr[22]), .B1(n105156), .B2(n110228), .ZN(n82183) );
  AOI22_X1 U67468 ( .A1(n105891), .A2(n110445), .B1(n82186), .B2(n105045), 
        .ZN(n82185) );
  AOI22_X1 U67469 ( .A1(n105158), .A2(\DLX_Datapath/next_A_IDEX[22] ), .B1(
        n105897), .B2(n82187), .ZN(n82184) );
  OR2_X1 U67470 ( .A1(n82188), .A2(n82189), .ZN(n60302) );
  OAI21_X1 U67471 ( .B1(n62191), .B2(n104753), .A(n82190), .ZN(n82189) );
  AOI22_X1 U67472 ( .A1(n105894), .A2(DataAddr[23]), .B1(n105157), .B2(n106824), .ZN(n82190) );
  NAND2_X1 U67473 ( .A1(n82191), .A2(n82192), .ZN(n82188) );
  AOI22_X1 U67474 ( .A1(n105896), .A2(n82193), .B1(n105892), .B2(n110446), 
        .ZN(n82192) );
  AOI22_X1 U67475 ( .A1(n82194), .A2(n105050), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[23] ), .ZN(n82191) );
  OR2_X1 U67476 ( .A1(n82196), .A2(n82195), .ZN(n60301) );
  OAI21_X1 U67477 ( .B1(n59477), .B2(net113091), .A(n82197), .ZN(n82196) );
  AOI22_X1 U67478 ( .A1(n105895), .A2(DataAddr[24]), .B1(n105157), .B2(
        net2410613), .ZN(n82197) );
  NAND2_X1 U67479 ( .A1(n82199), .A2(n82198), .ZN(n82195) );
  AOI22_X1 U67480 ( .A1(n105896), .A2(n80128), .B1(n105891), .B2(n62197), .ZN(
        n82199) );
  OR2_X1 U67482 ( .A1(n82203), .A2(n105020), .ZN(n82202) );
  AOI21_X1 U67483 ( .B1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [0]), 
        .B2(n111133), .A(n82200), .ZN(n82203) );
  AOI22_X1 U67484 ( .A1(n106816), .A2(n105051), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[24] ), .ZN(n82198) );
  OR2_X1 U67485 ( .A1(n82204), .A2(n82205), .ZN(n60300) );
  OAI21_X1 U67486 ( .B1(n57428), .B2(net113081), .A(n82206), .ZN(n82205) );
  AOI22_X1 U67487 ( .A1(n105894), .A2(DataAddr[25]), .B1(n105157), .B2(n108049), .ZN(n82206) );
  NAND2_X1 U67488 ( .A1(n82207), .A2(n82208), .ZN(n82204) );
  AOI22_X1 U67489 ( .A1(n105896), .A2(n104800), .B1(n105891), .B2(net2411291), 
        .ZN(n82208) );
  AOI22_X1 U67492 ( .A1(n82211), .A2(n105889), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[25] ), .ZN(n82207) );
  OR2_X1 U67493 ( .A1(n82212), .A2(n82213), .ZN(n60299) );
  AOI22_X1 U67495 ( .A1(n105895), .A2(DataAddr[26]), .B1(n105156), .B2(n108051), .ZN(n82214) );
  NAND2_X1 U67496 ( .A1(n82216), .A2(n82215), .ZN(n82212) );
  AOI22_X1 U67497 ( .A1(n80148), .A2(n105896), .B1(n105892), .B2(n66263), .ZN(
        n82216) );
  OAI21_X1 U67502 ( .B1(n104797), .B2(n82223), .A(n82224), .ZN(n82217) );
  AOI22_X1 U67503 ( .A1(n106815), .A2(n105051), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[26] ), .ZN(n82215) );
  OR2_X1 U67504 ( .A1(n82225), .A2(n82226), .ZN(n60298) );
  OAI21_X1 U67505 ( .B1(n59478), .B2(net113091), .A(n82227), .ZN(n82226) );
  AOI22_X1 U67506 ( .A1(n105894), .A2(DataAddr[27]), .B1(n105156), .B2(n107747), .ZN(n82227) );
  NAND2_X1 U67507 ( .A1(n82228), .A2(n82229), .ZN(n82225) );
  AOI22_X1 U67508 ( .A1(n105897), .A2(n80106), .B1(n105891), .B2(n62198), .ZN(
        n82229) );
  OAI21_X1 U67509 ( .B1(n105020), .B2(n82230), .A(n82231), .ZN(n80106) );
  NAND2_X1 U67510 ( .A1(n82232), .A2(n105020), .ZN(n82231) );
  XOR2_X1 U67511 ( .A(n82233), .B(n82234), .Z(n82232) );
  NAND2_X1 U67512 ( .A1(n82235), .A2(n82218), .ZN(n82233) );
  OAI21_X1 U67513 ( .B1(n111132), .B2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [2]), .A(n82223), .ZN(
        n82235) );
  OAI21_X1 U67514 ( .B1(n82236), .B2(n82237), .A(n82238), .ZN(n82223) );
  NAND2_X1 U67515 ( .A1(n111133), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [0]), .ZN(n82237) );
  XNOR2_X1 U67516 ( .A(n82239), .B(n82234), .ZN(n82230) );
  XOR2_X1 U67517 ( .A(n111132), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [3]), .Z(n82234) );
  NAND2_X1 U67518 ( .A1(n82240), .A2(n82218), .ZN(n82239) );
  NAND2_X1 U67519 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [2]), 
        .A2(n111132), .ZN(n82218) );
  OAI21_X1 U67520 ( .B1(n111132), .B2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [2]), .A(n82224), .ZN(
        n82240) );
  OAI21_X1 U67521 ( .B1(n82200), .B2(n82236), .A(n82238), .ZN(n82224) );
  NAND2_X1 U67522 ( .A1(n111132), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [1]), .ZN(n82238) );
  NOR2_X1 U67523 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [1]), 
        .A2(n111132), .ZN(n82236) );
  AOI22_X1 U67524 ( .A1(n82241), .A2(n105890), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[27] ), .ZN(n82228) );
  OAI21_X1 U67526 ( .B1(n57426), .B2(n104753), .A(n82244), .ZN(n82243) );
  AOI22_X1 U67527 ( .A1(n82022), .A2(DataAddr[28]), .B1(n105155), .B2(n106827), 
        .ZN(n82244) );
  AOI22_X1 U67529 ( .A1(n105891), .A2(n110964), .B1(n80124), .B2(n105897), 
        .ZN(n82246) );
  AOI22_X1 U67532 ( .A1(n82250), .A2(n105045), .B1(n104699), .B2(
        \DLX_Datapath/next_A_IDEX[28] ), .ZN(n82245) );
  OR2_X1 U67533 ( .A1(n82251), .A2(n82252), .ZN(n60296) );
  OAI21_X1 U67534 ( .B1(n57429), .B2(net113091), .A(n82253), .ZN(n82252) );
  AOI22_X1 U67535 ( .A1(n105894), .A2(DataAddr[29]), .B1(n105157), .B2(n106828), .ZN(n82253) );
  NAND2_X1 U67536 ( .A1(n82255), .A2(n82254), .ZN(n82251) );
  AOI22_X1 U67537 ( .A1(n80150), .A2(n104706), .B1(n105891), .B2(net2411318), 
        .ZN(n82255) );
  AOI21_X1 U67541 ( .B1(n82260), .B2(n105153), .A(n57426), .ZN(n82259) );
  AOI22_X1 U67542 ( .A1(n82261), .A2(n105889), .B1(n105159), .B2(
        \DLX_Datapath/next_A_IDEX[29] ), .ZN(n82254) );
  OAI21_X1 U67544 ( .B1(n57430), .B2(net113091), .A(n82264), .ZN(n82263) );
  AOI22_X1 U67545 ( .A1(n82022), .A2(DataAddr[30]), .B1(n105155), .B2(n106826), 
        .ZN(n82264) );
  AOI22_X1 U67547 ( .A1(n105891), .A2(n110965), .B1(n82267), .B2(n105051), 
        .ZN(n82266) );
  AOI22_X1 U67548 ( .A1(n105026), .A2(n82021), .B1(n105158), .B2(
        \DLX_Datapath/next_A_IDEX[30] ), .ZN(n82265) );
  OAI21_X1 U67551 ( .B1(n57430), .B2(n105153), .A(n82272), .ZN(n82268) );
  AOI22_X1 U67554 ( .A1(n82022), .A2(DataAddr[31]), .B1(n105155), .B2(n106825), 
        .ZN(n82275) );
  AOI21_X1 U67556 ( .B1(n82277), .B2(n82278), .A(n106807), .ZN(n82276) );
  AOI22_X1 U67560 ( .A1(n105891), .A2(n110966), .B1(n82284), .B2(n105890), 
        .ZN(n82283) );
  AOI21_X1 U67564 ( .B1(n82289), .B2(n82290), .A(n82291), .ZN(n82287) );
  AOI22_X1 U67565 ( .A1(n106843), .A2(n104839), .B1(n106844), .B2(n105041), 
        .ZN(n82291) );
  AOI22_X1 U67566 ( .A1(n105158), .A2(\DLX_Datapath/next_A_IDEX[31] ), .B1(
        n80136), .B2(n105896), .ZN(n82282) );
  OAI21_X1 U67567 ( .B1(n82293), .B2(n82294), .A(n82295), .ZN(n80136) );
  OAI21_X1 U67568 ( .B1(n82296), .B2(n82297), .A(n82294), .ZN(n82295) );
  XOR2_X1 U67572 ( .A(n105153), .B(n57431), .Z(n82294) );
  AOI22_X1 U67573 ( .A1(n82298), .A2(n82272), .B1(n105018), .B2(n82299), .ZN(
        n82293) );
  OAI21_X1 U67574 ( .B1(n57430), .B2(n105153), .A(n110963), .ZN(n82299) );
  AOI21_X1 U67575 ( .B1(n57426), .B2(n57429), .A(n105153), .ZN(n82300) );
  NAND2_X1 U67576 ( .A1(n57430), .A2(n105153), .ZN(n82272) );
  NAND2_X1 U67578 ( .A1(n82260), .A2(n82258), .ZN(n82249) );
  OR2_X1 U67579 ( .A1(n82301), .A2(n105153), .ZN(n82258) );
  NOR3_X1 U67582 ( .A1(n57427), .A2(n59478), .A3(n57428), .ZN(n82302) );
  NOR2_X1 U67584 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [0]), 
        .A2(n111133), .ZN(n82200) );
  OAI21_X1 U67592 ( .B1(IR_in[15]), .B2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [3]), .A(n82319), .ZN(
        n82315) );
  NOR2_X1 U67593 ( .A1(n82320), .A2(n82321), .ZN(n82319) );
  OAI21_X1 U67594 ( .B1(n82322), .B2(n82313), .A(n82323), .ZN(n82309) );
  AOI22_X1 U67595 ( .A1(n82324), .A2(n108275), .B1(n62199), .B2(n111155), .ZN(
        n82322) );
  NOR4_X1 U67597 ( .A1(n62182), .A2(n82321), .A3(n111154), .A4(n82317), .ZN(
        n82313) );
  NOR2_X1 U67598 ( .A1(n82311), .A2(n82312), .ZN(n82308) );
  AOI21_X1 U67599 ( .B1(n82325), .B2(n82326), .A(n82321), .ZN(n82312) );
  OAI21_X1 U67600 ( .B1(n82327), .B2(n82328), .A(n82323), .ZN(n82325) );
  AOI22_X1 U67601 ( .A1(n62191), .A2(n82304), .B1(n62196), .B2(n111136), .ZN(
        n82306) );
  AOI21_X1 U67602 ( .B1(IR_in[24]), .B2(n111134), .A(n111135), .ZN(n82303) );
  NAND2_X1 U67603 ( .A1(n105153), .A2(n82329), .ZN(n82271) );
  AOI21_X1 U67604 ( .B1(IR_in[25]), .B2(n111134), .A(n111135), .ZN(n82248) );
  NOR2_X1 U67605 ( .A1(n82330), .A2(n105150), .ZN(n82021) );
  NAND2_X1 U67606 ( .A1(n82280), .A2(n82286), .ZN(n82330) );
  OAI21_X1 U67607 ( .B1(n82331), .B2(n82332), .A(n82333), .ZN(n82286) );
  NAND2_X1 U67608 ( .A1(n82334), .A2(IR_in[27]), .ZN(n82333) );
  NOR3_X1 U67609 ( .A1(n82335), .A2(n82336), .A3(n82337), .ZN(n82331) );
  AOI21_X1 U67610 ( .B1(n82338), .B2(n82339), .A(n82340), .ZN(n82337) );
  AOI22_X1 U67611 ( .A1(n82341), .A2(n111001), .B1(n82342), .B2(n110973), .ZN(
        n82339) );
  AOI22_X1 U67612 ( .A1(n105074), .A2(n110995), .B1(n104835), .B2(n110980), 
        .ZN(n82338) );
  AOI21_X1 U67613 ( .B1(n82344), .B2(n82345), .A(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [0]), .ZN(n82336) );
  NAND2_X1 U67614 ( .A1(n105076), .A2(n82346), .ZN(n82345) );
  NAND2_X1 U67615 ( .A1(n82347), .A2(n82348), .ZN(n82346) );
  AOI22_X1 U67616 ( .A1(n82341), .A2(n110998), .B1(n82342), .B2(n110970), .ZN(
        n82348) );
  AOI22_X1 U67617 ( .A1(n105074), .A2(n110992), .B1(n104835), .B2(n110977), 
        .ZN(n82347) );
  AOI22_X1 U67618 ( .A1(n82349), .A2(n104912), .B1(n105075), .B2(n82350), .ZN(
        n82344) );
  OR2_X1 U67619 ( .A1(n82351), .A2(n82352), .ZN(n82350) );
  AOI21_X1 U67620 ( .B1(n82353), .B2(n82354), .A(PC_out[3]), .ZN(n82352) );
  AOI22_X1 U67621 ( .A1(n82341), .A2(n111009), .B1(n82342), .B2(n110960), .ZN(
        n82354) );
  AOI22_X1 U67622 ( .A1(n105074), .A2(n111002), .B1(n104835), .B2(n110982), 
        .ZN(n82353) );
  AOI21_X1 U67623 ( .B1(n82355), .B2(n82356), .A(n104912), .ZN(n82351) );
  AOI22_X1 U67624 ( .A1(n82341), .A2(n111011), .B1(n82342), .B2(n110961), .ZN(
        n82356) );
  AOI22_X1 U67625 ( .A1(n105074), .A2(n111004), .B1(n104835), .B2(n110984), 
        .ZN(n82355) );
  AOI21_X1 U67626 ( .B1(n82357), .B2(n82358), .A(n105075), .ZN(n82349) );
  AOI22_X1 U67627 ( .A1(n82341), .A2(n110996), .B1(n82342), .B2(n110968), .ZN(
        n82358) );
  AOI22_X1 U67628 ( .A1(n105074), .A2(n110990), .B1(n104835), .B2(n110975), 
        .ZN(n82357) );
  AOI21_X1 U67629 ( .B1(n82359), .B2(n82360), .A(net2465400), .ZN(n82335) );
  NAND2_X1 U67630 ( .A1(n82361), .A2(n104912), .ZN(n82360) );
  AOI21_X1 U67631 ( .B1(n82362), .B2(n82363), .A(n105075), .ZN(n82361) );
  AOI22_X1 U67632 ( .A1(n82341), .A2(n111000), .B1(n82342), .B2(n110972), .ZN(
        n82363) );
  AOI22_X1 U67633 ( .A1(n105074), .A2(n110994), .B1(n104835), .B2(n110979), 
        .ZN(n82362) );
  OAI21_X1 U67634 ( .B1(n82364), .B2(n82365), .A(n105075), .ZN(n82359) );
  AOI21_X1 U67635 ( .B1(n82366), .B2(n82367), .A(PC_out[3]), .ZN(n82365) );
  AOI22_X1 U67636 ( .A1(n82341), .A2(n111013), .B1(n82342), .B2(n110962), .ZN(
        n82367) );
  AOI22_X1 U67637 ( .A1(n105074), .A2(n111006), .B1(n104835), .B2(n110986), 
        .ZN(n82366) );
  AOI21_X1 U67638 ( .B1(n82368), .B2(n82369), .A(n104912), .ZN(n82364) );
  AOI22_X1 U67639 ( .A1(n82341), .A2(n111015), .B1(n82342), .B2(n106812), .ZN(
        n82369) );
  NOR2_X1 U67640 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_0/S_0[1] ), 
        .A2(n105072), .ZN(n82342) );
  NOR2_X1 U67641 ( .A1(PC_out[0]), .A2(n105073), .ZN(n82341) );
  AOI22_X1 U67642 ( .A1(n105074), .A2(n111008), .B1(n104835), .B2(n110988), 
        .ZN(n82368) );
  OAI21_X1 U67646 ( .B1(n104734), .B2(n82023), .A(n82371), .ZN(n60293) );
  NAND2_X1 U67647 ( .A1(n106347), .A2(n108615), .ZN(n82371) );
  XNOR2_X1 U67648 ( .A(PC_out[0]), .B(IR_in[0]), .ZN(n82023) );
  OAI21_X1 U67649 ( .B1(n104735), .B2(n106803), .A(n82372), .ZN(n60292) );
  NAND2_X1 U67650 ( .A1(n106347), .A2(n108616), .ZN(n82372) );
  OAI21_X1 U67651 ( .B1(n104736), .B2(n106802), .A(n82373), .ZN(n60291) );
  NAND2_X1 U67652 ( .A1(n106347), .A2(n108617), .ZN(n82373) );
  OAI21_X1 U67653 ( .B1(n104734), .B2(n106801), .A(n82374), .ZN(n60290) );
  NAND2_X1 U67654 ( .A1(n106347), .A2(n108618), .ZN(n82374) );
  OAI21_X1 U67655 ( .B1(n104734), .B2(n106782), .A(n82375), .ZN(n60273) );
  NAND2_X1 U67656 ( .A1(n106347), .A2(n110443), .ZN(n82375) );
  XOR2_X1 U67657 ( .A(n82376), .B(n82377), .Z(n82174) );
  NAND2_X1 U67658 ( .A1(n82323), .A2(n110441), .ZN(n82376) );
  OAI21_X1 U67659 ( .B1(n106779), .B2(n104734), .A(n82378), .ZN(n60272) );
  NAND2_X1 U67660 ( .A1(n106347), .A2(n110444), .ZN(n82378) );
  OAI21_X1 U67663 ( .B1(n82328), .B2(n106780), .A(n82323), .ZN(n82381) );
  OAI21_X1 U67664 ( .B1(n106778), .B2(n104734), .A(n82382), .ZN(n60271) );
  NAND2_X1 U67665 ( .A1(n106347), .A2(n110445), .ZN(n82382) );
  AOI21_X1 U67667 ( .B1(n82385), .B2(n62196), .A(n82386), .ZN(n82384) );
  NOR3_X1 U67668 ( .A1(n82387), .A2(n62196), .A3(n104794), .ZN(n82386) );
  OAI21_X1 U67671 ( .B1(n106781), .B2(n104737), .A(n82390), .ZN(n60270) );
  NAND2_X1 U67672 ( .A1(n106347), .A2(n110446), .ZN(n82390) );
  OAI21_X1 U67673 ( .B1(n82377), .B2(n82391), .A(n82392), .ZN(n82193) );
  NAND2_X1 U67674 ( .A1(n82393), .A2(n82377), .ZN(n82392) );
  XOR2_X1 U67675 ( .A(n82394), .B(n82395), .Z(n82393) );
  AOI21_X1 U67676 ( .B1(n82388), .B2(n82396), .A(n82311), .ZN(n82395) );
  OAI21_X1 U67677 ( .B1(n82321), .B2(n110441), .A(n82326), .ZN(n82388) );
  NOR2_X1 U67678 ( .A1(n62185), .A2(n82397), .ZN(n82328) );
  XNOR2_X1 U67680 ( .A(n82304), .B(n62191), .ZN(n82394) );
  AOI21_X1 U67681 ( .B1(IR_in[23]), .B2(n111134), .A(n111135), .ZN(n82304) );
  AOI21_X1 U67682 ( .B1(n82389), .B2(n82396), .A(n82311), .ZN(n82398) );
  NOR2_X1 U67683 ( .A1(n62196), .A2(n111136), .ZN(n82311) );
  NAND2_X1 U67684 ( .A1(n62196), .A2(n111136), .ZN(n82396) );
  OAI21_X1 U67685 ( .B1(n111152), .B2(n82399), .A(n82400), .ZN(n82387) );
  OAI21_X1 U67686 ( .B1(n82321), .B2(n110442), .A(n82326), .ZN(n82389) );
  NAND2_X1 U67687 ( .A1(n82380), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [1]), .ZN(n82326) );
  NAND2_X1 U67688 ( .A1(n62185), .A2(n82397), .ZN(n82323) );
  AOI21_X1 U67689 ( .B1(IR_in[20]), .B2(n111134), .A(n111135), .ZN(n82397) );
  NOR2_X1 U67690 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [1]), 
        .A2(n82380), .ZN(n82321) );
  OAI21_X1 U67691 ( .B1(n111153), .B2(n82399), .A(n82400), .ZN(n82380) );
  AOI21_X1 U67692 ( .B1(n82142), .B2(n106823), .A(n82327), .ZN(n82377) );
  OAI21_X1 U67693 ( .B1(n57424), .B2(n82166), .A(n82401), .ZN(n82327) );
  NAND2_X1 U67694 ( .A1(n82402), .A2(n82403), .ZN(n82401) );
  OAI21_X1 U67695 ( .B1(n82404), .B2(n82405), .A(n107745), .ZN(n82402) );
  NOR2_X1 U67696 ( .A1(n57425), .A2(n82167), .ZN(n82164) );
  AOI22_X1 U67697 ( .A1(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[1] ), .A2(n82406), .B1(n111131), .B2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [1]), .ZN(n82404) );
  NAND4_X2 U67698 ( .A1(n82403), .A2(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[1] ), .A3(n82406), .A4(n107746), .ZN(n82317) );
  XNOR2_X1 U67699 ( .A(n82167), .B(n57425), .ZN(n82405) );
  AOI21_X1 U67700 ( .B1(IR_in[18]), .B2(n111134), .A(n111135), .ZN(n82167) );
  XOR2_X1 U67701 ( .A(n82407), .B(n59472), .Z(n82406) );
  NAND2_X1 U67702 ( .A1(n57424), .A2(n82166), .ZN(n82403) );
  AOI21_X1 U67703 ( .B1(IR_in[19]), .B2(n111134), .A(n111135), .ZN(n82166) );
  NAND2_X1 U67705 ( .A1(n82410), .A2(n82409), .ZN(n82408) );
  AOI21_X1 U67706 ( .B1(n82411), .B2(n108275), .A(n82320), .ZN(n82410) );
  OAI21_X1 U67708 ( .B1(IR_in[13]), .B2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [1]), .A(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[1] ), .ZN(n82412) );
  OAI21_X1 U67709 ( .B1(n62199), .B2(n111155), .A(n82413), .ZN(n82318) );
  NAND2_X1 U67710 ( .A1(IR_in[13]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [1]), .ZN(n82413) );
  NOR2_X1 U67711 ( .A1(n104368), .A2(net71745), .ZN(n82411) );
  NAND2_X1 U67719 ( .A1(IR_in[8]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [0]), .ZN(n81255) );
  AOI21_X1 U67726 ( .B1(n82429), .B2(n82428), .A(n104371), .ZN(n82427) );
  NOR2_X1 U67727 ( .A1(n111158), .A2(net2465400), .ZN(n104371) );
  OAI21_X1 U67728 ( .B1(n105075), .B2(n111160), .A(net2465244), .ZN(n82429) );
  AOI21_X1 U67729 ( .B1(n82430), .B2(n111159), .A(n104808), .ZN(n82428) );
  NAND2_X1 U67730 ( .A1(n105071), .A2(PC_out[2]), .ZN(n82430) );
  AOI22_X1 U67731 ( .A1(n82431), .A2(n82432), .B1(IR_in[5]), .B2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [1]), .ZN(n82426) );
  NOR3_X1 U67732 ( .A1(n82077), .A2(n82076), .A3(n104808), .ZN(n82432) );
  NOR2_X1 U67733 ( .A1(n82343), .A2(IR_in[1]), .ZN(n82076) );
  NOR2_X1 U67734 ( .A1(net2465147), .A2(net2465273), .ZN(n82343) );
  NOR2_X1 U67735 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_0/S_0[1] ), 
        .A2(PC_out[0]), .ZN(n82077) );
  OAI21_X1 U67737 ( .B1(n74605), .B2(IR_in[2]), .A(n82433), .ZN(n82075) );
  OAI21_X1 U67738 ( .B1(net67008), .B2(net2465147), .A(net67007), .ZN(n82433)
         );
  NOR2_X1 U67739 ( .A1(n111156), .A2(n104494), .ZN(n104368) );
  AOI22_X1 U67740 ( .A1(n62199), .A2(n111155), .B1(n62182), .B2(n111154), .ZN(
        n82409) );
  AOI22_X1 U67741 ( .A1(n105888), .A2(PC_out[0]), .B1(n105161), .B2(n106765), 
        .ZN(n82434) );
  AOI22_X1 U67742 ( .A1(n105887), .A2(PC_out[1]), .B1(n105161), .B2(n108619), 
        .ZN(n82436) );
  AOI22_X1 U67743 ( .A1(n105887), .A2(n105078), .B1(n105160), .B2(n108621), 
        .ZN(n82437) );
  AOI22_X1 U67744 ( .A1(n105887), .A2(n82043), .B1(n105161), .B2(n108631), 
        .ZN(n82438) );
  XOR2_X1 U67745 ( .A(n105078), .B(n104912), .Z(n82043) );
  AOI22_X1 U67746 ( .A1(n105888), .A2(n82050), .B1(n105160), .B2(n109092), 
        .ZN(n82439) );
  XOR2_X1 U67747 ( .A(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [0]), .B(
        n105076), .Z(n82050) );
  AOI22_X1 U67748 ( .A1(n82435), .A2(n82057), .B1(n105161), .B2(n109094), .ZN(
        n82440) );
  XOR2_X1 U67749 ( .A(n82340), .B(n62201), .Z(n82057) );
  AOI22_X1 U67750 ( .A1(n82435), .A2(n82063), .B1(n105160), .B2(n109096), .ZN(
        n82441) );
  XOR2_X1 U67751 ( .A(n62200), .B(n82442), .Z(n82063) );
  AOI22_X1 U67752 ( .A1(n105888), .A2(n82078), .B1(n105160), .B2(n108972), 
        .ZN(n82443) );
  XOR2_X1 U67753 ( .A(n82444), .B(n62183), .Z(n82078) );
  AOI22_X1 U67754 ( .A1(n82435), .A2(n82085), .B1(n105160), .B2(n109435), .ZN(
        n82445) );
  XOR2_X1 U67755 ( .A(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [0]), .B(
        n82446), .Z(n82085) );
  AOI22_X1 U67756 ( .A1(n105888), .A2(n82092), .B1(n105161), .B2(n109437), 
        .ZN(n82447) );
  XOR2_X1 U67757 ( .A(n82448), .B(n104502), .Z(n82092) );
  AOI22_X1 U67758 ( .A1(n82435), .A2(n104507), .B1(n105161), .B2(n108508), 
        .ZN(n82449) );
  AOI22_X1 U67760 ( .A1(n105887), .A2(n82104), .B1(n105160), .B2(n107621), 
        .ZN(n82451) );
  XOR2_X1 U67761 ( .A(n82452), .B(n104499), .Z(n82104) );
  AOI22_X1 U67762 ( .A1(n105888), .A2(n82112), .B1(n105160), .B2(n108276), 
        .ZN(n82453) );
  AOI21_X1 U67763 ( .B1(n82454), .B2(n104494), .A(n82455), .ZN(n82112) );
  AOI22_X1 U67764 ( .A1(n105887), .A2(n106821), .B1(n105160), .B2(n108278), 
        .ZN(n82456) );
  OAI21_X1 U67765 ( .B1(n82455), .B2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [1]), .A(n82458), .ZN(
        n82457) );
  AOI22_X1 U67766 ( .A1(n105887), .A2(n82123), .B1(n105161), .B2(n108280), 
        .ZN(n82459) );
  AOI21_X1 U67767 ( .B1(n82458), .B2(n62199), .A(n105063), .ZN(n82123) );
  AOI22_X1 U67768 ( .A1(n105888), .A2(n106820), .B1(n105160), .B2(n108158), 
        .ZN(n82461) );
  AOI22_X1 U67770 ( .A1(n82435), .A2(n82136), .B1(n105161), .B2(n109899), .ZN(
        n82464) );
  AOI21_X1 U67771 ( .B1(n82463), .B2(n59471), .A(n82465), .ZN(n82136) );
  AOI22_X1 U67772 ( .A1(n105887), .A2(n106819), .B1(n105160), .B2(n109901), 
        .ZN(n82466) );
  AOI22_X1 U67774 ( .A1(n105888), .A2(n82153), .B1(n105161), .B2(n109783), 
        .ZN(n82469) );
  AOI21_X1 U67775 ( .B1(n82468), .B2(n57425), .A(n105033), .ZN(n82153) );
  AOI22_X1 U67776 ( .A1(n105887), .A2(n106818), .B1(n105160), .B2(n106822), 
        .ZN(n82471) );
  AOI22_X1 U67778 ( .A1(n105888), .A2(n82173), .B1(n105161), .B2(n110334), 
        .ZN(n82474) );
  AOI21_X1 U67779 ( .B1(n82473), .B2(n62185), .A(n82475), .ZN(n82173) );
  AOI22_X1 U67780 ( .A1(n82435), .A2(n106817), .B1(n105161), .B2(n110336), 
        .ZN(n82476) );
  AOI22_X1 U67782 ( .A1(n82435), .A2(n82186), .B1(n105160), .B2(n110228), .ZN(
        n82479) );
  XOR2_X1 U67783 ( .A(n62196), .B(n82478), .Z(n82186) );
  AOI22_X1 U67784 ( .A1(n82435), .A2(n82194), .B1(n105161), .B2(n106824), .ZN(
        n82480) );
  AOI21_X1 U67785 ( .B1(n82481), .B2(n62191), .A(n82482), .ZN(n82194) );
  OR2_X1 U67786 ( .A1(n62196), .A2(n82478), .ZN(n82481) );
  AOI22_X1 U67787 ( .A1(n105888), .A2(n106816), .B1(n105160), .B2(net2410613), 
        .ZN(n82483) );
  OAI21_X1 U67788 ( .B1(n82482), .B2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [0]), .A(n82485), .ZN(
        n82484) );
  AOI22_X1 U67789 ( .A1(n105887), .A2(n82211), .B1(n105161), .B2(n108049), 
        .ZN(n82486) );
  AOI21_X1 U67790 ( .B1(n82485), .B2(n57428), .A(n82487), .ZN(n82211) );
  AOI22_X1 U67791 ( .A1(n105887), .A2(n106815), .B1(n105160), .B2(n108051), 
        .ZN(n82488) );
  AOI22_X1 U67793 ( .A1(n105888), .A2(n82241), .B1(n105161), .B2(n107747), 
        .ZN(n82491) );
  AOI22_X1 U67795 ( .A1(n82435), .A2(n82250), .B1(n105160), .B2(n106827), .ZN(
        n82493) );
  XOR2_X1 U67796 ( .A(n105088), .B(n57426), .Z(n82250) );
  AOI22_X1 U67797 ( .A1(n82435), .A2(n82261), .B1(n105161), .B2(n106828), .ZN(
        n82494) );
  NOR2_X1 U67798 ( .A1(n106814), .A2(n82495), .ZN(n82261) );
  OAI21_X1 U67799 ( .B1(n57426), .B2(n105088), .A(n57429), .ZN(n82496) );
  AOI22_X1 U67800 ( .A1(n105888), .A2(n82267), .B1(n105160), .B2(n106826), 
        .ZN(n82497) );
  XOR2_X1 U67801 ( .A(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0 [2]), .B(
        n82495), .Z(n82267) );
  AOI22_X1 U67802 ( .A1(n105887), .A2(n82284), .B1(n105161), .B2(n106825), 
        .ZN(n82498) );
  NOR2_X1 U67805 ( .A1(n82490), .A2(n105068), .ZN(n82495) );
  NAND2_X1 U67807 ( .A1(n82487), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [2]), .ZN(n82490) );
  NOR2_X1 U67808 ( .A1(n82485), .A2(n57428), .ZN(n82487) );
  NOR2_X1 U67810 ( .A1(n82500), .A2(n82478), .ZN(n82482) );
  NAND2_X1 U67811 ( .A1(n82475), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [1]), .ZN(n82478) );
  NAND2_X1 U67813 ( .A1(n105033), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [3]), .ZN(n82473) );
  NAND2_X1 U67815 ( .A1(n82465), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [1]), .ZN(n82468) );
  NAND2_X1 U67817 ( .A1(n105063), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [3]), .ZN(n82463) );
  NOR2_X1 U67820 ( .A1(n82454), .A2(n104494), .ZN(n82455) );
  OR2_X1 U67821 ( .A1(n82452), .A2(n104499), .ZN(n82454) );
  NOR2_X1 U67823 ( .A1(n82448), .A2(n104502), .ZN(n82450) );
  NAND2_X1 U67824 ( .A1(n82446), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [0]), .ZN(n82448) );
  NOR2_X1 U67825 ( .A1(n82444), .A2(n62183), .ZN(n82446) );
  OR2_X1 U67826 ( .A1(n82442), .A2(n62200), .ZN(n82444) );
  OR2_X1 U67827 ( .A1(n82340), .A2(n62201), .ZN(n82442) );
  NAND2_X1 U67828 ( .A1(n105032), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [0]), .ZN(n82340) );
  AOI21_X1 U67834 ( .B1(n111147), .B2(n82334), .A(n80086), .ZN(n81922) );
  OAI21_X1 U67835 ( .B1(n105072), .B2(n104736), .A(n82502), .ZN(n60229) );
  NAND2_X1 U67836 ( .A1(n106347), .A2(n106809), .ZN(n82502) );
  OAI21_X1 U67837 ( .B1(n105073), .B2(n104734), .A(n82503), .ZN(n60228) );
  NAND2_X1 U67838 ( .A1(n106347), .A2(n110967), .ZN(n82503) );
  OAI21_X1 U67839 ( .B1(n105078), .B2(n104736), .A(n82504), .ZN(n60227) );
  NAND2_X1 U67840 ( .A1(n106347), .A2(n110959), .ZN(n82504) );
  OAI21_X1 U67841 ( .B1(n104912), .B2(n104734), .A(n82505), .ZN(n60226) );
  NAND2_X1 U67842 ( .A1(n106347), .A2(n108971), .ZN(n82505) );
  OAI21_X1 U67843 ( .B1(net2465400), .B2(n104737), .A(n82506), .ZN(n60225) );
  NAND2_X1 U67844 ( .A1(n106347), .A2(n109317), .ZN(n82506) );
  OAI21_X1 U67846 ( .B1(n111130), .B2(n104920), .A(net113153), .ZN(n80104) );
  OAI21_X1 U67847 ( .B1(n82507), .B2(n82508), .A(n82509), .ZN(n60224) );
  OAI21_X1 U67848 ( .B1(n82510), .B2(n82507), .A(n111045), .ZN(n82509) );
  OAI21_X1 U67849 ( .B1(n82507), .B2(n82511), .A(n82512), .ZN(n60223) );
  OAI21_X1 U67850 ( .B1(n82513), .B2(n82507), .A(n110995), .ZN(n82512) );
  OAI21_X1 U67851 ( .B1(n82508), .B2(n82514), .A(n82515), .ZN(n60222) );
  OAI21_X1 U67852 ( .B1(n82510), .B2(n82514), .A(n111046), .ZN(n82515) );
  OAI21_X1 U67853 ( .B1(n82511), .B2(n82514), .A(n82516), .ZN(n60221) );
  OAI21_X1 U67854 ( .B1(n82513), .B2(n82514), .A(n111001), .ZN(n82516) );
  OAI21_X1 U67855 ( .B1(n82508), .B2(n82517), .A(n82518), .ZN(n60220) );
  OAI21_X1 U67856 ( .B1(n82510), .B2(n82517), .A(n111047), .ZN(n82518) );
  OAI21_X1 U67857 ( .B1(n82511), .B2(n82517), .A(n82519), .ZN(n60219) );
  OAI21_X1 U67858 ( .B1(n82513), .B2(n82517), .A(n110973), .ZN(n82519) );
  OAI21_X1 U67859 ( .B1(n82508), .B2(n82520), .A(n82521), .ZN(n60218) );
  OAI21_X1 U67860 ( .B1(n82510), .B2(n82520), .A(n111048), .ZN(n82521) );
  OAI21_X1 U67861 ( .B1(n82511), .B2(n82520), .A(n82522), .ZN(n60217) );
  OAI21_X1 U67862 ( .B1(n82513), .B2(n82520), .A(n110980), .ZN(n82522) );
  OAI21_X1 U67863 ( .B1(n82508), .B2(n82523), .A(n82524), .ZN(n60216) );
  OAI21_X1 U67864 ( .B1(n82510), .B2(n82523), .A(n111007), .ZN(n82524) );
  OAI21_X1 U67865 ( .B1(n82511), .B2(n82523), .A(n82525), .ZN(n60215) );
  OAI21_X1 U67866 ( .B1(n82513), .B2(n82523), .A(n111008), .ZN(n82525) );
  OAI21_X1 U67867 ( .B1(n82508), .B2(n82526), .A(n82527), .ZN(n60214) );
  OAI21_X1 U67868 ( .B1(n82510), .B2(n82526), .A(n111014), .ZN(n82527) );
  OAI21_X1 U67869 ( .B1(n82511), .B2(n82526), .A(n82528), .ZN(n60213) );
  OAI21_X1 U67870 ( .B1(n82513), .B2(n82526), .A(n111015), .ZN(n82528) );
  OAI21_X1 U67871 ( .B1(n82508), .B2(n82529), .A(n82530), .ZN(n60212) );
  OAI21_X1 U67872 ( .B1(n82510), .B2(n82529), .A(n107150), .ZN(n82530) );
  OAI21_X1 U67873 ( .B1(n82511), .B2(n82529), .A(n82531), .ZN(n60211) );
  OAI21_X1 U67874 ( .B1(n82513), .B2(n82529), .A(n106812), .ZN(n82531) );
  OAI21_X1 U67875 ( .B1(n82508), .B2(n82532), .A(n82533), .ZN(n60210) );
  OAI21_X1 U67876 ( .B1(n82510), .B2(n82532), .A(n110987), .ZN(n82533) );
  NAND2_X1 U67877 ( .A1(n82534), .A2(n105148), .ZN(n82510) );
  NAND2_X1 U67878 ( .A1(n106552), .A2(n105148), .ZN(n82508) );
  OAI21_X1 U67879 ( .B1(n82511), .B2(n82532), .A(n82536), .ZN(n60209) );
  OAI21_X1 U67880 ( .B1(n82513), .B2(n82532), .A(n110988), .ZN(n82536) );
  NAND2_X1 U67881 ( .A1(n82537), .A2(n105148), .ZN(n82513) );
  NAND2_X1 U67882 ( .A1(n106551), .A2(n105147), .ZN(n82511) );
  OAI21_X1 U67883 ( .B1(n82507), .B2(n82538), .A(n82539), .ZN(n60208) );
  OAI21_X1 U67884 ( .B1(n82507), .B2(n82540), .A(n110993), .ZN(n82539) );
  OAI21_X1 U67885 ( .B1(n82507), .B2(n82541), .A(n82542), .ZN(n60207) );
  OAI21_X1 U67886 ( .B1(n82507), .B2(n82543), .A(n110994), .ZN(n82542) );
  OAI21_X1 U67887 ( .B1(n82514), .B2(n82538), .A(n82544), .ZN(n60206) );
  OAI21_X1 U67888 ( .B1(n82514), .B2(n82540), .A(n110999), .ZN(n82544) );
  OAI21_X1 U67889 ( .B1(n82514), .B2(n82541), .A(n82545), .ZN(n60205) );
  OAI21_X1 U67890 ( .B1(n82514), .B2(n82543), .A(n111000), .ZN(n82545) );
  OAI21_X1 U67891 ( .B1(n82517), .B2(n82538), .A(n82546), .ZN(n60204) );
  OAI21_X1 U67892 ( .B1(n82517), .B2(n82540), .A(n110971), .ZN(n82546) );
  OAI21_X1 U67893 ( .B1(n82517), .B2(n82541), .A(n82547), .ZN(n60203) );
  OAI21_X1 U67894 ( .B1(n82517), .B2(n82543), .A(n110972), .ZN(n82547) );
  OAI21_X1 U67895 ( .B1(n82520), .B2(n82538), .A(n82548), .ZN(n60202) );
  OAI21_X1 U67896 ( .B1(n82520), .B2(n82540), .A(n110978), .ZN(n82548) );
  OAI21_X1 U67897 ( .B1(n82520), .B2(n82541), .A(n82549), .ZN(n60201) );
  OAI21_X1 U67898 ( .B1(n82520), .B2(n82543), .A(n110979), .ZN(n82549) );
  OAI21_X1 U67899 ( .B1(n82523), .B2(n82538), .A(n82550), .ZN(n60200) );
  OAI21_X1 U67900 ( .B1(n82523), .B2(n82540), .A(n111005), .ZN(n82550) );
  OAI21_X1 U67901 ( .B1(n82523), .B2(n82541), .A(n82551), .ZN(n60199) );
  OAI21_X1 U67902 ( .B1(n82523), .B2(n82543), .A(n111006), .ZN(n82551) );
  OAI21_X1 U67903 ( .B1(n82526), .B2(n82538), .A(n82552), .ZN(n60198) );
  OAI21_X1 U67904 ( .B1(n82526), .B2(n82540), .A(n111012), .ZN(n82552) );
  OAI21_X1 U67905 ( .B1(n82526), .B2(n82541), .A(n82553), .ZN(n60197) );
  OAI21_X1 U67906 ( .B1(n82526), .B2(n82543), .A(n111013), .ZN(n82553) );
  OAI21_X1 U67907 ( .B1(n82529), .B2(n82538), .A(n82554), .ZN(n60196) );
  OAI21_X1 U67908 ( .B1(n82529), .B2(n82540), .A(n109320), .ZN(n82554) );
  OAI21_X1 U67909 ( .B1(n82529), .B2(n82541), .A(n82555), .ZN(n60195) );
  OAI21_X1 U67910 ( .B1(n82529), .B2(n82543), .A(n110962), .ZN(n82555) );
  OAI21_X1 U67911 ( .B1(n82532), .B2(n82538), .A(n82556), .ZN(n60194) );
  OAI21_X1 U67912 ( .B1(n82532), .B2(n82540), .A(n110985), .ZN(n82556) );
  NAND2_X1 U67913 ( .A1(n82534), .A2(n82557), .ZN(n82540) );
  NAND2_X1 U67914 ( .A1(n106552), .A2(n82557), .ZN(n82538) );
  OAI21_X1 U67915 ( .B1(n82532), .B2(n82541), .A(n82558), .ZN(n60193) );
  OAI21_X1 U67916 ( .B1(n82532), .B2(n82543), .A(n110986), .ZN(n82558) );
  NAND2_X1 U67917 ( .A1(n82537), .A2(n82557), .ZN(n82543) );
  NAND2_X1 U67918 ( .A1(n106551), .A2(n105149), .ZN(n82541) );
  OAI21_X1 U67919 ( .B1(n82507), .B2(n82559), .A(n82560), .ZN(n60192) );
  OAI21_X1 U67920 ( .B1(n82507), .B2(n82561), .A(n110991), .ZN(n82560) );
  OAI21_X1 U67921 ( .B1(n82507), .B2(n82562), .A(n82563), .ZN(n60191) );
  OAI21_X1 U67922 ( .B1(n82507), .B2(n82564), .A(n110992), .ZN(n82563) );
  OAI21_X1 U67923 ( .B1(n82514), .B2(n82559), .A(n82565), .ZN(n60190) );
  OAI21_X1 U67924 ( .B1(n82514), .B2(n82561), .A(n110997), .ZN(n82565) );
  OAI21_X1 U67925 ( .B1(n82514), .B2(n82562), .A(n82566), .ZN(n60189) );
  OAI21_X1 U67926 ( .B1(n82514), .B2(n82564), .A(n110998), .ZN(n82566) );
  OAI21_X1 U67927 ( .B1(n82517), .B2(n82559), .A(n82567), .ZN(n60188) );
  OAI21_X1 U67928 ( .B1(n82517), .B2(n82561), .A(n110969), .ZN(n82567) );
  OAI21_X1 U67929 ( .B1(n82517), .B2(n82562), .A(n82568), .ZN(n60187) );
  OAI21_X1 U67930 ( .B1(n82517), .B2(n82564), .A(n110970), .ZN(n82568) );
  OAI21_X1 U67931 ( .B1(n82520), .B2(n82559), .A(n82569), .ZN(n60186) );
  OAI21_X1 U67932 ( .B1(n82520), .B2(n82561), .A(n110976), .ZN(n82569) );
  OAI21_X1 U67933 ( .B1(n82520), .B2(n82562), .A(n82570), .ZN(n60185) );
  OAI21_X1 U67934 ( .B1(n82520), .B2(n82564), .A(n110977), .ZN(n82570) );
  OAI21_X1 U67935 ( .B1(n82523), .B2(n82559), .A(n82571), .ZN(n60184) );
  OAI21_X1 U67936 ( .B1(n82523), .B2(n82561), .A(n111003), .ZN(n82571) );
  OAI21_X1 U67937 ( .B1(n82523), .B2(n82562), .A(n82572), .ZN(n60183) );
  OAI21_X1 U67938 ( .B1(n82523), .B2(n82564), .A(n111004), .ZN(n82572) );
  OAI21_X1 U67939 ( .B1(n82526), .B2(n82559), .A(n82573), .ZN(n60182) );
  OAI21_X1 U67940 ( .B1(n82526), .B2(n82561), .A(n111010), .ZN(n82573) );
  OAI21_X1 U67941 ( .B1(n82526), .B2(n82562), .A(n82574), .ZN(n60181) );
  OAI21_X1 U67942 ( .B1(n82526), .B2(n82564), .A(n111011), .ZN(n82574) );
  OAI21_X1 U67943 ( .B1(n82529), .B2(n82559), .A(n82575), .ZN(n60180) );
  OAI21_X1 U67944 ( .B1(n82529), .B2(n82561), .A(n109318), .ZN(n82575) );
  OAI21_X1 U67945 ( .B1(n82529), .B2(n82562), .A(n82576), .ZN(n60179) );
  OAI21_X1 U67946 ( .B1(n82529), .B2(n82564), .A(n110961), .ZN(n82576) );
  OAI21_X1 U67947 ( .B1(n82532), .B2(n82559), .A(n82577), .ZN(n60178) );
  OAI21_X1 U67948 ( .B1(n82532), .B2(n82561), .A(n110983), .ZN(n82577) );
  NAND2_X1 U67949 ( .A1(n82534), .A2(n82578), .ZN(n82561) );
  NAND2_X1 U67950 ( .A1(n106552), .A2(n105145), .ZN(n82559) );
  OAI21_X1 U67951 ( .B1(n82532), .B2(n82562), .A(n82579), .ZN(n60177) );
  OAI21_X1 U67952 ( .B1(n82532), .B2(n82564), .A(n110984), .ZN(n82579) );
  NAND2_X1 U67953 ( .A1(n82537), .A2(n82578), .ZN(n82564) );
  NAND2_X1 U67954 ( .A1(n106551), .A2(n105145), .ZN(n82562) );
  OAI21_X1 U67955 ( .B1(n82507), .B2(n82580), .A(n82581), .ZN(n60176) );
  OAI21_X1 U67956 ( .B1(n82507), .B2(n82582), .A(n110989), .ZN(n82581) );
  OAI21_X1 U67957 ( .B1(n82507), .B2(n82583), .A(n82584), .ZN(n60175) );
  OAI21_X1 U67958 ( .B1(n82507), .B2(n82585), .A(n110990), .ZN(n82584) );
  NAND2_X1 U67959 ( .A1(n106808), .A2(n110959), .ZN(n82507) );
  OAI21_X1 U67960 ( .B1(n82514), .B2(n82580), .A(n82586), .ZN(n60174) );
  OAI21_X1 U67961 ( .B1(n82514), .B2(n82582), .A(n111041), .ZN(n82586) );
  OAI21_X1 U67962 ( .B1(n82514), .B2(n82583), .A(n82587), .ZN(n60173) );
  OAI21_X1 U67963 ( .B1(n82514), .B2(n82585), .A(n110996), .ZN(n82587) );
  NAND2_X1 U67964 ( .A1(n106810), .A2(n110959), .ZN(n82514) );
  OAI21_X1 U67965 ( .B1(n82517), .B2(n82580), .A(n82588), .ZN(n60172) );
  OAI21_X1 U67966 ( .B1(n82517), .B2(n82582), .A(n111042), .ZN(n82588) );
  OAI21_X1 U67967 ( .B1(n82517), .B2(n82583), .A(n82589), .ZN(n60171) );
  OAI21_X1 U67968 ( .B1(n82517), .B2(n82585), .A(n110968), .ZN(n82589) );
  NAND2_X1 U67969 ( .A1(n106804), .A2(n110959), .ZN(n82517) );
  OAI21_X1 U67970 ( .B1(n82520), .B2(n82580), .A(n82590), .ZN(n60170) );
  OAI21_X1 U67971 ( .B1(n82520), .B2(n82582), .A(n110974), .ZN(n82590) );
  OAI21_X1 U67972 ( .B1(n82520), .B2(n82583), .A(n82591), .ZN(n60169) );
  OAI21_X1 U67973 ( .B1(n82520), .B2(n82585), .A(n110975), .ZN(n82591) );
  NAND2_X1 U67974 ( .A1(n106811), .A2(n110959), .ZN(n82520) );
  OAI21_X1 U67975 ( .B1(n82523), .B2(n82580), .A(n82592), .ZN(n60168) );
  OAI21_X1 U67976 ( .B1(n82523), .B2(n82582), .A(n111043), .ZN(n82592) );
  OAI21_X1 U67977 ( .B1(n82523), .B2(n82583), .A(n82593), .ZN(n60167) );
  OAI21_X1 U67978 ( .B1(n82523), .B2(n82585), .A(n111002), .ZN(n82593) );
  NAND2_X1 U67979 ( .A1(n61666), .A2(n106808), .ZN(n82523) );
  OAI21_X1 U67980 ( .B1(n82526), .B2(n82580), .A(n82595), .ZN(n60166) );
  OAI21_X1 U67981 ( .B1(n82526), .B2(n82582), .A(n111044), .ZN(n82595) );
  OAI21_X1 U67982 ( .B1(n82526), .B2(n82583), .A(n82596), .ZN(n60165) );
  OAI21_X1 U67983 ( .B1(n82526), .B2(n82585), .A(n111009), .ZN(n82596) );
  NAND2_X1 U67984 ( .A1(n61666), .A2(n106810), .ZN(n82526) );
  OAI21_X1 U67985 ( .B1(n82529), .B2(n82580), .A(n82598), .ZN(n60164) );
  OAI21_X1 U67986 ( .B1(n82529), .B2(n82582), .A(n109319), .ZN(n82598) );
  OAI21_X1 U67987 ( .B1(n82529), .B2(n82583), .A(n82599), .ZN(n60163) );
  OAI21_X1 U67988 ( .B1(n82529), .B2(n82585), .A(n110960), .ZN(n82599) );
  NAND2_X1 U67989 ( .A1(n61666), .A2(n106804), .ZN(n82529) );
  OAI21_X1 U67990 ( .B1(n82532), .B2(n82580), .A(n82601), .ZN(n60162) );
  OAI21_X1 U67991 ( .B1(n82532), .B2(n82582), .A(n110981), .ZN(n82601) );
  NAND2_X1 U67992 ( .A1(n82534), .A2(n105146), .ZN(n82582) );
  NOR2_X1 U67993 ( .A1(n82603), .A2(n82289), .ZN(n82534) );
  NAND2_X1 U67994 ( .A1(n106552), .A2(n82602), .ZN(n82580) );
  OAI21_X1 U67995 ( .B1(n82605), .B2(n82606), .A(n82607), .ZN(n82604) );
  NAND2_X1 U67996 ( .A1(n82608), .A2(n82609), .ZN(n82607) );
  AOI22_X1 U67997 ( .A1(n104907), .A2(n82608), .B1(n104821), .B2(n82609), .ZN(
        n82606) );
  OAI21_X1 U67998 ( .B1(n82532), .B2(n82583), .A(n82610), .ZN(n60161) );
  OAI21_X1 U67999 ( .B1(n82532), .B2(n82585), .A(n110982), .ZN(n82610) );
  NAND2_X1 U68000 ( .A1(n82537), .A2(n82602), .ZN(n82585) );
  OAI21_X1 U68002 ( .B1(n106844), .B2(n106843), .A(net113081), .ZN(n82603) );
  AOI22_X1 U68003 ( .A1(n106553), .A2(n105023), .B1(n106550), .B2(n82613), 
        .ZN(n82611) );
  NAND2_X1 U68004 ( .A1(n106551), .A2(n82602), .ZN(n82583) );
  OAI21_X1 U68005 ( .B1(n82605), .B2(n106806), .A(n82615), .ZN(n82614) );
  AOI22_X1 U68006 ( .A1(n82608), .A2(n104839), .B1(n105041), .B2(n82609), .ZN(
        n82615) );
  NAND2_X1 U68009 ( .A1(n61666), .A2(n106811), .ZN(n82532) );
  NOR4_X1 U68010 ( .A1(n106369), .A2(n106368), .A3(n105123), .A4(n82617), .ZN(
        n60158) );
  OAI21_X1 U68011 ( .B1(n107130), .B2(n81923), .A(n82618), .ZN(n59220) );
  OR2_X1 U68012 ( .A1(n105898), .A2(n100633), .ZN(n82618) );
  OAI21_X1 U68013 ( .B1(n104501), .B2(n81923), .A(n82619), .ZN(n59219) );
  OR2_X1 U68014 ( .A1(n81925), .A2(n100634), .ZN(n82619) );
  OAI21_X1 U68015 ( .B1(n57382), .B2(n81923), .A(n82620), .ZN(n59218) );
  OR2_X1 U68016 ( .A1(n81925), .A2(n100635), .ZN(n82620) );
  OAI21_X1 U68017 ( .B1(n57381), .B2(n81923), .A(n82621), .ZN(n59217) );
  OR2_X1 U68018 ( .A1(n81925), .A2(n100636), .ZN(n82621) );
  OAI21_X1 U68019 ( .B1(n57380), .B2(n81923), .A(n82622), .ZN(n59216) );
  OR2_X1 U68020 ( .A1(n105898), .A2(n100637), .ZN(n82622) );
  NAND2_X1 U68021 ( .A1(net113153), .A2(n107416), .ZN(n81925) );
  NAND2_X1 U68022 ( .A1(n82623), .A2(n61540), .ZN(n81923) );
  NOR2_X1 U68023 ( .A1(n100767), .A2(net113154), .ZN(n82623) );
  OAI21_X1 U68024 ( .B1(n82624), .B2(n82625), .A(n82626), .ZN(n59098) );
  NAND2_X1 U68025 ( .A1(n100767), .A2(net113155), .ZN(n82626) );
  NAND2_X1 U68026 ( .A1(n111147), .A2(n105163), .ZN(n82625) );
  OAI21_X1 U68027 ( .B1(n57390), .B2(n104753), .A(n106596), .ZN(n59093) );
  NOR4_X1 U68028 ( .A1(IR_in[30]), .A2(n82628), .A3(n105152), .A4(n82629), 
        .ZN(n82627) );
  OAI21_X1 U68029 ( .B1(n82630), .B2(n105152), .A(n82631), .ZN(n59090) );
  NAND2_X1 U68030 ( .A1(net113157), .A2(\DLX_ControlUnit/ALUop2 [2]), .ZN(
        n82631) );
  NOR4_X1 U68031 ( .A1(n82632), .A2(n82633), .A3(n111127), .A4(n82634), .ZN(
        n82630) );
  NOR4_X1 U68032 ( .A1(IR_in[4]), .A2(n82635), .A3(n82636), .A4(n81967), .ZN(
        n82634) );
  AOI21_X1 U68033 ( .B1(n111160), .B2(n111159), .A(n82015), .ZN(n82635) );
  OAI21_X1 U68034 ( .B1(net67007), .B2(n111161), .A(n81965), .ZN(n82015) );
  NAND2_X1 U68035 ( .A1(IR_in[2]), .A2(net67008), .ZN(n81965) );
  OAI21_X1 U68036 ( .B1(n111158), .B2(n82007), .A(n82637), .ZN(n82633) );
  OAI21_X1 U68037 ( .B1(n82638), .B2(n111128), .A(n82639), .ZN(n82637) );
  NOR3_X1 U68038 ( .A1(n111123), .A2(IR_in[30]), .A3(IR_in[28]), .ZN(n82638)
         );
  NAND2_X1 U68039 ( .A1(n82640), .A2(n111138), .ZN(n82007) );
  NAND2_X1 U68040 ( .A1(n81998), .A2(n111139), .ZN(n81977) );
  NAND2_X1 U68041 ( .A1(n82641), .A2(n82642), .ZN(n82636) );
  NOR3_X1 U68042 ( .A1(IR_in[7]), .A2(IR_in[9]), .A3(IR_in[8]), .ZN(n82642) );
  NOR2_X1 U68043 ( .A1(IR_in[10]), .A2(n80100), .ZN(n82641) );
  NOR2_X1 U68044 ( .A1(n81967), .A2(n111159), .ZN(n81998) );
  NOR2_X1 U68046 ( .A1(IR_in[0]), .A2(n111161), .ZN(n82640) );
  NOR2_X1 U68047 ( .A1(net67008), .A2(IR_in[2]), .ZN(n81962) );
  OR2_X1 U68048 ( .A1(n82643), .A2(n111121), .ZN(n82632) );
  OAI21_X1 U68050 ( .B1(n80039), .B2(n82646), .A(n82647), .ZN(n82643) );
  OAI21_X1 U68051 ( .B1(n82648), .B2(n105152), .A(n82649), .ZN(n59088) );
  NAND2_X1 U68052 ( .A1(n61670), .A2(net113159), .ZN(n82649) );
  NOR4_X1 U68053 ( .A1(n82650), .A2(n80071), .A3(n80056), .A4(n82006), .ZN(
        n82648) );
  OAI21_X1 U68054 ( .B1(IR_in[26]), .B2(n81976), .A(n82647), .ZN(n82650) );
  OAI21_X1 U68055 ( .B1(n104753), .B2(n107416), .A(n104781), .ZN(n59085) );
  OAI21_X1 U68056 ( .B1(n57393), .B2(net113081), .A(n104781), .ZN(n59084) );
  OAI21_X1 U68057 ( .B1(n80056), .B2(n111118), .A(n105165), .ZN(n81878) );
  NOR3_X1 U68058 ( .A1(n80092), .A2(n111128), .A3(n80071), .ZN(n80099) );
  NAND2_X1 U68059 ( .A1(n111129), .A2(IR_in[28]), .ZN(n82624) );
  OAI21_X1 U68060 ( .B1(n82651), .B2(n105150), .A(n82652), .ZN(n59082) );
  NAND2_X1 U68061 ( .A1(n100496), .A2(net113156), .ZN(n82652) );
  NAND2_X1 U68062 ( .A1(n81921), .A2(net113153), .ZN(n80041) );
  NOR2_X1 U68063 ( .A1(n82654), .A2(n82653), .ZN(n81921) );
  AOI21_X1 U68064 ( .B1(n106769), .B2(n82655), .A(n82277), .ZN(n82654) );
  NAND2_X1 U68065 ( .A1(n82656), .A2(n106942), .ZN(n82277) );
  OAI21_X1 U68066 ( .B1(n105065), .B2(n82290), .A(n82657), .ZN(n82612) );
  AOI22_X1 U68069 ( .A1(n82605), .A2(n105065), .B1(n106806), .B2(n105041), 
        .ZN(n82655) );
  AOI21_X1 U68070 ( .B1(n104910), .B2(n82660), .A(n82278), .ZN(n82653) );
  NAND2_X1 U68071 ( .A1(n82656), .A2(n69325), .ZN(n82278) );
  NAND2_X1 U68073 ( .A1(n82662), .A2(n106770), .ZN(n82661) );
  NOR2_X1 U68074 ( .A1(n106807), .A2(n106805), .ZN(n82662) );
  NAND2_X1 U68075 ( .A1(n106807), .A2(n106805), .ZN(n82290) );
  AOI22_X1 U68076 ( .A1(n82605), .A2(n105041), .B1(n106806), .B2(n105065), 
        .ZN(n82660) );
  NAND2_X1 U68077 ( .A1(n106807), .A2(n82659), .ZN(n82289) );
  OAI21_X1 U68078 ( .B1(n82663), .B2(n82281), .A(n82664), .ZN(n82292) );
  NOR4_X1 U68080 ( .A1(n82666), .A2(n82667), .A3(n82668), .A4(n82669), .ZN(
        n82665) );
  NAND2_X1 U68081 ( .A1(n82670), .A2(n82671), .ZN(n82669) );
  NOR4_X1 U68082 ( .A1(DataAddr[26]), .A2(DataAddr[27]), .A3(DataAddr[30]), 
        .A4(DataAddr[31]), .ZN(n82671) );
  NOR4_X1 U68083 ( .A1(DataAddr[28]), .A2(DataAddr[12]), .A3(DataAddr[29]), 
        .A4(DataAddr[0]), .ZN(n82670) );
  NAND2_X1 U68084 ( .A1(n82672), .A2(n82673), .ZN(n82668) );
  NOR4_X1 U68085 ( .A1(DataAddr[3]), .A2(DataAddr[10]), .A3(DataAddr[11]), 
        .A4(DataAddr[13]), .ZN(n82673) );
  NOR4_X1 U68086 ( .A1(DataAddr[14]), .A2(DataAddr[15]), .A3(DataAddr[24]), 
        .A4(DataAddr[25]), .ZN(n82672) );
  NAND2_X1 U68087 ( .A1(n82674), .A2(n82675), .ZN(n82667) );
  NOR4_X1 U68088 ( .A1(DataAddr[8]), .A2(DataAddr[9]), .A3(DataAddr[5]), .A4(
        DataAddr[4]), .ZN(n82675) );
  NOR4_X1 U68089 ( .A1(DataAddr[6]), .A2(DataAddr[7]), .A3(DataAddr[2]), .A4(
        DataAddr[1]), .ZN(n82674) );
  NAND2_X1 U68090 ( .A1(n82676), .A2(n82677), .ZN(n82666) );
  NOR4_X1 U68091 ( .A1(DataAddr[20]), .A2(DataAddr[21]), .A3(DataAddr[22]), 
        .A4(DataAddr[23]), .ZN(n82677) );
  NOR4_X1 U68092 ( .A1(DataAddr[16]), .A2(DataAddr[17]), .A3(DataAddr[18]), 
        .A4(DataAddr[19]), .ZN(n82676) );
  OAI21_X1 U68093 ( .B1(n82678), .B2(n106939), .A(n82679), .ZN(n82281) );
  NAND2_X1 U68094 ( .A1(n82681), .A2(n82680), .ZN(n82679) );
  NOR4_X1 U68099 ( .A1(n82691), .A2(n82690), .A3(n82692), .A4(n82693), .ZN(
        n82680) );
  XOR2_X1 U68100 ( .A(n100420), .B(n59451), .Z(n82693) );
  XOR2_X1 U68101 ( .A(n100418), .B(n59445), .Z(n82692) );
  XOR2_X1 U68103 ( .A(n62662), .B(n59453), .Z(n82690) );
  NOR4_X1 U68104 ( .A1(n82695), .A2(n82696), .A3(n82697), .A4(n82698), .ZN(
        n82663) );
  NAND2_X1 U68105 ( .A1(n82699), .A2(n82700), .ZN(n82698) );
  NOR4_X1 U68106 ( .A1(\DLX_Datapath/next_A_IDEX[16] ), .A2(
        \DLX_Datapath/next_A_IDEX[15] ), .A3(\DLX_Datapath/next_A_IDEX[14] ), 
        .A4(\DLX_Datapath/next_A_IDEX[13] ), .ZN(n82700) );
  NOR4_X1 U68107 ( .A1(\DLX_Datapath/next_A_IDEX[12] ), .A2(
        \DLX_Datapath/next_A_IDEX[11] ), .A3(\DLX_Datapath/next_A_IDEX[10] ), 
        .A4(\DLX_Datapath/next_A_IDEX[0] ), .ZN(n82699) );
  NAND2_X1 U68108 ( .A1(n82701), .A2(n82702), .ZN(n82697) );
  NOR4_X1 U68109 ( .A1(\DLX_Datapath/next_A_IDEX[23] ), .A2(
        \DLX_Datapath/next_A_IDEX[22] ), .A3(\DLX_Datapath/next_A_IDEX[21] ), 
        .A4(\DLX_Datapath/next_A_IDEX[20] ), .ZN(n82702) );
  NOR4_X1 U68110 ( .A1(\DLX_Datapath/next_A_IDEX[1] ), .A2(
        \DLX_Datapath/next_A_IDEX[19] ), .A3(\DLX_Datapath/next_A_IDEX[18] ), 
        .A4(\DLX_Datapath/next_A_IDEX[17] ), .ZN(n82701) );
  NAND2_X1 U68111 ( .A1(n82703), .A2(n82704), .ZN(n82696) );
  NOR4_X1 U68112 ( .A1(\DLX_Datapath/next_A_IDEX[30] ), .A2(
        \DLX_Datapath/next_A_IDEX[2] ), .A3(\DLX_Datapath/next_A_IDEX[29] ), 
        .A4(\DLX_Datapath/next_A_IDEX[28] ), .ZN(n82704) );
  NOR4_X1 U68113 ( .A1(\DLX_Datapath/next_A_IDEX[27] ), .A2(
        \DLX_Datapath/next_A_IDEX[26] ), .A3(\DLX_Datapath/next_A_IDEX[25] ), 
        .A4(\DLX_Datapath/next_A_IDEX[24] ), .ZN(n82703) );
  NAND2_X1 U68114 ( .A1(n82705), .A2(n82706), .ZN(n82695) );
  NOR4_X1 U68115 ( .A1(\DLX_Datapath/next_A_IDEX[9] ), .A2(
        \DLX_Datapath/next_A_IDEX[8] ), .A3(\DLX_Datapath/next_A_IDEX[7] ), 
        .A4(\DLX_Datapath/next_A_IDEX[6] ), .ZN(n82706) );
  NOR4_X1 U68116 ( .A1(\DLX_Datapath/next_A_IDEX[5] ), .A2(
        \DLX_Datapath/next_A_IDEX[4] ), .A3(\DLX_Datapath/next_A_IDEX[3] ), 
        .A4(\DLX_Datapath/next_A_IDEX[31] ), .ZN(n82705) );
  NOR2_X1 U68117 ( .A1(n82659), .A2(n106807), .ZN(n82605) );
  OAI21_X1 U68118 ( .B1(n61666), .B2(n82708), .A(n82709), .ZN(n82707) );
  OR2_X1 U68119 ( .A1(n82710), .A2(n110959), .ZN(n82709) );
  NOR4_X1 U68120 ( .A1(n82711), .A2(n82712), .A3(n82713), .A4(n82714), .ZN(
        n82710) );
  AOI21_X1 U68121 ( .B1(n82715), .B2(n82716), .A(n82594), .ZN(n82714) );
  AOI22_X1 U68122 ( .A1(n105147), .A2(n111008), .B1(n105149), .B2(n111006), 
        .ZN(n82716) );
  AOI22_X1 U68123 ( .A1(n82578), .A2(n111004), .B1(n105146), .B2(n111002), 
        .ZN(n82715) );
  AOI21_X1 U68124 ( .B1(n82717), .B2(n82718), .A(n82597), .ZN(n82713) );
  AOI22_X1 U68125 ( .A1(n105148), .A2(n111015), .B1(n105149), .B2(n111013), 
        .ZN(n82718) );
  AOI22_X1 U68126 ( .A1(n82578), .A2(n111011), .B1(n105146), .B2(n111009), 
        .ZN(n82717) );
  AOI21_X1 U68127 ( .B1(n82719), .B2(n82720), .A(n82600), .ZN(n82712) );
  AOI22_X1 U68128 ( .A1(n105147), .A2(n106812), .B1(n105149), .B2(n110962), 
        .ZN(n82720) );
  AOI22_X1 U68129 ( .A1(n105145), .A2(n110961), .B1(n105146), .B2(n110960), 
        .ZN(n82719) );
  AOI21_X1 U68130 ( .B1(n82721), .B2(n82722), .A(n82616), .ZN(n82711) );
  AOI22_X1 U68131 ( .A1(n105148), .A2(n110988), .B1(n105149), .B2(n110986), 
        .ZN(n82722) );
  AOI22_X1 U68132 ( .A1(n105145), .A2(n110984), .B1(n105146), .B2(n110982), 
        .ZN(n82721) );
  NOR4_X1 U68133 ( .A1(n82723), .A2(n82724), .A3(n82725), .A4(n82726), .ZN(
        n82708) );
  AOI21_X1 U68134 ( .B1(n82727), .B2(n82728), .A(n82594), .ZN(n82726) );
  AOI22_X1 U68135 ( .A1(n105147), .A2(n110995), .B1(n105149), .B2(n110994), 
        .ZN(n82728) );
  AOI22_X1 U68136 ( .A1(n105145), .A2(n110992), .B1(n105146), .B2(n110990), 
        .ZN(n82727) );
  AOI21_X1 U68137 ( .B1(n82729), .B2(n82730), .A(n82597), .ZN(n82725) );
  AOI22_X1 U68138 ( .A1(n105147), .A2(n111001), .B1(n105149), .B2(n111000), 
        .ZN(n82730) );
  AOI22_X1 U68139 ( .A1(n82578), .A2(n110998), .B1(n105146), .B2(n110996), 
        .ZN(n82729) );
  AOI21_X1 U68140 ( .B1(n82731), .B2(n82732), .A(n82600), .ZN(n82724) );
  AOI22_X1 U68141 ( .A1(n105147), .A2(n110973), .B1(n82557), .B2(n110972), 
        .ZN(n82732) );
  AOI22_X1 U68142 ( .A1(n105145), .A2(n110970), .B1(n82602), .B2(n110968), 
        .ZN(n82731) );
  AOI21_X1 U68143 ( .B1(n82733), .B2(n82734), .A(n82616), .ZN(n82723) );
  AOI22_X1 U68144 ( .A1(n105147), .A2(n110980), .B1(n82557), .B2(n110979), 
        .ZN(n82734) );
  AOI22_X1 U68145 ( .A1(n82578), .A2(n110977), .B1(n82602), .B2(n110975), .ZN(
        n82733) );
  OAI21_X1 U68146 ( .B1(n61666), .B2(n82735), .A(n82736), .ZN(n82659) );
  OR2_X1 U68147 ( .A1(n82737), .A2(n110959), .ZN(n82736) );
  NOR4_X1 U68148 ( .A1(n82738), .A2(n82739), .A3(n82740), .A4(n82741), .ZN(
        n82737) );
  AOI21_X1 U68149 ( .B1(n82742), .B2(n82743), .A(n82594), .ZN(n82741) );
  AOI22_X1 U68150 ( .A1(n105148), .A2(n111007), .B1(n82557), .B2(n111005), 
        .ZN(n82743) );
  AOI22_X1 U68151 ( .A1(n105145), .A2(n111003), .B1(n82602), .B2(n111043), 
        .ZN(n82742) );
  AOI21_X1 U68152 ( .B1(n82744), .B2(n82745), .A(n82597), .ZN(n82740) );
  AOI22_X1 U68153 ( .A1(n105148), .A2(n111014), .B1(n105149), .B2(n111012), 
        .ZN(n82745) );
  AOI22_X1 U68154 ( .A1(n82578), .A2(n111010), .B1(n105146), .B2(n111044), 
        .ZN(n82744) );
  AOI21_X1 U68155 ( .B1(n82746), .B2(n82747), .A(n82600), .ZN(n82739) );
  AOI22_X1 U68156 ( .A1(n105148), .A2(n107150), .B1(n82557), .B2(n109320), 
        .ZN(n82747) );
  AOI22_X1 U68157 ( .A1(n105145), .A2(n109318), .B1(n82602), .B2(n109319), 
        .ZN(n82746) );
  AOI21_X1 U68158 ( .B1(n82748), .B2(n82749), .A(n82616), .ZN(n82738) );
  AOI22_X1 U68159 ( .A1(n105147), .A2(n110987), .B1(n82557), .B2(n110985), 
        .ZN(n82749) );
  AOI22_X1 U68160 ( .A1(n105145), .A2(n110983), .B1(n82602), .B2(n110981), 
        .ZN(n82748) );
  NOR4_X1 U68161 ( .A1(n82750), .A2(n82751), .A3(n82752), .A4(n82753), .ZN(
        n82735) );
  AOI21_X1 U68162 ( .B1(n82754), .B2(n82755), .A(n82594), .ZN(n82753) );
  NAND2_X1 U68163 ( .A1(n106809), .A2(n110967), .ZN(n82594) );
  AOI22_X1 U68164 ( .A1(n105148), .A2(n111045), .B1(n105149), .B2(n110993), 
        .ZN(n82755) );
  AOI22_X1 U68165 ( .A1(n82578), .A2(n110991), .B1(n105146), .B2(n110989), 
        .ZN(n82754) );
  AOI21_X1 U68166 ( .B1(n82756), .B2(n82757), .A(n82597), .ZN(n82752) );
  NAND2_X1 U68167 ( .A1(n59420), .A2(n110967), .ZN(n82597) );
  AOI22_X1 U68168 ( .A1(n105147), .A2(n111046), .B1(n105149), .B2(n110999), 
        .ZN(n82757) );
  AOI22_X1 U68169 ( .A1(n105145), .A2(n110997), .B1(n82602), .B2(n111041), 
        .ZN(n82756) );
  AOI21_X1 U68170 ( .B1(n82758), .B2(n82759), .A(n82600), .ZN(n82751) );
  NAND2_X1 U68171 ( .A1(n59421), .A2(n106809), .ZN(n82600) );
  AOI22_X1 U68172 ( .A1(n105148), .A2(n111047), .B1(n105149), .B2(n110971), 
        .ZN(n82759) );
  AOI22_X1 U68173 ( .A1(n82578), .A2(n110969), .B1(n105146), .B2(n111042), 
        .ZN(n82758) );
  AOI21_X1 U68174 ( .B1(n82760), .B2(n82761), .A(n82616), .ZN(n82750) );
  NAND2_X1 U68175 ( .A1(n59421), .A2(n59420), .ZN(n82616) );
  AOI22_X1 U68176 ( .A1(n105147), .A2(n111048), .B1(n82557), .B2(n110978), 
        .ZN(n82761) );
  NOR2_X1 U68177 ( .A1(n108971), .A2(n59423), .ZN(n82557) );
  AOI22_X1 U68179 ( .A1(n105145), .A2(n110976), .B1(n82602), .B2(n110974), 
        .ZN(n82760) );
  NOR2_X1 U68180 ( .A1(n109317), .A2(n108971), .ZN(n82602) );
  NOR2_X1 U68181 ( .A1(n109317), .A2(n59422), .ZN(n82578) );
  NOR4_X1 U68182 ( .A1(n111130), .A2(n80086), .A3(n111140), .A4(n80073), .ZN(
        n82651) );
  NAND2_X1 U68183 ( .A1(n82762), .A2(n82763), .ZN(n80073) );
  AOI21_X1 U68184 ( .B1(n111129), .B2(n111146), .A(n80071), .ZN(n82763) );
  NOR2_X1 U68185 ( .A1(n80039), .A2(n111144), .ZN(n80071) );
  OAI21_X1 U68186 ( .B1(IR_in[28]), .B2(n80064), .A(n82646), .ZN(n82764) );
  AOI21_X1 U68187 ( .B1(n111146), .B2(IR_in[28]), .A(n111145), .ZN(n82646) );
  NAND2_X1 U68188 ( .A1(n82765), .A2(IR_in[31]), .ZN(n80039) );
  NOR2_X1 U68189 ( .A1(IR_in[30]), .A2(IR_in[29]), .ZN(n82765) );
  NOR2_X1 U68190 ( .A1(n80092), .A2(n80069), .ZN(n82762) );
  NOR2_X1 U68192 ( .A1(n82766), .A2(n82629), .ZN(n80056) );
  NAND2_X1 U68193 ( .A1(n111141), .A2(n82639), .ZN(n82766) );
  NAND2_X1 U68194 ( .A1(n80064), .A2(n82628), .ZN(n82639) );
  NAND2_X1 U68195 ( .A1(n82334), .A2(n111145), .ZN(n80100) );
  NAND2_X1 U68196 ( .A1(n82767), .A2(n82768), .ZN(n80092) );
  NOR3_X1 U68197 ( .A1(n82769), .A2(n82006), .A3(n111127), .ZN(n82768) );
  NAND2_X1 U68198 ( .A1(n111129), .A2(n111143), .ZN(n81976) );
  OAI21_X1 U68199 ( .B1(n80042), .B2(n111124), .A(n82645), .ZN(n82769) );
  NAND2_X1 U68200 ( .A1(n82771), .A2(n111148), .ZN(n82645) );
  NOR2_X1 U68201 ( .A1(n82629), .A2(n111141), .ZN(n82771) );
  NOR4_X1 U68202 ( .A1(IR_in[31]), .A2(IR_in[29]), .A3(n111143), .A4(n111141), 
        .ZN(n81974) );
  NOR2_X1 U68203 ( .A1(n82016), .A2(n82772), .ZN(n82767) );
  OAI21_X1 U68204 ( .B1(IR_in[26]), .B2(n82770), .A(n82647), .ZN(n82772) );
  AOI21_X1 U68205 ( .B1(n111147), .B2(n82006), .A(n82005), .ZN(n82647) );
  NOR4_X1 U68208 ( .A1(IR_in[31]), .A2(IR_in[28]), .A3(n111142), .A4(n111141), 
        .ZN(n82006) );
  NAND2_X1 U68209 ( .A1(n82775), .A2(IR_in[29]), .ZN(n82770) );
  NOR2_X1 U68210 ( .A1(IR_in[31]), .A2(IR_in[30]), .ZN(n82775) );
  OAI33_X1 U68211 ( .A1(n80064), .A2(n82629), .A3(n111141), .B1(n81993), .B2(
        n82774), .B3(n111123), .ZN(n82016) );
  NOR2_X1 U68212 ( .A1(n111145), .A2(n80042), .ZN(n82774) );
  NOR2_X1 U68213 ( .A1(n111149), .A2(IR_in[27]), .ZN(n80042) );
  NAND2_X1 U68214 ( .A1(n111149), .A2(n111146), .ZN(n82628) );
  NAND2_X1 U68215 ( .A1(n82776), .A2(IR_in[30]), .ZN(n81993) );
  NOR2_X1 U68216 ( .A1(n111143), .A2(n111142), .ZN(n82776) );
  NAND2_X1 U68217 ( .A1(n82777), .A2(IR_in[29]), .ZN(n82629) );
  NOR2_X1 U68218 ( .A1(IR_in[28]), .A2(n111123), .ZN(n82777) );
  NAND2_X1 U68219 ( .A1(n82778), .A2(n111148), .ZN(n81887) );
  NOR2_X1 U68220 ( .A1(n80067), .A2(n111141), .ZN(n82778) );
  NAND2_X1 U68223 ( .A1(n82780), .A2(n82781), .ZN(n82332) );
  NOR3_X1 U68224 ( .A1(IR_in[29]), .A2(IR_in[31]), .A3(IR_in[30]), .ZN(n82781)
         );
  NOR2_X1 U68225 ( .A1(IR_in[27]), .A2(n111143), .ZN(n82780) );
  OAI21_X1 U68226 ( .B1(n100416), .B2(n105221), .A(n82782), .ZN(n59081) );
  NAND2_X1 U68227 ( .A1(n105221), .A2(n69289), .ZN(n82782) );
  OAI21_X1 U68228 ( .B1(n64652), .B2(n111106), .A(n82783), .ZN(n59080) );
  NAND2_X1 U68229 ( .A1(n82784), .A2(n106766), .ZN(n82783) );
  OAI21_X1 U68230 ( .B1(n100417), .B2(n61904), .A(n82785), .ZN(n59078) );
  NAND2_X1 U68231 ( .A1(n100417), .A2(n69303), .ZN(n82785) );
  OAI21_X1 U68232 ( .B1(n64652), .B2(n106837), .A(n82786), .ZN(n59077) );
  AOI22_X1 U68233 ( .A1(n82787), .A2(n61904), .B1(n107155), .B2(n106830), .ZN(
        n82786) );
  NOR2_X1 U68234 ( .A1(n58713), .A2(n82789), .ZN(n82787) );
  OAI21_X1 U68235 ( .B1(n59516), .B2(n106509), .A(n82790), .ZN(n59073) );
  NAND2_X1 U68236 ( .A1(n69346), .A2(n106509), .ZN(n82790) );
  OAI21_X1 U68237 ( .B1(n58722), .B2(Rst), .A(n82791), .ZN(n59072) );
  NAND2_X1 U68238 ( .A1(Rst), .A2(n69346), .ZN(n82791) );
  OAI21_X1 U68239 ( .B1(n105012), .B2(n106509), .A(n82792), .ZN(n59071) );
  NAND2_X1 U68240 ( .A1(n69347), .A2(n106514), .ZN(n82792) );
  OAI21_X1 U68241 ( .B1(n58720), .B2(Rst), .A(n82793), .ZN(n59070) );
  NAND2_X1 U68242 ( .A1(Rst), .A2(n69347), .ZN(n82793) );
  OAI21_X1 U68243 ( .B1(n59518), .B2(n106509), .A(n82794), .ZN(n59069) );
  NAND2_X1 U68244 ( .A1(n69348), .A2(n106509), .ZN(n82794) );
  OAI21_X1 U68245 ( .B1(Rst), .B2(n107109), .A(n82795), .ZN(n59068) );
  NAND2_X1 U68246 ( .A1(Rst), .A2(n69348), .ZN(n82795) );
  OAI21_X1 U68247 ( .B1(n100417), .B2(n100794), .A(n82796), .ZN(n59061) );
  NAND2_X1 U68248 ( .A1(n105221), .A2(n69413), .ZN(n82796) );
  OAI21_X1 U68249 ( .B1(n100417), .B2(n100800), .A(n82797), .ZN(n59060) );
  NAND2_X1 U68250 ( .A1(n105221), .A2(n69414), .ZN(n82797) );
  OAI21_X1 U68251 ( .B1(n100417), .B2(n58713), .A(n82798), .ZN(n59059) );
  NAND2_X1 U68252 ( .A1(n105221), .A2(n69415), .ZN(n82798) );
  OAI21_X1 U68253 ( .B1(n100417), .B2(n59346), .A(n82799), .ZN(n59058) );
  NAND2_X1 U68254 ( .A1(n105221), .A2(n69416), .ZN(n82799) );
  OAI21_X1 U68255 ( .B1(n100417), .B2(n59342), .A(n82800), .ZN(n59057) );
  NAND2_X1 U68256 ( .A1(n105221), .A2(n69417), .ZN(n82800) );
  OAI21_X1 U68257 ( .B1(n105222), .B2(n100653), .A(n82801), .ZN(n59054) );
  NAND2_X1 U68258 ( .A1(n100414), .A2(DataAddr[29]), .ZN(n82801) );
  OAI21_X1 U68259 ( .B1(n105222), .B2(n100711), .A(n82802), .ZN(n59053) );
  NAND2_X1 U68260 ( .A1(n105222), .A2(DataAddr[0]), .ZN(n82802) );
  NAND2_X1 U68261 ( .A1(n82803), .A2(n82804), .ZN(n59050) );
  AOI22_X1 U68262 ( .A1(DataIn_hw[6]), .A2(n105144), .B1(DataIn_b[6]), .B2(
        n111052), .ZN(n82804) );
  AOI22_X1 U68263 ( .A1(DataIn_w[6]), .A2(n105886), .B1(n69699), .B2(n111053), 
        .ZN(n82803) );
  NAND2_X1 U68264 ( .A1(n82807), .A2(n82808), .ZN(n59049) );
  AOI22_X1 U68265 ( .A1(DataIn_hw[5]), .A2(n82805), .B1(DataIn_b[5]), .B2(
        n111052), .ZN(n82808) );
  AOI22_X1 U68266 ( .A1(DataIn_w[5]), .A2(n105886), .B1(n69700), .B2(n111053), 
        .ZN(n82807) );
  NAND2_X1 U68267 ( .A1(n82809), .A2(n82810), .ZN(n59048) );
  AOI22_X1 U68268 ( .A1(DataIn_hw[4]), .A2(n105144), .B1(DataIn_b[4]), .B2(
        n111052), .ZN(n82810) );
  AOI22_X1 U68269 ( .A1(DataIn_w[4]), .A2(n105886), .B1(n69701), .B2(n111053), 
        .ZN(n82809) );
  NAND2_X1 U68270 ( .A1(n82811), .A2(n82812), .ZN(n59047) );
  AOI22_X1 U68271 ( .A1(DataIn_hw[3]), .A2(n82805), .B1(DataIn_b[3]), .B2(
        n111052), .ZN(n82812) );
  AOI22_X1 U68272 ( .A1(DataIn_w[3]), .A2(n105886), .B1(n69702), .B2(n111053), 
        .ZN(n82811) );
  NAND2_X1 U68273 ( .A1(n82813), .A2(n82814), .ZN(n59046) );
  AOI22_X1 U68274 ( .A1(DataIn_hw[2]), .A2(n105144), .B1(DataIn_b[2]), .B2(
        n111052), .ZN(n82814) );
  AOI22_X1 U68275 ( .A1(DataIn_w[2]), .A2(n105886), .B1(n69703), .B2(n111053), 
        .ZN(n82813) );
  NAND2_X1 U68276 ( .A1(n82815), .A2(n82816), .ZN(n59045) );
  AOI22_X1 U68277 ( .A1(DataIn_hw[1]), .A2(n82805), .B1(DataIn_b[1]), .B2(
        n111052), .ZN(n82816) );
  AOI22_X1 U68278 ( .A1(DataIn_w[1]), .A2(n105886), .B1(n69704), .B2(n111053), 
        .ZN(n82815) );
  NAND2_X1 U68279 ( .A1(n82817), .A2(n82818), .ZN(n59044) );
  AOI22_X1 U68280 ( .A1(DataIn_hw[0]), .A2(n105144), .B1(DataIn_b[0]), .B2(
        n111052), .ZN(n82818) );
  AOI22_X1 U68281 ( .A1(DataIn_w[0]), .A2(n105886), .B1(n69705), .B2(n111053), 
        .ZN(n82817) );
  NAND2_X1 U68282 ( .A1(n82819), .A2(n82820), .ZN(n59043) );
  AOI21_X1 U68283 ( .B1(DataIn_hw[9]), .B2(n105144), .A(n82821), .ZN(n82820)
         );
  AOI22_X1 U68284 ( .A1(DataIn_w[9]), .A2(n105886), .B1(n69706), .B2(n111053), 
        .ZN(n82819) );
  NAND2_X1 U68285 ( .A1(n82822), .A2(n82823), .ZN(n59042) );
  AOI21_X1 U68286 ( .B1(DataIn_hw[8]), .B2(n82805), .A(n82821), .ZN(n82823) );
  AOI22_X1 U68287 ( .A1(DataIn_w[8]), .A2(n105886), .B1(n69707), .B2(n111053), 
        .ZN(n82822) );
  OAI21_X1 U68288 ( .B1(n69697), .B2(n107370), .A(n82824), .ZN(n59041) );
  AOI21_X1 U68289 ( .B1(DataIn_w[31]), .B2(n82806), .A(n82821), .ZN(n82824) );
  OAI21_X1 U68290 ( .B1(n69697), .B2(n107372), .A(n82825), .ZN(n59040) );
  AOI21_X1 U68291 ( .B1(DataIn_w[30]), .B2(n82806), .A(n82821), .ZN(n82825) );
  OAI21_X1 U68292 ( .B1(n69697), .B2(n107374), .A(n82826), .ZN(n59039) );
  AOI21_X1 U68293 ( .B1(DataIn_w[29]), .B2(n82806), .A(n82821), .ZN(n82826) );
  OAI21_X1 U68294 ( .B1(n69697), .B2(n107375), .A(n82827), .ZN(n59038) );
  AOI21_X1 U68295 ( .B1(DataIn_w[28]), .B2(n82806), .A(n82821), .ZN(n82827) );
  OAI21_X1 U68296 ( .B1(n69697), .B2(n107377), .A(n82828), .ZN(n59037) );
  AOI21_X1 U68297 ( .B1(DataIn_w[27]), .B2(n82806), .A(n82821), .ZN(n82828) );
  OAI21_X1 U68298 ( .B1(n69697), .B2(n107379), .A(n82829), .ZN(n59036) );
  AOI21_X1 U68299 ( .B1(DataIn_w[26]), .B2(n82806), .A(n82821), .ZN(n82829) );
  OAI21_X1 U68300 ( .B1(n69697), .B2(n107381), .A(n82830), .ZN(n59035) );
  AOI21_X1 U68301 ( .B1(DataIn_w[25]), .B2(n105886), .A(n82821), .ZN(n82830)
         );
  OAI21_X1 U68302 ( .B1(n69697), .B2(n107383), .A(n82831), .ZN(n59034) );
  AOI21_X1 U68303 ( .B1(DataIn_w[24]), .B2(n82806), .A(n82821), .ZN(n82831) );
  OAI21_X1 U68304 ( .B1(n69697), .B2(n107385), .A(n82832), .ZN(n59033) );
  AOI21_X1 U68305 ( .B1(DataIn_w[23]), .B2(n105886), .A(n82821), .ZN(n82832)
         );
  OAI21_X1 U68306 ( .B1(n69697), .B2(n107387), .A(n82833), .ZN(n59032) );
  AOI21_X1 U68307 ( .B1(DataIn_w[22]), .B2(n105886), .A(n82821), .ZN(n82833)
         );
  OAI21_X1 U68308 ( .B1(n69697), .B2(n107389), .A(n82834), .ZN(n59031) );
  AOI21_X1 U68309 ( .B1(DataIn_w[21]), .B2(n105886), .A(n82821), .ZN(n82834)
         );
  OAI21_X1 U68310 ( .B1(n69697), .B2(n107391), .A(n82835), .ZN(n59030) );
  AOI21_X1 U68311 ( .B1(DataIn_w[20]), .B2(n82806), .A(n82821), .ZN(n82835) );
  OAI21_X1 U68312 ( .B1(n69697), .B2(n107393), .A(n82836), .ZN(n59029) );
  AOI21_X1 U68313 ( .B1(DataIn_w[19]), .B2(n105886), .A(n82821), .ZN(n82836)
         );
  OAI21_X1 U68314 ( .B1(n69697), .B2(n107395), .A(n82837), .ZN(n59028) );
  AOI21_X1 U68315 ( .B1(DataIn_w[18]), .B2(n82806), .A(n82821), .ZN(n82837) );
  OAI21_X1 U68316 ( .B1(n69697), .B2(n107397), .A(n82838), .ZN(n59027) );
  AOI21_X1 U68317 ( .B1(DataIn_w[17]), .B2(n82806), .A(n82821), .ZN(n82838) );
  OAI21_X1 U68318 ( .B1(n69697), .B2(n107399), .A(n82839), .ZN(n59026) );
  AOI21_X1 U68319 ( .B1(DataIn_w[16]), .B2(n82806), .A(n82821), .ZN(n82839) );
  NAND2_X1 U68320 ( .A1(n82840), .A2(n82841), .ZN(n59025) );
  AOI21_X1 U68321 ( .B1(DataIn_hw[15]), .B2(n105144), .A(n82821), .ZN(n82841)
         );
  AOI22_X1 U68322 ( .A1(DataIn_w[15]), .A2(n105886), .B1(n69724), .B2(n111053), 
        .ZN(n82840) );
  NAND2_X1 U68323 ( .A1(n82842), .A2(n82843), .ZN(n59024) );
  AOI21_X1 U68324 ( .B1(DataIn_hw[14]), .B2(n82805), .A(n82821), .ZN(n82843)
         );
  AOI22_X1 U68325 ( .A1(DataIn_w[14]), .A2(n105886), .B1(n69725), .B2(n111053), 
        .ZN(n82842) );
  NAND2_X1 U68326 ( .A1(n82844), .A2(n82845), .ZN(n59023) );
  AOI21_X1 U68327 ( .B1(DataIn_hw[13]), .B2(n105144), .A(n82821), .ZN(n82845)
         );
  AOI22_X1 U68328 ( .A1(DataIn_w[13]), .A2(n105886), .B1(n69726), .B2(n111053), 
        .ZN(n82844) );
  NAND2_X1 U68329 ( .A1(n82846), .A2(n82847), .ZN(n59022) );
  AOI21_X1 U68330 ( .B1(DataIn_hw[12]), .B2(n82805), .A(n82821), .ZN(n82847)
         );
  AOI22_X1 U68331 ( .A1(DataIn_w[12]), .A2(n105886), .B1(n69727), .B2(n111053), 
        .ZN(n82846) );
  NAND2_X1 U68332 ( .A1(n82848), .A2(n82849), .ZN(n59021) );
  AOI21_X1 U68333 ( .B1(DataIn_hw[11]), .B2(n105144), .A(n82821), .ZN(n82849)
         );
  AOI22_X1 U68334 ( .A1(DataIn_w[11]), .A2(n105886), .B1(n69728), .B2(n111053), 
        .ZN(n82848) );
  NAND2_X1 U68335 ( .A1(n82850), .A2(n82851), .ZN(n59020) );
  AOI21_X1 U68336 ( .B1(DataIn_hw[10]), .B2(n82805), .A(n82821), .ZN(n82851)
         );
  NOR2_X1 U68338 ( .A1(n111065), .A2(n82853), .ZN(n82852) );
  AOI22_X1 U68339 ( .A1(DataIn_w[10]), .A2(n105886), .B1(n69729), .B2(n111053), 
        .ZN(n82850) );
  NAND2_X1 U68340 ( .A1(n82854), .A2(n82855), .ZN(n59019) );
  AOI22_X1 U68341 ( .A1(DataIn_hw[7]), .A2(n82805), .B1(DataIn_b[7]), .B2(
        n111052), .ZN(n82855) );
  NAND2_X1 U68342 ( .A1(n69698), .A2(n69697), .ZN(n82853) );
  NOR2_X1 U68343 ( .A1(n82856), .A2(n111053), .ZN(n82805) );
  AOI22_X1 U68345 ( .A1(DataIn_w[7]), .A2(n105886), .B1(n69730), .B2(n111053), 
        .ZN(n82854) );
  NOR2_X1 U68346 ( .A1(n82857), .A2(n111053), .ZN(n82806) );
  NAND2_X1 U68348 ( .A1(n82858), .A2(n82859), .ZN(n59013) );
  AOI22_X1 U68349 ( .A1(n82860), .A2(n111070), .B1(n82861), .B2(n69710), .ZN(
        n82859) );
  AOI22_X1 U68350 ( .A1(n82862), .A2(n69307), .B1(n107413), .B2(n107414), .ZN(
        n82858) );
  NAND2_X1 U68351 ( .A1(n82863), .A2(n82864), .ZN(n59012) );
  AOI22_X1 U68352 ( .A1(n82860), .A2(n111087), .B1(n82861), .B2(n69705), .ZN(
        n82864) );
  AOI22_X1 U68353 ( .A1(n82862), .A2(n69292), .B1(n107413), .B2(n107415), .ZN(
        n82863) );
  OAI21_X1 U68354 ( .B1(n100417), .B2(n59334), .A(n82865), .ZN(n59009) );
  NAND2_X1 U68355 ( .A1(n105221), .A2(n69991), .ZN(n82865) );
  OAI21_X1 U68356 ( .B1(n64652), .B2(n107631), .A(n82866), .ZN(n59008) );
  AOI22_X1 U68357 ( .A1(n107630), .A2(n108277), .B1(n59335), .B2(n82867), .ZN(
        n82866) );
  OAI21_X1 U68358 ( .B1(n100414), .B2(n100687), .A(n82869), .ZN(n59006) );
  NAND2_X1 U68359 ( .A1(n100414), .A2(DataAddr[12]), .ZN(n82869) );
  NAND2_X1 U68360 ( .A1(n82870), .A2(n82871), .ZN(n59005) );
  AOI22_X1 U68361 ( .A1(n82860), .A2(n111097), .B1(n82861), .B2(n69727), .ZN(
        n82871) );
  AOI22_X1 U68362 ( .A1(n82862), .A2(n70130), .B1(n107413), .B2(n107741), .ZN(
        n82870) );
  OAI21_X1 U68363 ( .B1(n100417), .B2(n59350), .A(n82872), .ZN(n59004) );
  NAND2_X1 U68364 ( .A1(n105221), .A2(n70142), .ZN(n82872) );
  OAI21_X1 U68365 ( .B1(n64652), .B2(n107749), .A(n82873), .ZN(n59003) );
  AOI21_X1 U68366 ( .B1(n82874), .B2(n107152), .A(n82875), .ZN(n82873) );
  NOR3_X1 U68367 ( .A1(n107152), .A2(n100800), .A3(n106831), .ZN(n82875) );
  OAI21_X1 U68368 ( .B1(n82789), .B2(n107153), .A(n106829), .ZN(n82874) );
  OAI21_X1 U68369 ( .B1(n64652), .B2(n107750), .A(n82878), .ZN(n59002) );
  AOI22_X1 U68370 ( .A1(n100800), .A2(n82876), .B1(n82877), .B2(n107153), .ZN(
        n82878) );
  OAI21_X1 U68371 ( .B1(n82789), .B2(n106830), .A(n82788), .ZN(n82877) );
  AOI21_X1 U68372 ( .B1(n107160), .B2(n58713), .A(n82879), .ZN(n82788) );
  NOR3_X1 U68373 ( .A1(n82789), .A2(n61904), .A3(n58713), .ZN(n82876) );
  OAI21_X1 U68374 ( .B1(n64652), .B2(n107751), .A(n82880), .ZN(n59001) );
  AOI22_X1 U68375 ( .A1(n82879), .A2(n107154), .B1(n58713), .B2(n107160), .ZN(
        n82880) );
  NAND2_X1 U68376 ( .A1(n82881), .A2(n82882), .ZN(n82789) );
  NOR2_X1 U68377 ( .A1(n59350), .A2(n82883), .ZN(n82881) );
  OAI21_X1 U68378 ( .B1(n82884), .B2(n82885), .A(n82886), .ZN(n82879) );
  NOR3_X1 U68379 ( .A1(n82883), .A2(n59350), .A3(n82887), .ZN(n82884) );
  OAI21_X1 U68380 ( .B1(n100414), .B2(n100655), .A(n82888), .ZN(n58999) );
  NAND2_X1 U68381 ( .A1(n100414), .A2(DataAddr[28]), .ZN(n82888) );
  NAND2_X1 U68382 ( .A1(n82889), .A2(n82890), .ZN(n58998) );
  AOI22_X1 U68383 ( .A1(n82860), .A2(n111091), .B1(n82861), .B2(n69711), .ZN(
        n82890) );
  AOI22_X1 U68384 ( .A1(n82862), .A2(n70283), .B1(n107413), .B2(n107853), .ZN(
        n82889) );
  OAI21_X1 U68385 ( .B1(n100414), .B2(n100649), .A(n82891), .ZN(n58996) );
  NAND2_X1 U68386 ( .A1(n100414), .A2(DataAddr[31]), .ZN(n82891) );
  NAND2_X1 U68387 ( .A1(n82892), .A2(n82893), .ZN(n58995) );
  AOI22_X1 U68388 ( .A1(n82860), .A2(n111069), .B1(n82861), .B2(n69708), .ZN(
        n82893) );
  AOI22_X1 U68389 ( .A1(n82862), .A2(n70427), .B1(n107413), .B2(n107948), .ZN(
        n82892) );
  OAI21_X1 U68390 ( .B1(n100414), .B2(n100651), .A(n82894), .ZN(n58993) );
  NAND2_X1 U68391 ( .A1(n100414), .A2(DataAddr[30]), .ZN(n82894) );
  NAND2_X1 U68392 ( .A1(n82895), .A2(n82896), .ZN(n58992) );
  AOI22_X1 U68393 ( .A1(n82860), .A2(n111090), .B1(n82861), .B2(n69709), .ZN(
        n82896) );
  AOI22_X1 U68394 ( .A1(n82862), .A2(n70569), .B1(n107413), .B2(n108044), .ZN(
        n82895) );
  OAI21_X1 U68395 ( .B1(n100414), .B2(n100657), .A(n82897), .ZN(n58990) );
  NAND2_X1 U68396 ( .A1(n100414), .A2(DataAddr[27]), .ZN(n82897) );
  OAI21_X1 U68397 ( .B1(n100414), .B2(n100659), .A(n82898), .ZN(n58988) );
  NAND2_X1 U68398 ( .A1(n100414), .A2(DataAddr[26]), .ZN(n82898) );
  OAI21_X1 U68399 ( .B1(n100417), .B2(n59347), .A(n82899), .ZN(n58987) );
  NAND2_X1 U68400 ( .A1(n105221), .A2(n70575), .ZN(n82899) );
  OAI21_X1 U68401 ( .B1(n100417), .B2(n59348), .A(n82900), .ZN(n58986) );
  NAND2_X1 U68402 ( .A1(n105221), .A2(n70576), .ZN(n82900) );
  OAI21_X1 U68403 ( .B1(n100417), .B2(n59349), .A(n82901), .ZN(n58985) );
  NAND2_X1 U68404 ( .A1(n105221), .A2(n70577), .ZN(n82901) );
  OAI21_X1 U68405 ( .B1(n64652), .B2(n108053), .A(n82902), .ZN(n58984) );
  AOI21_X1 U68406 ( .B1(n107158), .B2(n108052), .A(n82903), .ZN(n82902) );
  NOR4_X1 U68407 ( .A1(n59348), .A2(n59347), .A3(n107159), .A4(n108052), .ZN(
        n82903) );
  NAND2_X1 U68408 ( .A1(n82905), .A2(n82906), .ZN(n58983) );
  AOI22_X1 U68409 ( .A1(n82860), .A2(n111093), .B1(n82861), .B2(n69713), .ZN(
        n82906) );
  AOI22_X1 U68410 ( .A1(n82862), .A2(n70717), .B1(n107413), .B2(n108154), .ZN(
        n82905) );
  OAI21_X1 U68411 ( .B1(n105222), .B2(n100661), .A(n82907), .ZN(n58981) );
  NAND2_X1 U68412 ( .A1(n100414), .A2(DataAddr[25]), .ZN(n82907) );
  OAI21_X1 U68413 ( .B1(n105222), .B2(n100663), .A(n82908), .ZN(n58979) );
  NAND2_X1 U68414 ( .A1(n100414), .A2(DataAddr[24]), .ZN(n82908) );
  OAI21_X1 U68415 ( .B1(n105222), .B2(n100681), .A(n82909), .ZN(n58977) );
  NAND2_X1 U68416 ( .A1(n100414), .A2(DataAddr[15]), .ZN(n82909) );
  OAI21_X1 U68417 ( .B1(n100417), .B2(n59338), .A(n82910), .ZN(n58976) );
  NAND2_X1 U68418 ( .A1(n105221), .A2(n70726), .ZN(n82910) );
  OAI21_X1 U68419 ( .B1(n64652), .B2(n111116), .A(n82911), .ZN(n58975) );
  AOI21_X1 U68420 ( .B1(n82912), .B2(n108159), .A(n82913), .ZN(n82911) );
  NOR3_X1 U68421 ( .A1(n108159), .A2(n59337), .A3(n82914), .ZN(n82913) );
  OAI21_X1 U68422 ( .B1(n107628), .B2(n108281), .A(n82915), .ZN(n82912) );
  NAND2_X1 U68423 ( .A1(n82916), .A2(n82917), .ZN(n58974) );
  AOI22_X1 U68424 ( .A1(n82860), .A2(n111096), .B1(n82861), .B2(n69724), .ZN(
        n82917) );
  AOI22_X1 U68425 ( .A1(n82862), .A2(n70872), .B1(n107413), .B2(n108270), .ZN(
        n82916) );
  OAI21_X1 U68426 ( .B1(n105222), .B2(n100683), .A(n82918), .ZN(n58972) );
  NAND2_X1 U68427 ( .A1(n100414), .A2(DataAddr[14]), .ZN(n82918) );
  OAI21_X1 U68428 ( .B1(n100417), .B2(n59335), .A(n82919), .ZN(n58971) );
  NAND2_X1 U68429 ( .A1(n105221), .A2(n70880), .ZN(n82919) );
  OAI21_X1 U68430 ( .B1(n100417), .B2(n59336), .A(n82920), .ZN(n58970) );
  NAND2_X1 U68431 ( .A1(n100417), .A2(n70882), .ZN(n82920) );
  OAI21_X1 U68432 ( .B1(n100417), .B2(n59337), .A(n82921), .ZN(n58969) );
  NAND2_X1 U68433 ( .A1(n100417), .A2(n70884), .ZN(n82921) );
  OAI21_X1 U68434 ( .B1(n64652), .B2(n108282), .A(n82922), .ZN(n58968) );
  AOI22_X1 U68435 ( .A1(n82923), .A2(n59336), .B1(n82924), .B2(n108279), .ZN(
        n82922) );
  NOR2_X1 U68436 ( .A1(n59335), .A2(n107628), .ZN(n82923) );
  OAI21_X1 U68437 ( .B1(n64652), .B2(n111117), .A(n82925), .ZN(n58967) );
  AOI22_X1 U68438 ( .A1(n59337), .A2(n107629), .B1(n107627), .B2(n108281), 
        .ZN(n82925) );
  AOI21_X1 U68439 ( .B1(n82867), .B2(n59336), .A(n82924), .ZN(n82915) );
  OAI21_X1 U68440 ( .B1(n107628), .B2(n108277), .A(n82868), .ZN(n82924) );
  AOI21_X1 U68441 ( .B1(n82926), .B2(n111051), .A(n111049), .ZN(n82868) );
  NAND2_X1 U68442 ( .A1(n82927), .A2(n82867), .ZN(n82914) );
  NOR2_X1 U68443 ( .A1(n82885), .A2(n82926), .ZN(n82867) );
  NOR2_X1 U68444 ( .A1(n59336), .A2(n59335), .ZN(n82927) );
  NAND2_X1 U68445 ( .A1(n82928), .A2(n82929), .ZN(n58966) );
  AOI22_X1 U68446 ( .A1(n82860), .A2(n111079), .B1(n82861), .B2(n69725), .ZN(
        n82929) );
  AOI22_X1 U68447 ( .A1(n105885), .A2(n71026), .B1(n107413), .B2(n108391), 
        .ZN(n82928) );
  OAI21_X1 U68448 ( .B1(n105222), .B2(n100685), .A(n82930), .ZN(n58964) );
  NAND2_X1 U68449 ( .A1(n100414), .A2(DataAddr[13]), .ZN(n82930) );
  NAND2_X1 U68450 ( .A1(n82931), .A2(n82932), .ZN(n58963) );
  AOI22_X1 U68451 ( .A1(n82860), .A2(n111080), .B1(n82861), .B2(n69726), .ZN(
        n82932) );
  AOI22_X1 U68452 ( .A1(n82862), .A2(n71169), .B1(n107413), .B2(n108500), .ZN(
        n82931) );
  OAI21_X1 U68453 ( .B1(n105222), .B2(n100689), .A(n82933), .ZN(n58961) );
  NAND2_X1 U68454 ( .A1(n100414), .A2(DataAddr[11]), .ZN(n82933) );
  OAI21_X1 U68455 ( .B1(n105222), .B2(n100691), .A(n82934), .ZN(n58959) );
  NAND2_X1 U68456 ( .A1(n100414), .A2(DataAddr[10]), .ZN(n82934) );
  OAI21_X1 U68457 ( .B1(n100417), .B2(n59333), .A(n82935), .ZN(n58958) );
  NAND2_X1 U68458 ( .A1(n100417), .A2(n71179), .ZN(n82935) );
  OAI21_X1 U68459 ( .B1(n64652), .B2(n108510), .A(n82936), .ZN(n58957) );
  AOI22_X1 U68460 ( .A1(n59333), .A2(n108629), .B1(n108627), .B2(n108509), 
        .ZN(n82936) );
  OAI21_X1 U68461 ( .B1(n105222), .B2(n100705), .A(n82939), .ZN(n58955) );
  NAND2_X1 U68462 ( .A1(n100414), .A2(DataAddr[3]), .ZN(n82939) );
  OAI21_X1 U68463 ( .B1(n100413), .B2(n105221), .A(n82940), .ZN(n58954) );
  NAND2_X1 U68464 ( .A1(n100417), .A2(n71325), .ZN(n82940) );
  OAI21_X1 U68465 ( .B1(n100417), .B2(n58643), .A(n82941), .ZN(n58953) );
  NAND2_X1 U68466 ( .A1(n100417), .A2(n71327), .ZN(n82941) );
  OAI21_X1 U68467 ( .B1(n100417), .B2(n100799), .A(n82942), .ZN(n58952) );
  NAND2_X1 U68468 ( .A1(n100417), .A2(n71329), .ZN(n82942) );
  OAI21_X1 U68469 ( .B1(n64652), .B2(n111109), .A(n82943), .ZN(n58951) );
  NAND2_X1 U68470 ( .A1(n82784), .A2(n108620), .ZN(n82943) );
  NAND2_X1 U68471 ( .A1(n82886), .A2(n82885), .ZN(n82784) );
  OAI21_X1 U68472 ( .B1(n64652), .B2(n111108), .A(n82944), .ZN(n58950) );
  AOI22_X1 U68473 ( .A1(n58643), .A2(n111051), .B1(n111049), .B2(n108622), 
        .ZN(n82944) );
  OAI21_X1 U68474 ( .B1(n64652), .B2(n111107), .A(n82945), .ZN(n58949) );
  AOI22_X1 U68475 ( .A1(n82946), .A2(n100799), .B1(n82947), .B2(n108632), .ZN(
        n82945) );
  OAI21_X1 U68476 ( .B1(n82885), .B2(n108622), .A(n82886), .ZN(n82947) );
  NOR2_X1 U68477 ( .A1(n58643), .A2(n82885), .ZN(n82946) );
  NAND2_X1 U68478 ( .A1(n82948), .A2(n82949), .ZN(n58948) );
  AOI22_X1 U68479 ( .A1(n82860), .A2(n111084), .B1(n82861), .B2(n69702), .ZN(
        n82949) );
  AOI22_X1 U68480 ( .A1(n82862), .A2(n71469), .B1(n107413), .B2(n108739), .ZN(
        n82948) );
  OAI21_X1 U68481 ( .B1(n100414), .B2(n100709), .A(n82950), .ZN(n58946) );
  NAND2_X1 U68482 ( .A1(n100414), .A2(DataAddr[1]), .ZN(n82950) );
  NAND2_X1 U68483 ( .A1(n82951), .A2(n82952), .ZN(n58945) );
  AOI22_X1 U68484 ( .A1(n82860), .A2(n111086), .B1(n82861), .B2(n69704), .ZN(
        n82952) );
  AOI22_X1 U68485 ( .A1(n82862), .A2(n71618), .B1(n107413), .B2(n108854), .ZN(
        n82951) );
  OAI21_X1 U68486 ( .B1(n100414), .B2(n100707), .A(n82953), .ZN(n58943) );
  NAND2_X1 U68487 ( .A1(n100414), .A2(DataAddr[2]), .ZN(n82953) );
  NAND2_X1 U68488 ( .A1(n82954), .A2(n82955), .ZN(n58942) );
  AOI22_X1 U68489 ( .A1(n82860), .A2(n111085), .B1(n82861), .B2(n69703), .ZN(
        n82955) );
  AOI22_X1 U68490 ( .A1(n105885), .A2(n71762), .B1(n107413), .B2(n108965), 
        .ZN(n82954) );
  OAI21_X1 U68491 ( .B1(n105222), .B2(n100697), .A(n82956), .ZN(n58940) );
  NAND2_X1 U68492 ( .A1(n100414), .A2(DataAddr[7]), .ZN(n82956) );
  OAI21_X1 U68493 ( .B1(n100417), .B2(n59330), .A(n82957), .ZN(n58939) );
  NAND2_X1 U68494 ( .A1(n100417), .A2(n71772), .ZN(n82957) );
  OAI21_X1 U68495 ( .B1(n64652), .B2(n108975), .A(n82958), .ZN(n58938) );
  AOI21_X1 U68496 ( .B1(n82959), .B2(n108973), .A(n82960), .ZN(n82958) );
  NOR3_X1 U68497 ( .A1(n108973), .A2(n59329), .A3(n82961), .ZN(n82960) );
  OAI21_X1 U68498 ( .B1(n108625), .B2(n109097), .A(n108624), .ZN(n82959) );
  NAND2_X1 U68499 ( .A1(n82963), .A2(n82964), .ZN(n58937) );
  AOI22_X1 U68500 ( .A1(n82860), .A2(n111088), .B1(n82861), .B2(n69730), .ZN(
        n82964) );
  AOI22_X1 U68501 ( .A1(n105885), .A2(n71913), .B1(n107413), .B2(n109084), 
        .ZN(n82963) );
  OAI21_X1 U68502 ( .B1(n100414), .B2(n100699), .A(n82965), .ZN(n58935) );
  NAND2_X1 U68503 ( .A1(n100414), .A2(DataAddr[6]), .ZN(n82965) );
  OAI21_X1 U68504 ( .B1(n100417), .B2(n59327), .A(n82966), .ZN(n58934) );
  NAND2_X1 U68505 ( .A1(n100417), .A2(n71922), .ZN(n82966) );
  OAI21_X1 U68506 ( .B1(n100417), .B2(n59328), .A(n82967), .ZN(n58933) );
  NAND2_X1 U68507 ( .A1(n100417), .A2(n71924), .ZN(n82967) );
  OAI21_X1 U68508 ( .B1(n100417), .B2(n59329), .A(n82968), .ZN(n58932) );
  NAND2_X1 U68509 ( .A1(n100417), .A2(n71926), .ZN(n82968) );
  OAI21_X1 U68510 ( .B1(n64652), .B2(n111115), .A(n82969), .ZN(n58931) );
  AOI22_X1 U68511 ( .A1(n82970), .A2(n109093), .B1(n59327), .B2(n82971), .ZN(
        n82969) );
  OAI21_X1 U68512 ( .B1(n100414), .B2(n100703), .A(n82972), .ZN(n58929) );
  NAND2_X1 U68513 ( .A1(n100414), .A2(DataAddr[4]), .ZN(n82972) );
  NAND2_X1 U68514 ( .A1(n82973), .A2(n82974), .ZN(n58928) );
  AOI22_X1 U68515 ( .A1(n82860), .A2(n111089), .B1(n82861), .B2(n69701), .ZN(
        n82974) );
  AOI22_X1 U68516 ( .A1(n105885), .A2(n72065), .B1(n107413), .B2(n109203), 
        .ZN(n82973) );
  OAI21_X1 U68517 ( .B1(n64652), .B2(n111114), .A(n82975), .ZN(n58927) );
  AOI21_X1 U68518 ( .B1(n108623), .B2(n109095), .A(n82976), .ZN(n82975) );
  NOR3_X1 U68519 ( .A1(n109095), .A2(n59327), .A3(n108625), .ZN(n82976) );
  OAI21_X1 U68520 ( .B1(n100414), .B2(n100701), .A(n82978), .ZN(n58925) );
  NAND2_X1 U68521 ( .A1(n100414), .A2(DataAddr[5]), .ZN(n82978) );
  NAND2_X1 U68522 ( .A1(n82979), .A2(n82980), .ZN(n58924) );
  AOI22_X1 U68523 ( .A1(n82860), .A2(n111077), .B1(n82861), .B2(n69700), .ZN(
        n82980) );
  AOI22_X1 U68524 ( .A1(n105885), .A2(n72209), .B1(n107413), .B2(n109312), 
        .ZN(n82979) );
  OAI21_X1 U68525 ( .B1(n64652), .B2(n111113), .A(n82981), .ZN(n58923) );
  AOI22_X1 U68526 ( .A1(n59329), .A2(n108626), .B1(n82962), .B2(n109097), .ZN(
        n82981) );
  OAI21_X1 U68527 ( .B1(n108625), .B2(n109095), .A(n82977), .ZN(n82962) );
  AOI21_X1 U68528 ( .B1(n82971), .B2(n59327), .A(n82970), .ZN(n82977) );
  OAI21_X1 U68529 ( .B1(n82982), .B2(n82885), .A(n82886), .ZN(n82970) );
  NOR2_X1 U68530 ( .A1(n58643), .A2(n100799), .ZN(n82982) );
  NAND2_X1 U68531 ( .A1(n82983), .A2(n82971), .ZN(n82961) );
  NOR3_X1 U68532 ( .A1(n82885), .A2(n100799), .A3(n58643), .ZN(n82971) );
  NOR2_X1 U68533 ( .A1(n59328), .A2(n59327), .ZN(n82983) );
  NAND2_X1 U68534 ( .A1(n82984), .A2(n82985), .ZN(n58922) );
  AOI22_X1 U68535 ( .A1(n82860), .A2(n111083), .B1(n82861), .B2(n69699), .ZN(
        n82985) );
  AOI22_X1 U68536 ( .A1(n105885), .A2(n72362), .B1(n107413), .B2(n109431), 
        .ZN(n82984) );
  OAI21_X1 U68537 ( .B1(n100414), .B2(n100693), .A(n82986), .ZN(n58920) );
  NAND2_X1 U68538 ( .A1(n100414), .A2(DataAddr[9]), .ZN(n82986) );
  OAI21_X1 U68539 ( .B1(n100417), .B2(n59331), .A(n82987), .ZN(n58919) );
  NAND2_X1 U68540 ( .A1(n100417), .A2(n72370), .ZN(n82987) );
  OAI21_X1 U68541 ( .B1(n100417), .B2(n59332), .A(n82988), .ZN(n58918) );
  NAND2_X1 U68542 ( .A1(n100417), .A2(n72372), .ZN(n82988) );
  OAI21_X1 U68543 ( .B1(n64652), .B2(n111112), .A(n82989), .ZN(n58917) );
  AOI22_X1 U68544 ( .A1(n108630), .A2(n109436), .B1(n59331), .B2(n82990), .ZN(
        n82989) );
  OAI21_X1 U68545 ( .B1(n100414), .B2(n100695), .A(n82992), .ZN(n58915) );
  NAND2_X1 U68546 ( .A1(n100414), .A2(DataAddr[8]), .ZN(n82992) );
  NAND2_X1 U68547 ( .A1(n82993), .A2(n82994), .ZN(n58914) );
  AOI22_X1 U68548 ( .A1(n82860), .A2(n111076), .B1(n82861), .B2(n69707), .ZN(
        n82994) );
  AOI22_X1 U68549 ( .A1(n105885), .A2(n72511), .B1(n107413), .B2(n109544), 
        .ZN(n82993) );
  OAI21_X1 U68550 ( .B1(n64652), .B2(n111110), .A(n82995), .ZN(n58913) );
  AOI21_X1 U68551 ( .B1(n82996), .B2(n107622), .A(n82997), .ZN(n82995) );
  NOR3_X1 U68552 ( .A1(n107622), .A2(n59333), .A3(n82938), .ZN(n82997) );
  NAND2_X1 U68553 ( .A1(n82998), .A2(n82990), .ZN(n82938) );
  NOR2_X1 U68554 ( .A1(n59332), .A2(n59331), .ZN(n82998) );
  OAI21_X1 U68555 ( .B1(n108628), .B2(n108509), .A(n82937), .ZN(n82996) );
  AOI21_X1 U68556 ( .B1(n82990), .B2(n59332), .A(n82999), .ZN(n82937) );
  NAND2_X1 U68557 ( .A1(n83000), .A2(n83001), .ZN(n58912) );
  AOI22_X1 U68558 ( .A1(n82860), .A2(n111081), .B1(n82861), .B2(n69728), .ZN(
        n83001) );
  AOI22_X1 U68559 ( .A1(n105885), .A2(n72661), .B1(n107413), .B2(n109654), 
        .ZN(n83000) );
  OAI21_X1 U68560 ( .B1(n64652), .B2(n111111), .A(n83002), .ZN(n58911) );
  AOI22_X1 U68561 ( .A1(n83003), .A2(n59332), .B1(n82999), .B2(n109438), .ZN(
        n83002) );
  OAI21_X1 U68562 ( .B1(n108628), .B2(n109436), .A(n82991), .ZN(n82999) );
  AOI21_X1 U68563 ( .B1(n83004), .B2(n111051), .A(n111049), .ZN(n82991) );
  NOR2_X1 U68564 ( .A1(n59331), .A2(n108628), .ZN(n83003) );
  NOR2_X1 U68565 ( .A1(n82885), .A2(n83004), .ZN(n82990) );
  NAND2_X1 U68566 ( .A1(n83005), .A2(n83006), .ZN(n58910) );
  AOI22_X1 U68567 ( .A1(n82860), .A2(n111075), .B1(n82861), .B2(n69706), .ZN(
        n83006) );
  AOI22_X1 U68568 ( .A1(n105885), .A2(n72803), .B1(n107413), .B2(n109761), 
        .ZN(n83005) );
  NAND2_X1 U68569 ( .A1(n83007), .A2(n83008), .ZN(n58909) );
  AOI22_X1 U68570 ( .A1(n82860), .A2(n111082), .B1(n82861), .B2(n69729), .ZN(
        n83008) );
  AOI22_X1 U68571 ( .A1(n105885), .A2(n72808), .B1(n107413), .B2(n109766), 
        .ZN(n83007) );
  OAI21_X1 U68572 ( .B1(n100414), .B2(n100673), .A(n83009), .ZN(n58907) );
  NAND2_X1 U68573 ( .A1(n100414), .A2(DataAddr[19]), .ZN(n83009) );
  OAI21_X1 U68574 ( .B1(n105222), .B2(n100675), .A(n83010), .ZN(n58905) );
  NAND2_X1 U68575 ( .A1(n100414), .A2(DataAddr[18]), .ZN(n83010) );
  OAI21_X1 U68576 ( .B1(n105222), .B2(n100677), .A(n83011), .ZN(n58903) );
  NAND2_X1 U68577 ( .A1(n100414), .A2(DataAddr[17]), .ZN(n83011) );
  OAI21_X1 U68578 ( .B1(n100417), .B2(n59341), .A(n83012), .ZN(n58902) );
  NAND2_X1 U68579 ( .A1(n100417), .A2(n72830), .ZN(n83012) );
  OAI21_X1 U68580 ( .B1(n64652), .B2(n109785), .A(n83013), .ZN(n58901) );
  AOI22_X1 U68581 ( .A1(n107626), .A2(n109900), .B1(n59339), .B2(n83014), .ZN(
        n83013) );
  OAI21_X1 U68582 ( .B1(n105222), .B2(n100679), .A(n83016), .ZN(n58899) );
  NAND2_X1 U68583 ( .A1(n100414), .A2(DataAddr[16]), .ZN(n83016) );
  NAND2_X1 U68584 ( .A1(n83017), .A2(n83018), .ZN(n58898) );
  AOI22_X1 U68585 ( .A1(n82860), .A2(n111074), .B1(n82861), .B2(n69723), .ZN(
        n83018) );
  AOI22_X1 U68586 ( .A1(n105885), .A2(n72969), .B1(n107413), .B2(n109895), 
        .ZN(n83017) );
  OAI21_X1 U68587 ( .B1(n100417), .B2(n59339), .A(n83019), .ZN(n58897) );
  NAND2_X1 U68588 ( .A1(n100417), .A2(n72978), .ZN(n83019) );
  OAI21_X1 U68589 ( .B1(n100417), .B2(n59340), .A(n83020), .ZN(n58896) );
  NAND2_X1 U68590 ( .A1(n100417), .A2(n72980), .ZN(n83020) );
  OAI21_X1 U68591 ( .B1(n64652), .B2(n109903), .A(n83021), .ZN(n58895) );
  AOI22_X1 U68592 ( .A1(n83022), .A2(n59340), .B1(n83023), .B2(n109902), .ZN(
        n83021) );
  NOR2_X1 U68593 ( .A1(n59339), .A2(n107624), .ZN(n83022) );
  NAND2_X1 U68594 ( .A1(n83024), .A2(n83025), .ZN(n58894) );
  AOI22_X1 U68595 ( .A1(n82860), .A2(n111078), .B1(n82861), .B2(n69722), .ZN(
        n83025) );
  AOI22_X1 U68596 ( .A1(n105885), .A2(n73120), .B1(n107413), .B2(n110010), 
        .ZN(n83024) );
  OAI21_X1 U68597 ( .B1(n64652), .B2(n110012), .A(n83026), .ZN(n58893) );
  AOI21_X1 U68598 ( .B1(n83027), .B2(n107161), .A(n83028), .ZN(n83026) );
  NOR3_X1 U68599 ( .A1(n107161), .A2(n59341), .A3(n83029), .ZN(n83028) );
  OAI21_X1 U68600 ( .B1(n107624), .B2(n109784), .A(n83030), .ZN(n83027) );
  NAND2_X1 U68601 ( .A1(n83031), .A2(n83032), .ZN(n58892) );
  AOI22_X1 U68602 ( .A1(n82860), .A2(n111072), .B1(n82861), .B2(n69720), .ZN(
        n83032) );
  AOI22_X1 U68603 ( .A1(n105885), .A2(n73263), .B1(n107413), .B2(n110119), 
        .ZN(n83031) );
  OAI21_X1 U68604 ( .B1(n64652), .B2(n110120), .A(n83033), .ZN(n58891) );
  AOI22_X1 U68605 ( .A1(n59341), .A2(n107625), .B1(n107623), .B2(n109784), 
        .ZN(n83033) );
  AOI21_X1 U68606 ( .B1(n83014), .B2(n59340), .A(n83023), .ZN(n83030) );
  OAI21_X1 U68607 ( .B1(n107624), .B2(n109900), .A(n83015), .ZN(n83023) );
  AOI21_X1 U68608 ( .B1(n83034), .B2(n111051), .A(n111049), .ZN(n83015) );
  NAND2_X1 U68609 ( .A1(n83035), .A2(n83014), .ZN(n83029) );
  NOR2_X1 U68610 ( .A1(n82885), .A2(n83034), .ZN(n83014) );
  NOR2_X1 U68611 ( .A1(n59340), .A2(n59339), .ZN(n83035) );
  NAND2_X1 U68612 ( .A1(n83036), .A2(n83037), .ZN(n58890) );
  AOI22_X1 U68613 ( .A1(n82860), .A2(n111073), .B1(n82861), .B2(n69721), .ZN(
        n83037) );
  AOI22_X1 U68614 ( .A1(n105885), .A2(n73405), .B1(n107413), .B2(n110226), 
        .ZN(n83036) );
  OAI21_X1 U68615 ( .B1(n100414), .B2(n100665), .A(n83038), .ZN(n58888) );
  NAND2_X1 U68616 ( .A1(n100414), .A2(DataAddr[23]), .ZN(n83038) );
  OAI21_X1 U68617 ( .B1(n100414), .B2(n100667), .A(n83039), .ZN(n58886) );
  NAND2_X1 U68618 ( .A1(n100414), .A2(DataAddr[22]), .ZN(n83039) );
  OAI21_X1 U68619 ( .B1(n100417), .B2(n59345), .A(n83040), .ZN(n58885) );
  NAND2_X1 U68620 ( .A1(n100417), .A2(n73411), .ZN(n83040) );
  OAI21_X1 U68621 ( .B1(n64652), .B2(n110230), .A(n83041), .ZN(n58884) );
  AOI22_X1 U68622 ( .A1(n59345), .A2(n107164), .B1(n107162), .B2(n110229), 
        .ZN(n83041) );
  NAND2_X1 U68623 ( .A1(n83044), .A2(n83045), .ZN(n58883) );
  AOI22_X1 U68624 ( .A1(n82860), .A2(n111066), .B1(n82861), .B2(n69717), .ZN(
        n83045) );
  AOI22_X1 U68625 ( .A1(n105885), .A2(n73552), .B1(n107413), .B2(n110332), 
        .ZN(n83044) );
  OAI21_X1 U68626 ( .B1(n100414), .B2(n100669), .A(n83046), .ZN(n58881) );
  NAND2_X1 U68627 ( .A1(n100414), .A2(DataAddr[21]), .ZN(n83046) );
  OAI21_X1 U68628 ( .B1(n100417), .B2(n59343), .A(n83047), .ZN(n58880) );
  NAND2_X1 U68629 ( .A1(n100417), .A2(n73558), .ZN(n83047) );
  OAI21_X1 U68630 ( .B1(n100417), .B2(n59344), .A(n83048), .ZN(n58879) );
  NAND2_X1 U68631 ( .A1(n100417), .A2(n73560), .ZN(n83048) );
  OAI21_X1 U68632 ( .B1(n64652), .B2(n110338), .A(n83049), .ZN(n58878) );
  AOI22_X1 U68633 ( .A1(n107165), .A2(n110335), .B1(n59343), .B2(n83050), .ZN(
        n83049) );
  OAI21_X1 U68634 ( .B1(n100414), .B2(n100671), .A(n83052), .ZN(n58876) );
  NAND2_X1 U68635 ( .A1(n100414), .A2(DataAddr[20]), .ZN(n83052) );
  NAND2_X1 U68636 ( .A1(n83053), .A2(n83054), .ZN(n58875) );
  AOI22_X1 U68637 ( .A1(n82860), .A2(n111068), .B1(n82861), .B2(n69719), .ZN(
        n83054) );
  AOI22_X1 U68638 ( .A1(n105885), .A2(n73699), .B1(n107413), .B2(n110439), 
        .ZN(n83053) );
  OAI21_X1 U68639 ( .B1(n64652), .B2(n110447), .A(n83055), .ZN(n58874) );
  AOI21_X1 U68640 ( .B1(n83056), .B2(n107156), .A(n83057), .ZN(n83055) );
  NOR3_X1 U68641 ( .A1(n107156), .A2(n59345), .A3(n83043), .ZN(n83057) );
  NAND2_X1 U68642 ( .A1(n83058), .A2(n83050), .ZN(n83043) );
  NOR2_X1 U68643 ( .A1(n59344), .A2(n59343), .ZN(n83058) );
  OAI21_X1 U68644 ( .B1(n107163), .B2(n110229), .A(n83042), .ZN(n83056) );
  AOI21_X1 U68645 ( .B1(n83050), .B2(n59344), .A(n83059), .ZN(n83042) );
  NAND2_X1 U68646 ( .A1(n83060), .A2(n83061), .ZN(n58873) );
  AOI22_X1 U68647 ( .A1(n82860), .A2(n111071), .B1(n82861), .B2(n69716), .ZN(
        n83061) );
  AOI22_X1 U68648 ( .A1(n105885), .A2(n73847), .B1(n107413), .B2(n110546), 
        .ZN(n83060) );
  OAI21_X1 U68649 ( .B1(n64652), .B2(n110547), .A(n83062), .ZN(n58872) );
  AOI22_X1 U68650 ( .A1(n83063), .A2(n59344), .B1(n83059), .B2(n110337), .ZN(
        n83062) );
  OAI21_X1 U68651 ( .B1(n107163), .B2(n110335), .A(n83051), .ZN(n83059) );
  AOI21_X1 U68652 ( .B1(n83064), .B2(n111051), .A(n111049), .ZN(n83051) );
  NOR2_X1 U68653 ( .A1(n59343), .A2(n107163), .ZN(n83063) );
  NOR2_X1 U68654 ( .A1(n82885), .A2(n83064), .ZN(n83050) );
  NAND2_X1 U68655 ( .A1(n83065), .A2(n83066), .ZN(n58871) );
  AOI22_X1 U68656 ( .A1(n82860), .A2(n111067), .B1(n82861), .B2(n69718), .ZN(
        n83066) );
  AOI22_X1 U68657 ( .A1(n105885), .A2(n73988), .B1(n107413), .B2(n110652), 
        .ZN(n83065) );
  OAI21_X1 U68658 ( .B1(n64652), .B2(n110654), .A(n83067), .ZN(n58870) );
  AOI21_X1 U68659 ( .B1(n83068), .B2(n107748), .A(n83069), .ZN(n83067) );
  NOR3_X1 U68660 ( .A1(n107748), .A2(n82883), .A3(n107159), .ZN(n83069) );
  NAND2_X1 U68661 ( .A1(n83070), .A2(n108048), .ZN(n82883) );
  NOR2_X1 U68662 ( .A1(n59349), .A2(n59348), .ZN(n83070) );
  OAI21_X1 U68663 ( .B1(n107159), .B2(n108052), .A(n82904), .ZN(n83068) );
  AOI21_X1 U68664 ( .B1(n82882), .B2(n59348), .A(n83071), .ZN(n82904) );
  NAND2_X1 U68665 ( .A1(n83072), .A2(n83073), .ZN(n58869) );
  AOI22_X1 U68666 ( .A1(n82860), .A2(n111092), .B1(n82861), .B2(n69712), .ZN(
        n83073) );
  AOI22_X1 U68667 ( .A1(n105885), .A2(n74130), .B1(n107413), .B2(n110750), 
        .ZN(n83072) );
  OAI21_X1 U68668 ( .B1(n64652), .B2(n110751), .A(n83074), .ZN(n58868) );
  AOI21_X1 U68669 ( .B1(n83071), .B2(n108050), .A(n83075), .ZN(n83074) );
  NOR3_X1 U68670 ( .A1(n108050), .A2(n59347), .A3(n107159), .ZN(n83075) );
  OAI21_X1 U68671 ( .B1(n107159), .B2(n108048), .A(n83076), .ZN(n83071) );
  NAND2_X1 U68672 ( .A1(n83077), .A2(n83078), .ZN(n58867) );
  AOI22_X1 U68673 ( .A1(n82860), .A2(n111094), .B1(n82861), .B2(n69714), .ZN(
        n83078) );
  AOI22_X1 U68674 ( .A1(n105885), .A2(n74270), .B1(n107413), .B2(n110851), 
        .ZN(n83077) );
  OAI21_X1 U68675 ( .B1(n64652), .B2(n110852), .A(n83079), .ZN(n58866) );
  AOI22_X1 U68676 ( .A1(n107157), .A2(n108048), .B1(n59347), .B2(n82882), .ZN(
        n83079) );
  NOR2_X1 U68677 ( .A1(n82885), .A2(n82887), .ZN(n82882) );
  AOI21_X1 U68678 ( .B1(n82887), .B2(n111051), .A(n111049), .ZN(n83076) );
  NAND2_X1 U68679 ( .A1(n64652), .A2(n111050), .ZN(n82886) );
  NAND2_X1 U68680 ( .A1(n100415), .A2(n64652), .ZN(n82885) );
  NAND2_X1 U68681 ( .A1(n83080), .A2(n83081), .ZN(n82887) );
  NOR3_X1 U68682 ( .A1(n59344), .A2(n59346), .A3(n59345), .ZN(n83081) );
  NOR2_X1 U68683 ( .A1(n59343), .A2(n83064), .ZN(n83080) );
  NAND2_X1 U68684 ( .A1(n83082), .A2(n83083), .ZN(n83064) );
  NOR3_X1 U68685 ( .A1(n59340), .A2(n59342), .A3(n59341), .ZN(n83083) );
  NOR2_X1 U68686 ( .A1(n59339), .A2(n83034), .ZN(n83082) );
  NAND2_X1 U68687 ( .A1(n83084), .A2(n83085), .ZN(n83034) );
  NOR3_X1 U68688 ( .A1(n59336), .A2(n59338), .A3(n59337), .ZN(n83085) );
  NOR2_X1 U68689 ( .A1(n59335), .A2(n82926), .ZN(n83084) );
  NAND2_X1 U68690 ( .A1(n83086), .A2(n83087), .ZN(n82926) );
  NOR3_X1 U68691 ( .A1(n59332), .A2(n59334), .A3(n59333), .ZN(n83087) );
  NOR2_X1 U68692 ( .A1(n59331), .A2(n83004), .ZN(n83086) );
  NAND2_X1 U68693 ( .A1(n83088), .A2(n83089), .ZN(n83004) );
  NOR3_X1 U68694 ( .A1(n59329), .A2(n100799), .A3(n59330), .ZN(n83089) );
  NOR3_X1 U68695 ( .A1(n58643), .A2(n59328), .A3(n59327), .ZN(n83088) );
  NAND2_X1 U68696 ( .A1(n83090), .A2(n83091), .ZN(n58865) );
  AOI22_X1 U68697 ( .A1(n82860), .A2(n111095), .B1(n82861), .B2(n69715), .ZN(
        n83091) );
  AND2_X2 U68698 ( .A1(n83092), .A2(n83093), .ZN(n82861) );
  NOR3_X1 U68699 ( .A1(n83094), .A2(n83095), .A3(n106935), .ZN(n83093) );
  NOR2_X1 U68700 ( .A1(n83096), .A2(n107413), .ZN(n83092) );
  AND2_X2 U68701 ( .A1(n62027), .A2(n83097), .ZN(n82860) );
  AOI22_X1 U68702 ( .A1(n105885), .A2(n74410), .B1(n107413), .B2(n110952), 
        .ZN(n83090) );
  NOR2_X1 U68703 ( .A1(n83098), .A2(n107413), .ZN(n82862) );
  OR2_X1 U68704 ( .A1(n83097), .A2(n83099), .ZN(n83098) );
  NOR4_X1 U68705 ( .A1(n83095), .A2(n106935), .A3(n83094), .A4(n83096), .ZN(
        n83099) );
  NAND2_X1 U68707 ( .A1(n83101), .A2(n83102), .ZN(n83096) );
  NOR2_X1 U68708 ( .A1(n69322), .A2(n59419), .ZN(n83101) );
  OAI21_X1 U68710 ( .B1(n69326), .B2(n59415), .A(n83104), .ZN(n83094) );
  AOI21_X1 U68711 ( .B1(n107062), .B2(n83105), .A(n83106), .ZN(n83103) );
  NAND4_X2 U68712 ( .A1(n83107), .A2(n83108), .A3(n83109), .A4(n83110), .ZN(
        n58864) );
  NOR3_X1 U68713 ( .A1(n83111), .A2(n83112), .A3(n83113), .ZN(n83110) );
  AOI21_X1 U68715 ( .B1(n83115), .B2(n83116), .A(n106326), .ZN(n83112) );
  NOR4_X1 U68716 ( .A1(n83117), .A2(n83118), .A3(n83119), .A4(n83120), .ZN(
        n83116) );
  OAI21_X1 U68717 ( .B1(n100775), .B2(n105168), .A(n83121), .ZN(n83120) );
  AOI22_X1 U68718 ( .A1(n83122), .A2(n107878), .B1(n105883), .B2(n107882), 
        .ZN(n83121) );
  NAND2_X1 U68719 ( .A1(n83124), .A2(n83125), .ZN(n83119) );
  AOI22_X1 U68720 ( .A1(n105882), .A2(n107886), .B1(n105881), .B2(n70343), 
        .ZN(n83125) );
  AOI22_X1 U68721 ( .A1(n105880), .A2(n107918), .B1(n70331), .B2(n105879), 
        .ZN(n83124) );
  OAI21_X1 U68722 ( .B1(n100992), .B2(n105167), .A(n83130), .ZN(n83118) );
  AOI22_X1 U68723 ( .A1(n105878), .A2(n107907), .B1(n70355), .B2(n105877), 
        .ZN(n83130) );
  NAND2_X1 U68724 ( .A1(n83133), .A2(n83134), .ZN(n83117) );
  AOI22_X1 U68725 ( .A1(n83135), .A2(n107915), .B1(n70383), .B2(n105875), .ZN(
        n83134) );
  AOI22_X1 U68726 ( .A1(n70367), .A2(n105874), .B1(n105873), .B2(n107903), 
        .ZN(n83133) );
  NOR4_X1 U68727 ( .A1(n83139), .A2(n83140), .A3(n83141), .A4(n83142), .ZN(
        n83115) );
  OAI21_X1 U68728 ( .B1(n103912), .B2(n105872), .A(n83144), .ZN(n83142) );
  NAND2_X1 U68730 ( .A1(n83147), .A2(n83148), .ZN(n83141) );
  AOI22_X1 U68731 ( .A1(n83149), .A2(n107929), .B1(n70291), .B2(n83150), .ZN(
        n83148) );
  AOI22_X1 U68732 ( .A1(n83151), .A2(n107932), .B1(n83152), .B2(n107876), .ZN(
        n83147) );
  OAI21_X1 U68733 ( .B1(n103911), .B2(n106741), .A(n83153), .ZN(n83140) );
  AOI22_X1 U68734 ( .A1(n70303), .A2(n105866), .B1(n70295), .B2(n83155), .ZN(
        n83153) );
  NAND2_X1 U68735 ( .A1(n83156), .A2(n83157), .ZN(n83139) );
  AOI22_X1 U68736 ( .A1(n83158), .A2(n107891), .B1(n105862), .B2(n107874), 
        .ZN(n83157) );
  AOI22_X1 U68737 ( .A1(n105861), .A2(n107870), .B1(n105860), .B2(n107866), 
        .ZN(n83156) );
  AND2_X2 U68738 ( .A1(n105859), .A2(n70402), .ZN(n83111) );
  AOI22_X1 U68739 ( .A1(n83163), .A2(n107860), .B1(n105856), .B2(n107872), 
        .ZN(n83109) );
  AOI22_X1 U68740 ( .A1(n105855), .A2(n107910), .B1(n105854), .B2(n107940), 
        .ZN(n83108) );
  AOI22_X1 U68741 ( .A1(n106287), .A2(n107891), .B1(n70331), .B2(n106282), 
        .ZN(n83107) );
  NAND4_X2 U68742 ( .A1(n83167), .A2(n83168), .A3(n83169), .A4(n83170), .ZN(
        n58863) );
  NOR3_X1 U68743 ( .A1(n83171), .A2(n83172), .A3(n83173), .ZN(n83170) );
  NOR2_X1 U68744 ( .A1(n103890), .A2(n106737), .ZN(n83173) );
  AOI21_X1 U68745 ( .B1(n83174), .B2(n83175), .A(n106324), .ZN(n83172) );
  NOR4_X1 U68746 ( .A1(n83176), .A2(n83177), .A3(n83178), .A4(n83179), .ZN(
        n83175) );
  OAI21_X1 U68747 ( .B1(n103893), .B2(n106739), .A(n83180), .ZN(n83179) );
  AOI22_X1 U68748 ( .A1(n105884), .A2(n107975), .B1(n105883), .B2(n107977), 
        .ZN(n83180) );
  NAND2_X1 U68749 ( .A1(n83181), .A2(n83182), .ZN(n83178) );
  AOI22_X1 U68750 ( .A1(n105882), .A2(n107981), .B1(n70485), .B2(n105881), 
        .ZN(n83182) );
  AOI22_X1 U68751 ( .A1(n105880), .A2(n108015), .B1(n70473), .B2(n105879), 
        .ZN(n83181) );
  OAI21_X1 U68752 ( .B1(n100993), .B2(n105167), .A(n83183), .ZN(n83177) );
  AOI22_X1 U68753 ( .A1(n105878), .A2(n108003), .B1(n70497), .B2(n105877), 
        .ZN(n83183) );
  NAND2_X1 U68754 ( .A1(n83184), .A2(n83185), .ZN(n83176) );
  AOI22_X1 U68755 ( .A1(n83135), .A2(n108012), .B1(n70525), .B2(n105875), .ZN(
        n83185) );
  AOI22_X1 U68756 ( .A1(n105874), .A2(n107996), .B1(n105873), .B2(n107999), 
        .ZN(n83184) );
  NOR4_X1 U68757 ( .A1(n83186), .A2(n83187), .A3(n83188), .A4(n83189), .ZN(
        n83174) );
  OAI21_X1 U68758 ( .B1(n103901), .B2(n83143), .A(n83190), .ZN(n83189) );
  NAND2_X1 U68760 ( .A1(n83191), .A2(n83192), .ZN(n83188) );
  AOI22_X1 U68761 ( .A1(n83149), .A2(n108025), .B1(n70433), .B2(n83150), .ZN(
        n83192) );
  AOI22_X1 U68762 ( .A1(n83151), .A2(n108028), .B1(n83152), .B2(n107973), .ZN(
        n83191) );
  OAI21_X1 U68763 ( .B1(n103900), .B2(n106741), .A(n83193), .ZN(n83187) );
  AOI22_X1 U68764 ( .A1(n70445), .A2(n105866), .B1(n70437), .B2(n105865), .ZN(
        n83193) );
  NAND2_X1 U68765 ( .A1(n83194), .A2(n83195), .ZN(n83186) );
  AOI22_X1 U68766 ( .A1(n83158), .A2(n107986), .B1(n70461), .B2(n105862), .ZN(
        n83195) );
  AOI22_X1 U68767 ( .A1(n83160), .A2(n107967), .B1(n105860), .B2(n107963), 
        .ZN(n83194) );
  AND2_X2 U68768 ( .A1(n105859), .A2(n70544), .ZN(n83171) );
  AOI22_X1 U68769 ( .A1(n83163), .A2(n107957), .B1(n105856), .B2(n107969), 
        .ZN(n83169) );
  AOI22_X1 U68770 ( .A1(n105855), .A2(n108006), .B1(n105854), .B2(n108036), 
        .ZN(n83168) );
  AOI22_X1 U68771 ( .A1(n106287), .A2(n107986), .B1(n70473), .B2(n106282), 
        .ZN(n83167) );
  NAND4_X2 U68772 ( .A1(n83196), .A2(n83197), .A3(n83198), .A4(n83199), .ZN(
        n58862) );
  NOR3_X1 U68773 ( .A1(n83200), .A2(n83201), .A3(n83202), .ZN(n83199) );
  NOR2_X1 U68774 ( .A1(n103874), .A2(n106737), .ZN(n83202) );
  AOI21_X1 U68775 ( .B1(n83203), .B2(n83204), .A(n106324), .ZN(n83201) );
  NOR4_X1 U68776 ( .A1(n83205), .A2(n83206), .A3(n83207), .A4(n83208), .ZN(
        n83204) );
  OAI21_X1 U68777 ( .B1(n103878), .B2(n105168), .A(n83209), .ZN(n83208) );
  AOI22_X1 U68778 ( .A1(n105884), .A2(n107239), .B1(n105883), .B2(n107244), 
        .ZN(n83209) );
  NAND2_X1 U68779 ( .A1(n83210), .A2(n83211), .ZN(n83207) );
  AOI22_X1 U68780 ( .A1(n105882), .A2(n107248), .B1(n69538), .B2(n105881), 
        .ZN(n83211) );
  AOI22_X1 U68781 ( .A1(n105880), .A2(n107285), .B1(n83129), .B2(n69526), .ZN(
        n83210) );
  OAI21_X1 U68782 ( .B1(n100994), .B2(n106738), .A(n83212), .ZN(n83206) );
  AOI22_X1 U68783 ( .A1(n105878), .A2(n107274), .B1(n105877), .B2(n107259), 
        .ZN(n83212) );
  NAND2_X1 U68784 ( .A1(n83213), .A2(n83214), .ZN(n83205) );
  AOI22_X1 U68785 ( .A1(n83135), .A2(n107282), .B1(n69578), .B2(n105875), .ZN(
        n83214) );
  AOI22_X1 U68786 ( .A1(n105874), .A2(n107267), .B1(n105873), .B2(n107270), 
        .ZN(n83213) );
  NOR4_X1 U68787 ( .A1(n83215), .A2(n83216), .A3(n83217), .A4(n83218), .ZN(
        n83203) );
  OAI21_X1 U68788 ( .B1(n103886), .B2(n105872), .A(n83219), .ZN(n83218) );
  NAND2_X1 U68790 ( .A1(n83220), .A2(n83221), .ZN(n83217) );
  AOI22_X1 U68791 ( .A1(n83149), .A2(n107198), .B1(n69486), .B2(n83150), .ZN(
        n83221) );
  AOI22_X1 U68792 ( .A1(n83151), .A2(n107192), .B1(n83152), .B2(n107237), .ZN(
        n83220) );
  OAI21_X1 U68793 ( .B1(n103885), .B2(n106741), .A(n83222), .ZN(n83216) );
  AOI22_X1 U68794 ( .A1(n69498), .A2(n105866), .B1(n105865), .B2(n69490), .ZN(
        n83222) );
  NAND2_X1 U68795 ( .A1(n83223), .A2(n83224), .ZN(n83215) );
  AOI22_X1 U68796 ( .A1(n83158), .A2(n107254), .B1(n69514), .B2(n105862), .ZN(
        n83224) );
  AOI22_X1 U68797 ( .A1(n105861), .A2(n107230), .B1(n105860), .B2(n107226), 
        .ZN(n83223) );
  AND2_X2 U68798 ( .A1(n105859), .A2(n69469), .ZN(n83200) );
  AOI22_X1 U68799 ( .A1(n83163), .A2(n107219), .B1(n105856), .B2(n107232), 
        .ZN(n83198) );
  AOI22_X1 U68800 ( .A1(n105855), .A2(n107277), .B1(n105854), .B2(n107176), 
        .ZN(n83197) );
  AOI22_X1 U68801 ( .A1(n106287), .A2(n107254), .B1(n69526), .B2(n80260), .ZN(
        n83196) );
  NAND4_X2 U68802 ( .A1(n83225), .A2(n83226), .A3(n83227), .A4(n83228), .ZN(
        n58861) );
  NOR3_X1 U68803 ( .A1(n83229), .A2(n83230), .A3(n83231), .ZN(n83228) );
  NOR2_X1 U68804 ( .A1(n103855), .A2(n106737), .ZN(n83231) );
  AOI21_X1 U68805 ( .B1(n83232), .B2(n83233), .A(n106325), .ZN(n83230) );
  NOR4_X1 U68806 ( .A1(n83234), .A2(n83235), .A3(n83236), .A4(n83237), .ZN(
        n83233) );
  OAI21_X1 U68807 ( .B1(n103860), .B2(n105864), .A(n83238), .ZN(n83237) );
  AOI22_X1 U68808 ( .A1(n105883), .A2(n107783), .B1(n83239), .B2(n107795), 
        .ZN(n83238) );
  NAND2_X1 U68809 ( .A1(n83240), .A2(n83241), .ZN(n83236) );
  AOI22_X1 U68810 ( .A1(n70199), .A2(n83127), .B1(n83128), .B2(n107823), .ZN(
        n83241) );
  AOI22_X1 U68811 ( .A1(n70187), .A2(n105879), .B1(n105884), .B2(n107778), 
        .ZN(n83240) );
  NAND2_X1 U68812 ( .A1(n83242), .A2(n83243), .ZN(n83235) );
  AOI22_X1 U68813 ( .A1(n105878), .A2(n107811), .B1(n105877), .B2(n107796), 
        .ZN(n83243) );
  AOI22_X1 U68814 ( .A1(n83244), .A2(n107799), .B1(n83126), .B2(n107787), .ZN(
        n83242) );
  NAND2_X1 U68815 ( .A1(n83245), .A2(n83246), .ZN(n83234) );
  AOI22_X1 U68816 ( .A1(n83135), .A2(n107820), .B1(n70239), .B2(n105875), .ZN(
        n83246) );
  AOI22_X1 U68817 ( .A1(n105874), .A2(n107804), .B1(n105873), .B2(n107807), 
        .ZN(n83245) );
  NOR4_X1 U68818 ( .A1(n83247), .A2(n83248), .A3(n83249), .A4(n83250), .ZN(
        n83232) );
  OAI21_X1 U68819 ( .B1(n103869), .B2(n83143), .A(n83251), .ZN(n83250) );
  NAND2_X1 U68821 ( .A1(n83252), .A2(n83253), .ZN(n83249) );
  AOI22_X1 U68822 ( .A1(n83149), .A2(n107834), .B1(n70147), .B2(n83150), .ZN(
        n83253) );
  AOI22_X1 U68823 ( .A1(n83151), .A2(n107837), .B1(n83152), .B2(n107776), .ZN(
        n83252) );
  OAI21_X1 U68824 ( .B1(n83254), .B2(n107832), .A(n83255), .ZN(n83248) );
  AOI22_X1 U68825 ( .A1(n70151), .A2(n83155), .B1(n83256), .B2(n107828), .ZN(
        n83255) );
  NAND2_X1 U68826 ( .A1(n83257), .A2(n83258), .ZN(n83247) );
  AOI22_X1 U68827 ( .A1(n105862), .A2(n107773), .B1(n105861), .B2(n107768), 
        .ZN(n83258) );
  AOI22_X1 U68828 ( .A1(n105860), .A2(n107764), .B1(n70159), .B2(n83154), .ZN(
        n83257) );
  NOR2_X1 U68829 ( .A1(n103867), .A2(n105858), .ZN(n83229) );
  AOI22_X1 U68830 ( .A1(n105856), .A2(n107770), .B1(n83165), .B2(n107815), 
        .ZN(n83227) );
  AOI22_X1 U68831 ( .A1(n105854), .A2(n107845), .B1(n106286), .B2(n107793), 
        .ZN(n83226) );
  AOI22_X1 U68832 ( .A1(n70187), .A2(n80260), .B1(n83259), .B2(n70258), .ZN(
        n83225) );
  NAND4_X2 U68833 ( .A1(n83260), .A2(n83261), .A3(n83262), .A4(n83263), .ZN(
        n58860) );
  NOR3_X1 U68834 ( .A1(n83264), .A2(n83265), .A3(n83266), .ZN(n83263) );
  AOI21_X1 U68836 ( .B1(n83267), .B2(n83268), .A(n106326), .ZN(n83265) );
  NOR4_X1 U68837 ( .A1(n83269), .A2(n83270), .A3(n83271), .A4(n83272), .ZN(
        n83268) );
  OAI21_X1 U68838 ( .B1(n103843), .B2(n106739), .A(n83273), .ZN(n83272) );
  AOI22_X1 U68839 ( .A1(n105884), .A2(n110680), .B1(n105883), .B2(n110684), 
        .ZN(n83273) );
  NAND2_X1 U68840 ( .A1(n83274), .A2(n83275), .ZN(n83271) );
  AOI22_X1 U68841 ( .A1(n105882), .A2(n110688), .B1(n74045), .B2(n105881), 
        .ZN(n83275) );
  AOI22_X1 U68842 ( .A1(n105880), .A2(n110719), .B1(n83129), .B2(n74033), .ZN(
        n83274) );
  OAI21_X1 U68843 ( .B1(n106738), .B2(n104651), .A(n83276), .ZN(n83270) );
  AOI22_X1 U68844 ( .A1(n74077), .A2(n105878), .B1(n74057), .B2(n105877), .ZN(
        n83276) );
  NAND2_X1 U68845 ( .A1(n83277), .A2(n83278), .ZN(n83269) );
  AOI22_X1 U68846 ( .A1(n83135), .A2(n110716), .B1(n74085), .B2(n105875), .ZN(
        n83278) );
  AOI22_X1 U68847 ( .A1(n74069), .A2(n105874), .B1(n105873), .B2(n110704), 
        .ZN(n83277) );
  NOR4_X1 U68848 ( .A1(n83279), .A2(n83280), .A3(n83281), .A4(n83282), .ZN(
        n83267) );
  OAI21_X1 U68849 ( .B1(n103851), .B2(n105872), .A(n83283), .ZN(n83282) );
  NAND2_X1 U68851 ( .A1(n83284), .A2(n83285), .ZN(n83281) );
  AOI22_X1 U68852 ( .A1(n83149), .A2(n110729), .B1(n73993), .B2(n83150), .ZN(
        n83285) );
  AOI22_X1 U68853 ( .A1(n83151), .A2(n110732), .B1(n83152), .B2(n110678), .ZN(
        n83284) );
  OAI21_X1 U68854 ( .B1(n103850), .B2(n106741), .A(n83286), .ZN(n83280) );
  AOI22_X1 U68855 ( .A1(n74005), .A2(n105866), .B1(n73997), .B2(n105865), .ZN(
        n83286) );
  NAND2_X1 U68856 ( .A1(n83287), .A2(n83288), .ZN(n83279) );
  AOI22_X1 U68857 ( .A1(n83158), .A2(n110693), .B1(n74021), .B2(n105862), .ZN(
        n83288) );
  AOI22_X1 U68858 ( .A1(n83160), .A2(n110671), .B1(n105860), .B2(n110667), 
        .ZN(n83287) );
  AND2_X2 U68859 ( .A1(n105859), .A2(n74104), .ZN(n83264) );
  AOI22_X1 U68860 ( .A1(n83163), .A2(n110660), .B1(n105856), .B2(n110673), 
        .ZN(n83262) );
  AOI22_X1 U68861 ( .A1(n105855), .A2(n110711), .B1(n105854), .B2(n110740), 
        .ZN(n83261) );
  AOI22_X1 U68862 ( .A1(n106287), .A2(n110693), .B1(n74033), .B2(n106285), 
        .ZN(n83260) );
  NAND4_X2 U68863 ( .A1(n83289), .A2(n83290), .A3(n83291), .A4(n83292), .ZN(
        n58859) );
  NOR3_X1 U68864 ( .A1(n83293), .A2(n83294), .A3(n83295), .ZN(n83292) );
  AOI21_X1 U68866 ( .B1(n83296), .B2(n83297), .A(n106325), .ZN(n83294) );
  NOR4_X1 U68867 ( .A1(n83298), .A2(n83299), .A3(n83300), .A4(n83301), .ZN(
        n83297) );
  OAI21_X1 U68868 ( .B1(n103829), .B2(n105864), .A(n83302), .ZN(n83301) );
  AOI22_X1 U68869 ( .A1(n105883), .A2(n108084), .B1(n83239), .B2(n108095), 
        .ZN(n83302) );
  NAND2_X1 U68870 ( .A1(n83303), .A2(n83304), .ZN(n83300) );
  AOI22_X1 U68871 ( .A1(n70632), .A2(n83127), .B1(n83128), .B2(n108122), .ZN(
        n83304) );
  AOI22_X1 U68872 ( .A1(n70620), .A2(n105879), .B1(n105884), .B2(n108080), 
        .ZN(n83303) );
  NAND2_X1 U68873 ( .A1(n83305), .A2(n83306), .ZN(n83299) );
  AOI22_X1 U68874 ( .A1(n70664), .A2(n105878), .B1(n105877), .B2(n108098), 
        .ZN(n83306) );
  AOI22_X1 U68875 ( .A1(n83244), .A2(n108101), .B1(n83126), .B2(n108088), .ZN(
        n83305) );
  NAND2_X1 U68876 ( .A1(n83307), .A2(n83308), .ZN(n83298) );
  AOI22_X1 U68877 ( .A1(n83135), .A2(n108119), .B1(n70672), .B2(n105875), .ZN(
        n83308) );
  AOI22_X1 U68878 ( .A1(n70656), .A2(n105874), .B1(n105873), .B2(n108107), 
        .ZN(n83307) );
  NOR4_X1 U68879 ( .A1(n83309), .A2(n83310), .A3(n83311), .A4(n83312), .ZN(
        n83296) );
  OAI21_X1 U68880 ( .B1(n103837), .B2(n83143), .A(n83313), .ZN(n83312) );
  NAND2_X1 U68882 ( .A1(n83314), .A2(n83315), .ZN(n83311) );
  AOI22_X1 U68883 ( .A1(n83149), .A2(n108134), .B1(n70580), .B2(n83150), .ZN(
        n83315) );
  AOI22_X1 U68884 ( .A1(n83151), .A2(n108137), .B1(n83152), .B2(n108078), .ZN(
        n83314) );
  OAI21_X1 U68885 ( .B1(n83254), .B2(n108132), .A(n83316), .ZN(n83310) );
  AOI22_X1 U68886 ( .A1(n70584), .A2(n83155), .B1(n83256), .B2(n108128), .ZN(
        n83316) );
  NAND2_X1 U68887 ( .A1(n83317), .A2(n83318), .ZN(n83309) );
  AOI22_X1 U68888 ( .A1(n105862), .A2(n108075), .B1(n105861), .B2(n108070), 
        .ZN(n83318) );
  AOI22_X1 U68889 ( .A1(n105860), .A2(n108066), .B1(n70592), .B2(n83154), .ZN(
        n83317) );
  NOR2_X1 U68890 ( .A1(n103835), .A2(n105858), .ZN(n83293) );
  AOI22_X1 U68891 ( .A1(n105856), .A2(n108072), .B1(n83165), .B2(n108114), 
        .ZN(n83291) );
  AOI22_X1 U68892 ( .A1(n105854), .A2(n108145), .B1(n106289), .B2(n108093), 
        .ZN(n83290) );
  AOI22_X1 U68893 ( .A1(n70620), .A2(n80260), .B1(n70691), .B2(n83259), .ZN(
        n83289) );
  NAND4_X2 U68894 ( .A1(n83319), .A2(n83320), .A3(n83321), .A4(n83322), .ZN(
        n58858) );
  NOR3_X1 U68895 ( .A1(n83323), .A2(n83324), .A3(n83325), .ZN(n83322) );
  AOI21_X1 U68897 ( .B1(n83326), .B2(n83327), .A(n106323), .ZN(n83324) );
  NOR4_X1 U68898 ( .A1(n83328), .A2(n83329), .A3(n83330), .A4(n83331), .ZN(
        n83327) );
  OAI21_X1 U68899 ( .B1(n103812), .B2(n105168), .A(n83332), .ZN(n83331) );
  AOI22_X1 U68900 ( .A1(n105884), .A2(n110777), .B1(n105883), .B2(n110782), 
        .ZN(n83332) );
  NAND2_X1 U68901 ( .A1(n83333), .A2(n83334), .ZN(n83330) );
  AOI22_X1 U68902 ( .A1(n105882), .A2(n110786), .B1(n74186), .B2(n105881), 
        .ZN(n83334) );
  AOI22_X1 U68903 ( .A1(n105880), .A2(n110821), .B1(n74174), .B2(n105879), 
        .ZN(n83333) );
  OAI21_X1 U68904 ( .B1(n100997), .B2(n105167), .A(n83335), .ZN(n83329) );
  AOI22_X1 U68905 ( .A1(n74218), .A2(n105878), .B1(n105877), .B2(n110797), 
        .ZN(n83335) );
  NAND2_X1 U68906 ( .A1(n83336), .A2(n83337), .ZN(n83328) );
  AOI22_X1 U68907 ( .A1(n83135), .A2(n110818), .B1(n74226), .B2(n105875), .ZN(
        n83337) );
  AOI22_X1 U68908 ( .A1(n74210), .A2(n105874), .B1(n105873), .B2(n110806), 
        .ZN(n83336) );
  NOR4_X1 U68909 ( .A1(n83338), .A2(n83339), .A3(n83340), .A4(n83341), .ZN(
        n83326) );
  OAI21_X1 U68910 ( .B1(n103821), .B2(n105872), .A(n83342), .ZN(n83341) );
  NAND2_X1 U68912 ( .A1(n83343), .A2(n83344), .ZN(n83340) );
  AOI22_X1 U68913 ( .A1(n83149), .A2(n110832), .B1(n74134), .B2(n83150), .ZN(
        n83344) );
  AOI22_X1 U68914 ( .A1(n83151), .A2(n110835), .B1(n83152), .B2(n110775), .ZN(
        n83343) );
  OAI21_X1 U68915 ( .B1(n103820), .B2(n106741), .A(n83345), .ZN(n83339) );
  AOI22_X1 U68916 ( .A1(n74146), .A2(n105866), .B1(n105865), .B2(n74138), .ZN(
        n83345) );
  NAND2_X1 U68917 ( .A1(n83346), .A2(n83347), .ZN(n83338) );
  AOI22_X1 U68918 ( .A1(n83158), .A2(n110792), .B1(n105862), .B2(n74162), .ZN(
        n83347) );
  AOI22_X1 U68919 ( .A1(n83160), .A2(n110768), .B1(n105860), .B2(n110764), 
        .ZN(n83346) );
  AND2_X2 U68920 ( .A1(n105859), .A2(n74245), .ZN(n83323) );
  AOI22_X1 U68921 ( .A1(n83163), .A2(n110757), .B1(n105856), .B2(n110770), 
        .ZN(n83321) );
  AOI22_X1 U68922 ( .A1(n105855), .A2(n110813), .B1(n105854), .B2(n110843), 
        .ZN(n83320) );
  AOI22_X1 U68923 ( .A1(n106287), .A2(n110792), .B1(n74174), .B2(n106284), 
        .ZN(n83319) );
  NAND4_X2 U68924 ( .A1(n83348), .A2(n83349), .A3(n83350), .A4(n83351), .ZN(
        n58857) );
  NOR3_X1 U68925 ( .A1(n83352), .A2(n83353), .A3(n83354), .ZN(n83351) );
  NOR2_X1 U68926 ( .A1(n103793), .A2(n106737), .ZN(n83354) );
  AOI21_X1 U68927 ( .B1(n83355), .B2(n83356), .A(n106324), .ZN(n83353) );
  NOR4_X1 U68928 ( .A1(n83357), .A2(n83358), .A3(n83359), .A4(n83360), .ZN(
        n83356) );
  OAI21_X1 U68929 ( .B1(n103796), .B2(n105168), .A(n83361), .ZN(n83360) );
  AOI22_X1 U68930 ( .A1(n105884), .A2(n110878), .B1(n105883), .B2(n110883), 
        .ZN(n83361) );
  NAND2_X1 U68931 ( .A1(n83362), .A2(n83363), .ZN(n83359) );
  AOI22_X1 U68932 ( .A1(n105882), .A2(n110886), .B1(n74326), .B2(n105881), 
        .ZN(n83363) );
  AOI22_X1 U68933 ( .A1(n105880), .A2(n110922), .B1(n74314), .B2(n105879), 
        .ZN(n83362) );
  OAI21_X1 U68934 ( .B1(n105167), .B2(n104650), .A(n83364), .ZN(n83358) );
  AOI22_X1 U68935 ( .A1(n105878), .A2(n110909), .B1(n74338), .B2(n105877), 
        .ZN(n83364) );
  NAND2_X1 U68936 ( .A1(n83365), .A2(n83366), .ZN(n83357) );
  AOI22_X1 U68937 ( .A1(n83135), .A2(n110919), .B1(n74366), .B2(n105875), .ZN(
        n83366) );
  AOI22_X1 U68938 ( .A1(n105874), .A2(n110901), .B1(n105873), .B2(n110905), 
        .ZN(n83365) );
  NOR4_X1 U68939 ( .A1(n83367), .A2(n83368), .A3(n83369), .A4(n83370), .ZN(
        n83355) );
  OAI21_X1 U68940 ( .B1(n103805), .B2(n83143), .A(n83371), .ZN(n83370) );
  NAND2_X1 U68942 ( .A1(n83372), .A2(n83373), .ZN(n83369) );
  AOI22_X1 U68943 ( .A1(n83149), .A2(n110933), .B1(n74274), .B2(n83150), .ZN(
        n83373) );
  AOI22_X1 U68944 ( .A1(n83151), .A2(n110936), .B1(n83152), .B2(n110876), .ZN(
        n83372) );
  OAI21_X1 U68945 ( .B1(n103804), .B2(n106741), .A(n83374), .ZN(n83368) );
  AOI22_X1 U68946 ( .A1(n74286), .A2(n105866), .B1(n74278), .B2(n105865), .ZN(
        n83374) );
  NAND2_X1 U68947 ( .A1(n83375), .A2(n83376), .ZN(n83367) );
  AOI22_X1 U68948 ( .A1(n83158), .A2(n111016), .B1(n74302), .B2(n105862), .ZN(
        n83376) );
  AOI22_X1 U68949 ( .A1(n83160), .A2(n110869), .B1(n105860), .B2(n110865), 
        .ZN(n83375) );
  AOI22_X1 U68951 ( .A1(n83163), .A2(n110858), .B1(n105856), .B2(n110871), 
        .ZN(n83350) );
  AOI22_X1 U68952 ( .A1(n105855), .A2(n110913), .B1(n105854), .B2(n110944), 
        .ZN(n83349) );
  AOI22_X1 U68953 ( .A1(n106288), .A2(n111016), .B1(n74314), .B2(n106284), 
        .ZN(n83348) );
  NAND4_X2 U68954 ( .A1(n83377), .A2(n83378), .A3(n83379), .A4(n83380), .ZN(
        n58856) );
  NOR3_X1 U68955 ( .A1(n83381), .A2(n83382), .A3(n83383), .ZN(n83380) );
  NOR2_X1 U68956 ( .A1(n103776), .A2(n106737), .ZN(n83383) );
  AOI21_X1 U68957 ( .B1(n83384), .B2(n83385), .A(n106325), .ZN(n83382) );
  NOR4_X1 U68958 ( .A1(n83386), .A2(n83387), .A3(n83388), .A4(n83389), .ZN(
        n83385) );
  OAI21_X1 U68959 ( .B1(n103780), .B2(n105168), .A(n83390), .ZN(n83389) );
  AOI22_X1 U68960 ( .A1(n105884), .A2(n110472), .B1(n105883), .B2(n110477), 
        .ZN(n83390) );
  NAND2_X1 U68961 ( .A1(n83391), .A2(n83392), .ZN(n83388) );
  AOI22_X1 U68962 ( .A1(n105882), .A2(n110480), .B1(n73762), .B2(n105881), 
        .ZN(n83392) );
  AOI22_X1 U68963 ( .A1(n105880), .A2(n110516), .B1(n73750), .B2(n105879), 
        .ZN(n83391) );
  OAI21_X1 U68964 ( .B1(n100998), .B2(n105167), .A(n83393), .ZN(n83387) );
  AOI22_X1 U68965 ( .A1(n105878), .A2(n110504), .B1(n105877), .B2(n110490), 
        .ZN(n83393) );
  NAND2_X1 U68966 ( .A1(n83394), .A2(n83395), .ZN(n83386) );
  AOI22_X1 U68967 ( .A1(n83135), .A2(n110513), .B1(n73802), .B2(n105875), .ZN(
        n83395) );
  AOI22_X1 U68968 ( .A1(n105874), .A2(n110496), .B1(n105873), .B2(n110500), 
        .ZN(n83394) );
  NOR4_X1 U68969 ( .A1(n83396), .A2(n83397), .A3(n83398), .A4(n83399), .ZN(
        n83384) );
  OAI21_X1 U68970 ( .B1(n103788), .B2(n105872), .A(n83400), .ZN(n83399) );
  NAND2_X1 U68972 ( .A1(n83401), .A2(n83402), .ZN(n83398) );
  AOI22_X1 U68973 ( .A1(n83149), .A2(n110526), .B1(n73710), .B2(n83150), .ZN(
        n83402) );
  AOI22_X1 U68974 ( .A1(n83151), .A2(n110529), .B1(n83152), .B2(n110471), .ZN(
        n83401) );
  OAI21_X1 U68975 ( .B1(n103787), .B2(n106741), .A(n83403), .ZN(n83397) );
  AOI22_X1 U68976 ( .A1(n73722), .A2(n105866), .B1(n73714), .B2(n105865), .ZN(
        n83403) );
  NAND2_X1 U68977 ( .A1(n83404), .A2(n83405), .ZN(n83396) );
  AOI22_X1 U68978 ( .A1(n83158), .A2(n111017), .B1(n73738), .B2(n105862), .ZN(
        n83405) );
  AOI22_X1 U68979 ( .A1(n83160), .A2(n110464), .B1(n105860), .B2(n110460), 
        .ZN(n83404) );
  AOI22_X1 U68981 ( .A1(n83163), .A2(n110453), .B1(n105856), .B2(n110466), 
        .ZN(n83379) );
  AOI22_X1 U68982 ( .A1(n105855), .A2(n110508), .B1(n105854), .B2(n110537), 
        .ZN(n83378) );
  AOI22_X1 U68983 ( .A1(n106288), .A2(n111017), .B1(n73750), .B2(n106282), 
        .ZN(n83377) );
  NAND4_X2 U68984 ( .A1(n83406), .A2(n83407), .A3(n83408), .A4(n83409), .ZN(
        n58855) );
  NOR3_X1 U68985 ( .A1(n83410), .A2(n83411), .A3(n83412), .ZN(n83409) );
  NOR2_X1 U68986 ( .A1(n103759), .A2(n106737), .ZN(n83412) );
  AOI21_X1 U68987 ( .B1(n83413), .B2(n83414), .A(n106327), .ZN(n83411) );
  NOR4_X1 U68988 ( .A1(n83415), .A2(n83416), .A3(n83417), .A4(n83418), .ZN(
        n83414) );
  OAI21_X1 U68989 ( .B1(n103763), .B2(n105168), .A(n83419), .ZN(n83418) );
  AOI22_X1 U68990 ( .A1(n105884), .A2(n110254), .B1(n105883), .B2(n110259), 
        .ZN(n83419) );
  NAND2_X1 U68991 ( .A1(n83420), .A2(n83421), .ZN(n83417) );
  AOI22_X1 U68992 ( .A1(n105882), .A2(n110262), .B1(n73466), .B2(n105881), 
        .ZN(n83421) );
  AOI22_X1 U68993 ( .A1(n105880), .A2(n110300), .B1(n83129), .B2(n73454), .ZN(
        n83420) );
  OAI21_X1 U68994 ( .B1(n100999), .B2(n106738), .A(n83422), .ZN(n83416) );
  AOI22_X1 U68995 ( .A1(n105878), .A2(n110287), .B1(n105877), .B2(n110273), 
        .ZN(n83422) );
  NAND2_X1 U68996 ( .A1(n83423), .A2(n83424), .ZN(n83415) );
  AOI22_X1 U68997 ( .A1(n83135), .A2(n110297), .B1(n73506), .B2(n105875), .ZN(
        n83424) );
  AOI22_X1 U68998 ( .A1(n105874), .A2(n111039), .B1(n105873), .B2(n110283), 
        .ZN(n83423) );
  NOR4_X1 U68999 ( .A1(n83425), .A2(n83426), .A3(n83427), .A4(n83428), .ZN(
        n83413) );
  OAI21_X1 U69000 ( .B1(n103771), .B2(n105872), .A(n83429), .ZN(n83428) );
  NAND2_X1 U69002 ( .A1(n83430), .A2(n83431), .ZN(n83427) );
  AOI22_X1 U69003 ( .A1(n83149), .A2(n110311), .B1(n73414), .B2(n83150), .ZN(
        n83431) );
  AOI22_X1 U69004 ( .A1(n83151), .A2(n110314), .B1(n83152), .B2(n110253), .ZN(
        n83430) );
  OAI21_X1 U69005 ( .B1(n103770), .B2(n106741), .A(n83432), .ZN(n83426) );
  AOI22_X1 U69006 ( .A1(n73426), .A2(n105866), .B1(n73418), .B2(n105865), .ZN(
        n83432) );
  NAND2_X1 U69007 ( .A1(n83433), .A2(n83434), .ZN(n83425) );
  AOI22_X1 U69008 ( .A1(n83158), .A2(n110268), .B1(n73442), .B2(n105862), .ZN(
        n83434) );
  AOI22_X1 U69009 ( .A1(n83160), .A2(n110246), .B1(n105860), .B2(n110242), 
        .ZN(n83433) );
  AOI22_X1 U69011 ( .A1(n83163), .A2(n110235), .B1(n105856), .B2(n110248), 
        .ZN(n83408) );
  AOI22_X1 U69012 ( .A1(n105855), .A2(n110291), .B1(n105854), .B2(n110322), 
        .ZN(n83407) );
  AOI22_X1 U69013 ( .A1(n106289), .A2(n110268), .B1(n73454), .B2(n106283), 
        .ZN(n83406) );
  NAND4_X2 U69014 ( .A1(n83435), .A2(n83436), .A3(n83437), .A4(n83438), .ZN(
        n58854) );
  NOR3_X1 U69015 ( .A1(n83439), .A2(n83440), .A3(n83441), .ZN(n83438) );
  NOR2_X1 U69016 ( .A1(n103742), .A2(n106737), .ZN(n83441) );
  AOI21_X1 U69017 ( .B1(n83442), .B2(n83443), .A(n106327), .ZN(n83440) );
  NOR4_X1 U69018 ( .A1(n83444), .A2(n83445), .A3(n83446), .A4(n83447), .ZN(
        n83443) );
  OAI21_X1 U69019 ( .B1(n103746), .B2(n105168), .A(n83448), .ZN(n83447) );
  AOI22_X1 U69020 ( .A1(n105884), .A2(n110571), .B1(n105883), .B2(n110576), 
        .ZN(n83448) );
  NAND2_X1 U69021 ( .A1(n83449), .A2(n83450), .ZN(n83446) );
  AOI22_X1 U69022 ( .A1(n105882), .A2(n110580), .B1(n73903), .B2(n105881), 
        .ZN(n83450) );
  AOI22_X1 U69023 ( .A1(n105880), .A2(n110621), .B1(n73891), .B2(n105879), 
        .ZN(n83449) );
  OAI21_X1 U69024 ( .B1(n101000), .B2(n105167), .A(n83451), .ZN(n83445) );
  AOI22_X1 U69025 ( .A1(n105878), .A2(n110607), .B1(n105877), .B2(n110591), 
        .ZN(n83451) );
  NAND2_X1 U69026 ( .A1(n83452), .A2(n83453), .ZN(n83444) );
  AOI22_X1 U69027 ( .A1(n83135), .A2(n110617), .B1(n73943), .B2(n105875), .ZN(
        n83453) );
  AOI22_X1 U69028 ( .A1(n105874), .A2(n110599), .B1(n105873), .B2(n110603), 
        .ZN(n83452) );
  NOR4_X1 U69029 ( .A1(n83454), .A2(n83455), .A3(n83456), .A4(n83457), .ZN(
        n83442) );
  OAI21_X1 U69030 ( .B1(n103754), .B2(n105872), .A(n83458), .ZN(n83457) );
  NAND2_X1 U69032 ( .A1(n83459), .A2(n83460), .ZN(n83456) );
  AOI22_X1 U69033 ( .A1(n83149), .A2(n110631), .B1(n73851), .B2(n83150), .ZN(
        n83460) );
  AOI22_X1 U69034 ( .A1(n83151), .A2(n110634), .B1(n83152), .B2(n110570), .ZN(
        n83459) );
  OAI21_X1 U69035 ( .B1(n103753), .B2(n106741), .A(n83461), .ZN(n83455) );
  AOI22_X1 U69036 ( .A1(n73863), .A2(n105866), .B1(n73855), .B2(n105865), .ZN(
        n83461) );
  NAND2_X1 U69037 ( .A1(n83462), .A2(n83463), .ZN(n83454) );
  AOI22_X1 U69038 ( .A1(n83158), .A2(n110586), .B1(n73879), .B2(n105862), .ZN(
        n83463) );
  AOI22_X1 U69039 ( .A1(n83160), .A2(n110563), .B1(n105860), .B2(n110559), 
        .ZN(n83462) );
  AOI22_X1 U69041 ( .A1(n83163), .A2(n110552), .B1(n105856), .B2(n110565), 
        .ZN(n83437) );
  AOI22_X1 U69042 ( .A1(n105855), .A2(n110611), .B1(n105854), .B2(n110642), 
        .ZN(n83436) );
  AOI22_X1 U69043 ( .A1(n106288), .A2(n110586), .B1(n73891), .B2(n106284), 
        .ZN(n83435) );
  NAND4_X2 U69044 ( .A1(n83464), .A2(n83465), .A3(n83466), .A4(n83467), .ZN(
        n58853) );
  NOR3_X1 U69045 ( .A1(n83468), .A2(n83469), .A3(n83470), .ZN(n83467) );
  NOR2_X1 U69046 ( .A1(n103726), .A2(n106737), .ZN(n83470) );
  AOI21_X1 U69047 ( .B1(n83471), .B2(n83472), .A(n106327), .ZN(n83469) );
  NOR4_X1 U69048 ( .A1(n83473), .A2(n83474), .A3(n83475), .A4(n83476), .ZN(
        n83472) );
  OAI21_X1 U69049 ( .B1(n103729), .B2(n105168), .A(n83477), .ZN(n83476) );
  AOI22_X1 U69050 ( .A1(n105884), .A2(n110362), .B1(n105883), .B2(n110367), 
        .ZN(n83477) );
  NAND2_X1 U69051 ( .A1(n83478), .A2(n83479), .ZN(n83475) );
  AOI22_X1 U69052 ( .A1(n105882), .A2(n110371), .B1(n73615), .B2(n105881), 
        .ZN(n83479) );
  AOI22_X1 U69053 ( .A1(n105880), .A2(n110409), .B1(n83129), .B2(n73603), .ZN(
        n83478) );
  OAI21_X1 U69054 ( .B1(n101001), .B2(n106738), .A(n83480), .ZN(n83474) );
  AOI22_X1 U69055 ( .A1(n105878), .A2(n110396), .B1(n73627), .B2(n105877), 
        .ZN(n83480) );
  NAND2_X1 U69056 ( .A1(n83481), .A2(n83482), .ZN(n83473) );
  AOI22_X1 U69057 ( .A1(n105876), .A2(n110406), .B1(n73655), .B2(n105875), 
        .ZN(n83482) );
  AOI22_X1 U69058 ( .A1(n105874), .A2(n111038), .B1(n105873), .B2(n110392), 
        .ZN(n83481) );
  NOR4_X1 U69059 ( .A1(n83483), .A2(n83484), .A3(n83485), .A4(n83486), .ZN(
        n83471) );
  OAI21_X1 U69060 ( .B1(n103737), .B2(n105872), .A(n83487), .ZN(n83486) );
  NAND2_X1 U69062 ( .A1(n83488), .A2(n83489), .ZN(n83485) );
  AOI22_X1 U69063 ( .A1(n105870), .A2(n110420), .B1(n73563), .B2(n105869), 
        .ZN(n83489) );
  AOI22_X1 U69064 ( .A1(n105868), .A2(n110423), .B1(n83152), .B2(n110361), 
        .ZN(n83488) );
  OAI21_X1 U69065 ( .B1(n103736), .B2(n106741), .A(n83490), .ZN(n83484) );
  AOI22_X1 U69066 ( .A1(n73575), .A2(n105866), .B1(n73567), .B2(n105865), .ZN(
        n83490) );
  NAND2_X1 U69067 ( .A1(n83491), .A2(n83492), .ZN(n83483) );
  AOI22_X1 U69068 ( .A1(n83158), .A2(n110377), .B1(n73591), .B2(n105862), .ZN(
        n83492) );
  AOI22_X1 U69069 ( .A1(n83160), .A2(n110354), .B1(n105860), .B2(n110350), 
        .ZN(n83491) );
  AND2_X2 U69070 ( .A1(n105859), .A2(n73674), .ZN(n83468) );
  AOI22_X1 U69071 ( .A1(n83163), .A2(n110343), .B1(n105856), .B2(n110356), 
        .ZN(n83466) );
  AOI22_X1 U69072 ( .A1(n105855), .A2(n110400), .B1(n105854), .B2(n110431), 
        .ZN(n83465) );
  AOI22_X1 U69073 ( .A1(n106286), .A2(n110377), .B1(n73603), .B2(n106285), 
        .ZN(n83464) );
  NAND4_X2 U69074 ( .A1(n83493), .A2(n83494), .A3(n83495), .A4(n83496), .ZN(
        n58852) );
  NOR3_X1 U69075 ( .A1(n83497), .A2(n83498), .A3(n83499), .ZN(n83496) );
  NOR2_X1 U69076 ( .A1(n103708), .A2(n106737), .ZN(n83499) );
  AOI21_X1 U69077 ( .B1(n83500), .B2(n83501), .A(n106327), .ZN(n83498) );
  NOR4_X1 U69078 ( .A1(n83502), .A2(n83503), .A3(n83504), .A4(n83505), .ZN(
        n83501) );
  OAI21_X1 U69079 ( .B1(n103712), .B2(n105168), .A(n83506), .ZN(n83505) );
  AOI22_X1 U69080 ( .A1(n83122), .A2(n110038), .B1(n105883), .B2(n110043), 
        .ZN(n83506) );
  NAND2_X1 U69081 ( .A1(n83507), .A2(n83508), .ZN(n83504) );
  AOI22_X1 U69082 ( .A1(n105882), .A2(n110047), .B1(n73177), .B2(n105881), 
        .ZN(n83508) );
  AOI22_X1 U69083 ( .A1(n105880), .A2(n110087), .B1(n83129), .B2(n73165), .ZN(
        n83507) );
  OAI21_X1 U69084 ( .B1(n101002), .B2(n105167), .A(n83509), .ZN(n83503) );
  AOI22_X1 U69085 ( .A1(n105878), .A2(n110074), .B1(n105877), .B2(n110059), 
        .ZN(n83509) );
  NAND2_X1 U69086 ( .A1(n83510), .A2(n83511), .ZN(n83502) );
  AOI22_X1 U69087 ( .A1(n105876), .A2(n110084), .B1(n73217), .B2(n105875), 
        .ZN(n83511) );
  AOI22_X1 U69088 ( .A1(n105874), .A2(n111040), .B1(n105873), .B2(n110070), 
        .ZN(n83510) );
  NOR4_X1 U69089 ( .A1(n83512), .A2(n83513), .A3(n83514), .A4(n83515), .ZN(
        n83500) );
  OAI21_X1 U69090 ( .B1(n103721), .B2(n105872), .A(n83516), .ZN(n83515) );
  NAND2_X1 U69092 ( .A1(n83517), .A2(n83518), .ZN(n83514) );
  AOI22_X1 U69093 ( .A1(n105870), .A2(n110098), .B1(n73125), .B2(n105869), 
        .ZN(n83518) );
  AOI22_X1 U69094 ( .A1(n105868), .A2(n110101), .B1(n105867), .B2(n110037), 
        .ZN(n83517) );
  OAI21_X1 U69095 ( .B1(n103720), .B2(n106741), .A(n83519), .ZN(n83513) );
  AOI22_X1 U69096 ( .A1(n73137), .A2(n105866), .B1(n73129), .B2(n105865), .ZN(
        n83519) );
  NAND2_X1 U69097 ( .A1(n83520), .A2(n83521), .ZN(n83512) );
  AOI22_X1 U69098 ( .A1(n83158), .A2(n110053), .B1(n105862), .B2(n110034), 
        .ZN(n83521) );
  AOI22_X1 U69099 ( .A1(n83160), .A2(n110029), .B1(n105860), .B2(n110025), 
        .ZN(n83520) );
  AOI22_X1 U69101 ( .A1(n83163), .A2(n110018), .B1(n105856), .B2(n110031), 
        .ZN(n83495) );
  AOI22_X1 U69102 ( .A1(n105855), .A2(n110078), .B1(n105854), .B2(n110109), 
        .ZN(n83494) );
  AOI22_X1 U69103 ( .A1(n106287), .A2(n110053), .B1(n73165), .B2(n106284), 
        .ZN(n83493) );
  NAND4_X2 U69104 ( .A1(n83522), .A2(n83523), .A3(n83524), .A4(n83525), .ZN(
        n58851) );
  NOR3_X1 U69105 ( .A1(n83526), .A2(n83527), .A3(n83528), .ZN(n83525) );
  NOR2_X1 U69106 ( .A1(n103691), .A2(n106737), .ZN(n83528) );
  AOI21_X1 U69107 ( .B1(n83529), .B2(n83530), .A(n106327), .ZN(n83527) );
  NOR4_X1 U69108 ( .A1(n83531), .A2(n83532), .A3(n83533), .A4(n83534), .ZN(
        n83530) );
  OAI21_X1 U69109 ( .B1(n103695), .B2(n105168), .A(n83535), .ZN(n83534) );
  AOI22_X1 U69110 ( .A1(n83122), .A2(n110145), .B1(n105883), .B2(n110150), 
        .ZN(n83535) );
  NAND2_X1 U69111 ( .A1(n83536), .A2(n83537), .ZN(n83533) );
  AOI22_X1 U69112 ( .A1(n105882), .A2(n110154), .B1(n73319), .B2(n83127), .ZN(
        n83537) );
  AOI22_X1 U69113 ( .A1(n105880), .A2(n110194), .B1(n73307), .B2(n105879), 
        .ZN(n83536) );
  OAI21_X1 U69114 ( .B1(n101003), .B2(n106738), .A(n83538), .ZN(n83532) );
  AOI22_X1 U69115 ( .A1(n105878), .A2(n110181), .B1(n105877), .B2(n110166), 
        .ZN(n83538) );
  NAND2_X1 U69116 ( .A1(n83539), .A2(n83540), .ZN(n83531) );
  AOI22_X1 U69117 ( .A1(n105876), .A2(n110191), .B1(n73359), .B2(n105875), 
        .ZN(n83540) );
  AOI22_X1 U69118 ( .A1(n105874), .A2(n111035), .B1(n105873), .B2(n110177), 
        .ZN(n83539) );
  NOR4_X1 U69119 ( .A1(n83541), .A2(n83542), .A3(n83543), .A4(n83544), .ZN(
        n83529) );
  OAI21_X1 U69120 ( .B1(n103704), .B2(n105872), .A(n83545), .ZN(n83544) );
  NAND2_X1 U69122 ( .A1(n83546), .A2(n83547), .ZN(n83543) );
  AOI22_X1 U69123 ( .A1(n105870), .A2(n110205), .B1(n73267), .B2(n105869), 
        .ZN(n83547) );
  AOI22_X1 U69124 ( .A1(n105868), .A2(n110208), .B1(n105867), .B2(n110144), 
        .ZN(n83546) );
  OAI21_X1 U69125 ( .B1(n103703), .B2(n106741), .A(n83548), .ZN(n83542) );
  AOI22_X1 U69126 ( .A1(n73279), .A2(n105866), .B1(n73271), .B2(n83155), .ZN(
        n83548) );
  NAND2_X1 U69127 ( .A1(n83549), .A2(n83550), .ZN(n83541) );
  AOI22_X1 U69128 ( .A1(n105863), .A2(n110160), .B1(n105862), .B2(n110141), 
        .ZN(n83550) );
  AOI22_X1 U69129 ( .A1(n83160), .A2(n110136), .B1(n105860), .B2(n110132), 
        .ZN(n83549) );
  AND2_X2 U69130 ( .A1(n105859), .A2(n73378), .ZN(n83526) );
  AOI22_X1 U69131 ( .A1(n105857), .A2(n110125), .B1(n105856), .B2(n110138), 
        .ZN(n83524) );
  AOI22_X1 U69132 ( .A1(n105855), .A2(n110185), .B1(n105854), .B2(n110216), 
        .ZN(n83523) );
  AOI22_X1 U69133 ( .A1(n106289), .A2(n110160), .B1(n73307), .B2(n106283), 
        .ZN(n83522) );
  NAND4_X2 U69134 ( .A1(n83551), .A2(n83552), .A3(n83553), .A4(n83554), .ZN(
        n58850) );
  NOR3_X1 U69135 ( .A1(n83555), .A2(n83556), .A3(n83557), .ZN(n83554) );
  NOR2_X1 U69136 ( .A1(n103673), .A2(n106737), .ZN(n83557) );
  AOI21_X1 U69137 ( .B1(n83558), .B2(n83559), .A(n106327), .ZN(n83556) );
  NOR4_X1 U69138 ( .A1(n83560), .A2(n83561), .A3(n83562), .A4(n83563), .ZN(
        n83559) );
  OAI21_X1 U69139 ( .B1(n103677), .B2(n105168), .A(n83564), .ZN(n83563) );
  AOI22_X1 U69140 ( .A1(n105884), .A2(n109929), .B1(n105883), .B2(n109934), 
        .ZN(n83564) );
  NAND2_X1 U69141 ( .A1(n83565), .A2(n83566), .ZN(n83562) );
  AOI22_X1 U69142 ( .A1(n105882), .A2(n109938), .B1(n73035), .B2(n105881), 
        .ZN(n83566) );
  AOI22_X1 U69143 ( .A1(n105880), .A2(n109979), .B1(n73023), .B2(n105879), 
        .ZN(n83565) );
  OAI21_X1 U69144 ( .B1(n101004), .B2(n105167), .A(n83567), .ZN(n83561) );
  AOI22_X1 U69145 ( .A1(n105878), .A2(n109966), .B1(n105877), .B2(n109950), 
        .ZN(n83567) );
  NAND2_X1 U69146 ( .A1(n83568), .A2(n83569), .ZN(n83560) );
  AOI22_X1 U69147 ( .A1(n105876), .A2(n109976), .B1(n73075), .B2(n105875), 
        .ZN(n83569) );
  AOI22_X1 U69148 ( .A1(n105874), .A2(n109958), .B1(n105873), .B2(n109962), 
        .ZN(n83568) );
  NOR4_X1 U69149 ( .A1(n83570), .A2(n83571), .A3(n83572), .A4(n83573), .ZN(
        n83558) );
  OAI21_X1 U69150 ( .B1(n103687), .B2(n105872), .A(n83574), .ZN(n83573) );
  NAND2_X1 U69152 ( .A1(n83575), .A2(n83576), .ZN(n83572) );
  AOI22_X1 U69153 ( .A1(n105870), .A2(n109990), .B1(n72983), .B2(n105869), 
        .ZN(n83576) );
  AOI22_X1 U69154 ( .A1(n105868), .A2(n109993), .B1(n105867), .B2(n109928), 
        .ZN(n83575) );
  OAI21_X1 U69155 ( .B1(n103685), .B2(n105169), .A(n83577), .ZN(n83571) );
  AOI22_X1 U69156 ( .A1(n72995), .A2(n105866), .B1(n72987), .B2(n105865), .ZN(
        n83577) );
  NAND2_X1 U69157 ( .A1(n83578), .A2(n83579), .ZN(n83570) );
  AOI22_X1 U69158 ( .A1(n105863), .A2(n109944), .B1(n105862), .B2(n109925), 
        .ZN(n83579) );
  AOI22_X1 U69159 ( .A1(n105861), .A2(n109920), .B1(n105860), .B2(n109916), 
        .ZN(n83578) );
  AOI22_X1 U69161 ( .A1(n105857), .A2(n109909), .B1(n105856), .B2(n109922), 
        .ZN(n83553) );
  AOI22_X1 U69162 ( .A1(n105855), .A2(n109970), .B1(n105854), .B2(n110001), 
        .ZN(n83552) );
  AOI22_X1 U69163 ( .A1(n106288), .A2(n109944), .B1(n73023), .B2(n106285), 
        .ZN(n83551) );
  NAND4_X2 U69164 ( .A1(n83580), .A2(n83581), .A3(n83582), .A4(n83583), .ZN(
        n58849) );
  NOR3_X1 U69165 ( .A1(n83584), .A2(n83585), .A3(n83586), .ZN(n83583) );
  NOR2_X1 U69166 ( .A1(n103655), .A2(n106737), .ZN(n83586) );
  AOI21_X1 U69167 ( .B1(n83587), .B2(n83588), .A(n106327), .ZN(n83585) );
  NOR4_X1 U69168 ( .A1(n83589), .A2(n83590), .A3(n83591), .A4(n83592), .ZN(
        n83588) );
  OAI21_X1 U69169 ( .B1(n103659), .B2(n105168), .A(n83593), .ZN(n83592) );
  AOI22_X1 U69170 ( .A1(n83122), .A2(n109812), .B1(n105883), .B2(n109817), 
        .ZN(n83593) );
  NAND2_X1 U69171 ( .A1(n83594), .A2(n83595), .ZN(n83591) );
  AOI22_X1 U69172 ( .A1(n105882), .A2(n109821), .B1(n72885), .B2(n83127), .ZN(
        n83595) );
  AOI22_X1 U69173 ( .A1(n105880), .A2(n109862), .B1(n72873), .B2(n105879), 
        .ZN(n83594) );
  OAI21_X1 U69174 ( .B1(n101005), .B2(n106738), .A(n83596), .ZN(n83590) );
  AOI22_X1 U69175 ( .A1(n105878), .A2(n109849), .B1(n105877), .B2(n109833), 
        .ZN(n83596) );
  NAND2_X1 U69176 ( .A1(n83597), .A2(n83598), .ZN(n83589) );
  AOI22_X1 U69177 ( .A1(n105876), .A2(n109859), .B1(n72925), .B2(n105875), 
        .ZN(n83598) );
  AOI22_X1 U69178 ( .A1(n105874), .A2(n109841), .B1(n105873), .B2(n109845), 
        .ZN(n83597) );
  NOR4_X1 U69179 ( .A1(n83599), .A2(n83600), .A3(n83601), .A4(n83602), .ZN(
        n83587) );
  OAI21_X1 U69180 ( .B1(n103669), .B2(n105872), .A(n83603), .ZN(n83602) );
  NAND2_X1 U69182 ( .A1(n83604), .A2(n83605), .ZN(n83601) );
  AOI22_X1 U69183 ( .A1(n105870), .A2(n109873), .B1(n72833), .B2(n105869), 
        .ZN(n83605) );
  AOI22_X1 U69184 ( .A1(n105868), .A2(n109876), .B1(n105867), .B2(n109810), 
        .ZN(n83604) );
  OAI21_X1 U69185 ( .B1(n103667), .B2(n106741), .A(n83606), .ZN(n83600) );
  AOI22_X1 U69186 ( .A1(n72845), .A2(n105866), .B1(n72837), .B2(n83155), .ZN(
        n83606) );
  NAND2_X1 U69187 ( .A1(n83607), .A2(n83608), .ZN(n83599) );
  AOI22_X1 U69188 ( .A1(n105863), .A2(n109827), .B1(n105862), .B2(n109807), 
        .ZN(n83608) );
  AOI22_X1 U69189 ( .A1(n105861), .A2(n109802), .B1(n105860), .B2(n109798), 
        .ZN(n83607) );
  AND2_X2 U69190 ( .A1(n105859), .A2(n72944), .ZN(n83584) );
  AOI22_X1 U69191 ( .A1(n105857), .A2(n109791), .B1(n105856), .B2(n109804), 
        .ZN(n83582) );
  AOI22_X1 U69192 ( .A1(n105855), .A2(n109853), .B1(n105854), .B2(n109884), 
        .ZN(n83581) );
  AOI22_X1 U69193 ( .A1(n106289), .A2(n109827), .B1(n72873), .B2(n106282), 
        .ZN(n83580) );
  NAND4_X2 U69194 ( .A1(n83609), .A2(n83610), .A3(n83611), .A4(n83612), .ZN(
        n58848) );
  NOR3_X1 U69195 ( .A1(n83613), .A2(n83614), .A3(n83615), .ZN(n83612) );
  NOR2_X1 U69196 ( .A1(n103638), .A2(n105166), .ZN(n83615) );
  AOI21_X1 U69197 ( .B1(n83616), .B2(n83617), .A(n106327), .ZN(n83614) );
  NOR4_X1 U69198 ( .A1(n83618), .A2(n83619), .A3(n83620), .A4(n83621), .ZN(
        n83617) );
  OAI21_X1 U69199 ( .B1(n103642), .B2(n105168), .A(n83622), .ZN(n83621) );
  AOI22_X1 U69200 ( .A1(n105884), .A2(n108186), .B1(n105883), .B2(n108191), 
        .ZN(n83622) );
  NAND2_X1 U69201 ( .A1(n83623), .A2(n83624), .ZN(n83620) );
  AOI22_X1 U69202 ( .A1(n105882), .A2(n108195), .B1(n105881), .B2(n70781), 
        .ZN(n83624) );
  AOI22_X1 U69203 ( .A1(n105880), .A2(n108236), .B1(n83129), .B2(n70769), .ZN(
        n83623) );
  OAI21_X1 U69204 ( .B1(n101006), .B2(n106738), .A(n83625), .ZN(n83619) );
  AOI22_X1 U69205 ( .A1(n105878), .A2(n108223), .B1(n105877), .B2(n108207), 
        .ZN(n83625) );
  NAND2_X1 U69206 ( .A1(n83626), .A2(n83627), .ZN(n83618) );
  AOI22_X1 U69207 ( .A1(n105876), .A2(n108233), .B1(n83136), .B2(n70821), .ZN(
        n83627) );
  AOI22_X1 U69208 ( .A1(n105874), .A2(n108215), .B1(n105873), .B2(n108219), 
        .ZN(n83626) );
  NOR4_X1 U69209 ( .A1(n83628), .A2(n83629), .A3(n83630), .A4(n83631), .ZN(
        n83616) );
  OAI21_X1 U69210 ( .B1(n103651), .B2(n105872), .A(n83632), .ZN(n83631) );
  NAND2_X1 U69212 ( .A1(n83633), .A2(n83634), .ZN(n83630) );
  AOI22_X1 U69213 ( .A1(n105870), .A2(n108247), .B1(n70729), .B2(n105869), 
        .ZN(n83634) );
  AOI22_X1 U69214 ( .A1(n105868), .A2(n108250), .B1(n105867), .B2(n108184), 
        .ZN(n83633) );
  OAI21_X1 U69215 ( .B1(n103650), .B2(n105169), .A(n83635), .ZN(n83629) );
  AOI22_X1 U69216 ( .A1(n70741), .A2(n105866), .B1(n70733), .B2(n105865), .ZN(
        n83635) );
  NAND2_X1 U69217 ( .A1(n83636), .A2(n83637), .ZN(n83628) );
  AOI22_X1 U69218 ( .A1(n105863), .A2(n108201), .B1(n105862), .B2(n108181), 
        .ZN(n83637) );
  AOI22_X1 U69219 ( .A1(n105861), .A2(n108176), .B1(n105860), .B2(n108172), 
        .ZN(n83636) );
  AOI22_X1 U69221 ( .A1(n105857), .A2(n108165), .B1(n105856), .B2(n108178), 
        .ZN(n83611) );
  AOI22_X1 U69222 ( .A1(n105855), .A2(n108227), .B1(n105854), .B2(n108258), 
        .ZN(n83610) );
  AOI22_X1 U69223 ( .A1(n106286), .A2(n108201), .B1(n70769), .B2(n106283), 
        .ZN(n83609) );
  NAND4_X2 U69224 ( .A1(n83638), .A2(n83639), .A3(n83640), .A4(n83641), .ZN(
        n58847) );
  NOR3_X1 U69225 ( .A1(n83642), .A2(n83643), .A3(n83644), .ZN(n83641) );
  NOR2_X1 U69226 ( .A1(n103620), .A2(n106737), .ZN(n83644) );
  AOI21_X1 U69227 ( .B1(n83645), .B2(n83646), .A(n106327), .ZN(n83643) );
  NOR4_X1 U69228 ( .A1(n83647), .A2(n83648), .A3(n83649), .A4(n83650), .ZN(
        n83646) );
  OAI21_X1 U69229 ( .B1(n103624), .B2(n105168), .A(n83651), .ZN(n83650) );
  AOI22_X1 U69230 ( .A1(n105884), .A2(n108309), .B1(n105883), .B2(n108314), 
        .ZN(n83651) );
  NAND2_X1 U69231 ( .A1(n83652), .A2(n83653), .ZN(n83649) );
  AOI22_X1 U69232 ( .A1(n105882), .A2(n108318), .B1(n105881), .B2(n70940), 
        .ZN(n83653) );
  AOI22_X1 U69233 ( .A1(n105880), .A2(n108359), .B1(n70928), .B2(n105879), 
        .ZN(n83652) );
  OAI21_X1 U69234 ( .B1(n101007), .B2(n105167), .A(n83654), .ZN(n83648) );
  AOI22_X1 U69235 ( .A1(n105878), .A2(n108346), .B1(n105877), .B2(n108330), 
        .ZN(n83654) );
  NAND2_X1 U69236 ( .A1(n83655), .A2(n83656), .ZN(n83647) );
  AOI22_X1 U69237 ( .A1(n105876), .A2(n108356), .B1(n70980), .B2(n105875), 
        .ZN(n83656) );
  AOI22_X1 U69238 ( .A1(n105874), .A2(n108338), .B1(n83138), .B2(n108342), 
        .ZN(n83655) );
  NOR4_X1 U69239 ( .A1(n83657), .A2(n83658), .A3(n83659), .A4(n83660), .ZN(
        n83645) );
  OAI21_X1 U69240 ( .B1(n103634), .B2(n105872), .A(n83661), .ZN(n83660) );
  NAND2_X1 U69242 ( .A1(n83662), .A2(n83663), .ZN(n83659) );
  AOI22_X1 U69243 ( .A1(n105870), .A2(n108370), .B1(n70888), .B2(n105869), 
        .ZN(n83663) );
  AOI22_X1 U69244 ( .A1(n105868), .A2(n108373), .B1(n105867), .B2(n108307), 
        .ZN(n83662) );
  OAI21_X1 U69245 ( .B1(n103632), .B2(n106741), .A(n83664), .ZN(n83658) );
  AOI22_X1 U69246 ( .A1(n70900), .A2(n105866), .B1(n70892), .B2(n105865), .ZN(
        n83664) );
  NAND2_X1 U69247 ( .A1(n83665), .A2(n83666), .ZN(n83657) );
  AOI22_X1 U69248 ( .A1(n105863), .A2(n108324), .B1(n105862), .B2(n108304), 
        .ZN(n83666) );
  AOI22_X1 U69249 ( .A1(n105861), .A2(n108299), .B1(n105860), .B2(n108295), 
        .ZN(n83665) );
  AND2_X2 U69250 ( .A1(n105859), .A2(n70999), .ZN(n83642) );
  AOI22_X1 U69251 ( .A1(n105857), .A2(n108288), .B1(n105856), .B2(n108301), 
        .ZN(n83640) );
  AOI22_X1 U69252 ( .A1(n105855), .A2(n108350), .B1(n105854), .B2(n108381), 
        .ZN(n83639) );
  AOI22_X1 U69253 ( .A1(n106286), .A2(n108324), .B1(n70928), .B2(n106284), 
        .ZN(n83638) );
  NAND4_X2 U69254 ( .A1(n83667), .A2(n83668), .A3(n83669), .A4(n83670), .ZN(
        n58846) );
  NOR3_X1 U69255 ( .A1(n83671), .A2(n83672), .A3(n83673), .ZN(n83670) );
  NOR2_X1 U69256 ( .A1(n103601), .A2(n105166), .ZN(n83673) );
  AOI21_X1 U69257 ( .B1(n83674), .B2(n83675), .A(n106327), .ZN(n83672) );
  NOR4_X1 U69258 ( .A1(n83676), .A2(n83677), .A3(n83678), .A4(n83679), .ZN(
        n83675) );
  OAI21_X1 U69259 ( .B1(n103605), .B2(n105168), .A(n83680), .ZN(n83679) );
  AOI22_X1 U69260 ( .A1(n83122), .A2(n108420), .B1(n83123), .B2(n108425), .ZN(
        n83680) );
  NAND2_X1 U69261 ( .A1(n83681), .A2(n83682), .ZN(n83678) );
  AOI22_X1 U69262 ( .A1(n105882), .A2(n108429), .B1(n105881), .B2(n71085), 
        .ZN(n83682) );
  AOI22_X1 U69263 ( .A1(n105880), .A2(n108470), .B1(n105879), .B2(n71073), 
        .ZN(n83681) );
  OAI21_X1 U69264 ( .B1(n101008), .B2(n106738), .A(n83683), .ZN(n83677) );
  AOI22_X1 U69265 ( .A1(n83131), .A2(n108457), .B1(n83132), .B2(n108441), .ZN(
        n83683) );
  NAND2_X1 U69266 ( .A1(n83684), .A2(n83685), .ZN(n83676) );
  AOI22_X1 U69267 ( .A1(n105876), .A2(n108467), .B1(n83136), .B2(n71125), .ZN(
        n83685) );
  AOI22_X1 U69268 ( .A1(n105874), .A2(n108449), .B1(n83138), .B2(n108453), 
        .ZN(n83684) );
  NOR4_X1 U69269 ( .A1(n83686), .A2(n83687), .A3(n83688), .A4(n83689), .ZN(
        n83674) );
  OAI21_X1 U69270 ( .B1(n103616), .B2(n105872), .A(n83690), .ZN(n83689) );
  NAND2_X1 U69272 ( .A1(n83691), .A2(n83692), .ZN(n83688) );
  AOI22_X1 U69273 ( .A1(n105870), .A2(n108481), .B1(n71033), .B2(n105869), 
        .ZN(n83692) );
  AOI22_X1 U69274 ( .A1(n105868), .A2(n108484), .B1(n105867), .B2(n108418), 
        .ZN(n83691) );
  OAI21_X1 U69275 ( .B1(n103614), .B2(n105169), .A(n83693), .ZN(n83687) );
  AOI22_X1 U69276 ( .A1(n71045), .A2(n105866), .B1(n71037), .B2(n83155), .ZN(
        n83693) );
  NAND2_X1 U69277 ( .A1(n83694), .A2(n83695), .ZN(n83686) );
  AOI22_X1 U69278 ( .A1(n105863), .A2(n108435), .B1(n83159), .B2(n108415), 
        .ZN(n83695) );
  AOI22_X1 U69279 ( .A1(n105861), .A2(n108410), .B1(n83161), .B2(n108406), 
        .ZN(n83694) );
  AOI22_X1 U69281 ( .A1(n105857), .A2(n108399), .B1(n105856), .B2(n108412), 
        .ZN(n83669) );
  AOI22_X1 U69282 ( .A1(n105855), .A2(n108461), .B1(n105854), .B2(n108492), 
        .ZN(n83668) );
  AOI22_X1 U69283 ( .A1(n106286), .A2(n108435), .B1(n71073), .B2(n106285), 
        .ZN(n83667) );
  NAND4_X2 U69284 ( .A1(n83696), .A2(n83697), .A3(n83698), .A4(n83699), .ZN(
        n58845) );
  NOR3_X1 U69285 ( .A1(n83700), .A2(n83701), .A3(n83702), .ZN(n83699) );
  NOR2_X1 U69286 ( .A1(n103583), .A2(n106737), .ZN(n83702) );
  AOI21_X1 U69287 ( .B1(n83703), .B2(n83704), .A(n106327), .ZN(n83701) );
  NOR4_X1 U69288 ( .A1(n83705), .A2(n83706), .A3(n83707), .A4(n83708), .ZN(
        n83704) );
  OAI21_X1 U69289 ( .B1(n103587), .B2(n106739), .A(n83709), .ZN(n83708) );
  AOI22_X1 U69290 ( .A1(n83122), .A2(n107658), .B1(n83123), .B2(n107663), .ZN(
        n83709) );
  NAND2_X1 U69291 ( .A1(n83710), .A2(n83711), .ZN(n83707) );
  AOI22_X1 U69292 ( .A1(n105882), .A2(n107667), .B1(n70046), .B2(n83127), .ZN(
        n83711) );
  AOI22_X1 U69293 ( .A1(n105880), .A2(n107708), .B1(n70034), .B2(n105879), 
        .ZN(n83710) );
  OAI21_X1 U69294 ( .B1(n101009), .B2(n105167), .A(n83712), .ZN(n83706) );
  AOI22_X1 U69295 ( .A1(n83131), .A2(n107695), .B1(n83132), .B2(n107679), .ZN(
        n83712) );
  NAND2_X1 U69296 ( .A1(n83713), .A2(n83714), .ZN(n83705) );
  AOI22_X1 U69297 ( .A1(n105876), .A2(n107705), .B1(n70086), .B2(n105875), 
        .ZN(n83714) );
  AOI22_X1 U69298 ( .A1(n83137), .A2(n107687), .B1(n83138), .B2(n107691), .ZN(
        n83713) );
  NOR4_X1 U69299 ( .A1(n83715), .A2(n83716), .A3(n83717), .A4(n83718), .ZN(
        n83703) );
  OAI21_X1 U69300 ( .B1(n103597), .B2(n105872), .A(n83719), .ZN(n83718) );
  NAND2_X1 U69302 ( .A1(n83720), .A2(n83721), .ZN(n83717) );
  AOI22_X1 U69303 ( .A1(n105870), .A2(n107718), .B1(n69994), .B2(n105869), 
        .ZN(n83721) );
  AOI22_X1 U69304 ( .A1(n105868), .A2(n107721), .B1(n105867), .B2(n107656), 
        .ZN(n83720) );
  OAI21_X1 U69305 ( .B1(n103595), .B2(n105169), .A(n83722), .ZN(n83716) );
  AOI22_X1 U69306 ( .A1(n70006), .A2(n105866), .B1(n69998), .B2(n83155), .ZN(
        n83722) );
  NAND2_X1 U69307 ( .A1(n83723), .A2(n83724), .ZN(n83715) );
  AOI22_X1 U69308 ( .A1(n105863), .A2(n107673), .B1(n83159), .B2(n107653), 
        .ZN(n83724) );
  AOI22_X1 U69309 ( .A1(n105861), .A2(n107648), .B1(n83161), .B2(n107644), 
        .ZN(n83723) );
  AND2_X2 U69310 ( .A1(n83162), .A2(n70105), .ZN(n83700) );
  AOI22_X1 U69311 ( .A1(n105857), .A2(n107637), .B1(n83164), .B2(n107650), 
        .ZN(n83698) );
  AOI22_X1 U69312 ( .A1(n105855), .A2(n107699), .B1(n83166), .B2(n107729), 
        .ZN(n83697) );
  AOI22_X1 U69313 ( .A1(n106287), .A2(n107673), .B1(n70034), .B2(n106285), 
        .ZN(n83696) );
  NAND4_X2 U69314 ( .A1(n83725), .A2(n83726), .A3(n83727), .A4(n83728), .ZN(
        n58844) );
  NOR3_X1 U69315 ( .A1(n83729), .A2(n83730), .A3(n83731), .ZN(n83728) );
  NOR2_X1 U69316 ( .A1(n103566), .A2(n105166), .ZN(n83731) );
  AOI21_X1 U69317 ( .B1(n83732), .B2(n83733), .A(n106327), .ZN(n83730) );
  NOR4_X1 U69318 ( .A1(n83734), .A2(n83735), .A3(n83736), .A4(n83737), .ZN(
        n83733) );
  OAI21_X1 U69319 ( .B1(n103569), .B2(n106739), .A(n83738), .ZN(n83737) );
  AOI22_X1 U69320 ( .A1(n83122), .A2(n109576), .B1(n83123), .B2(n109581), .ZN(
        n83738) );
  NAND2_X1 U69321 ( .A1(n83739), .A2(n83740), .ZN(n83736) );
  AOI22_X1 U69322 ( .A1(n105882), .A2(n109585), .B1(n72575), .B2(n83127), .ZN(
        n83740) );
  AOI22_X1 U69323 ( .A1(n105880), .A2(n109623), .B1(n72563), .B2(n105879), 
        .ZN(n83739) );
  OAI21_X1 U69324 ( .B1(n101010), .B2(n106738), .A(n83741), .ZN(n83735) );
  AOI22_X1 U69325 ( .A1(n72607), .A2(n105878), .B1(n83132), .B2(n109597), .ZN(
        n83741) );
  NAND2_X1 U69326 ( .A1(n83742), .A2(n83743), .ZN(n83734) );
  AOI22_X1 U69327 ( .A1(n105876), .A2(n109620), .B1(n72615), .B2(n105875), 
        .ZN(n83743) );
  AOI22_X1 U69328 ( .A1(n83137), .A2(n109605), .B1(n72603), .B2(n105873), .ZN(
        n83742) );
  NOR4_X1 U69329 ( .A1(n83744), .A2(n83745), .A3(n83746), .A4(n83747), .ZN(
        n83732) );
  OAI21_X1 U69330 ( .B1(n103579), .B2(n83143), .A(n83748), .ZN(n83747) );
  NAND2_X1 U69332 ( .A1(n83749), .A2(n83750), .ZN(n83746) );
  AOI22_X1 U69333 ( .A1(n105870), .A2(n109633), .B1(n72523), .B2(n105869), 
        .ZN(n83750) );
  AOI22_X1 U69334 ( .A1(n105868), .A2(n109636), .B1(n105867), .B2(n109574), 
        .ZN(n83749) );
  OAI21_X1 U69335 ( .B1(n103578), .B2(n105169), .A(n83751), .ZN(n83745) );
  AOI22_X1 U69336 ( .A1(n72535), .A2(n105866), .B1(n72527), .B2(n83155), .ZN(
        n83751) );
  NAND2_X1 U69337 ( .A1(n83752), .A2(n83753), .ZN(n83744) );
  AOI22_X1 U69338 ( .A1(n105863), .A2(n109591), .B1(n83159), .B2(n109571), 
        .ZN(n83753) );
  AOI22_X1 U69339 ( .A1(n105861), .A2(n109566), .B1(n83161), .B2(n109562), 
        .ZN(n83752) );
  AND2_X2 U69340 ( .A1(n105859), .A2(n72634), .ZN(n83729) );
  AOI22_X1 U69341 ( .A1(n105857), .A2(n109555), .B1(n83164), .B2(n109568), 
        .ZN(n83727) );
  AOI22_X1 U69342 ( .A1(n105855), .A2(n109614), .B1(n83166), .B2(n109644), 
        .ZN(n83726) );
  AOI22_X1 U69343 ( .A1(n106287), .A2(n109591), .B1(n72563), .B2(n106285), 
        .ZN(n83725) );
  NAND4_X2 U69344 ( .A1(n83754), .A2(n83755), .A3(n83756), .A4(n83757), .ZN(
        n58843) );
  NOR3_X1 U69345 ( .A1(n83758), .A2(n83759), .A3(n83760), .ZN(n83757) );
  NOR2_X1 U69346 ( .A1(n103548), .A2(n105166), .ZN(n83760) );
  AOI21_X1 U69347 ( .B1(n83761), .B2(n83762), .A(n106323), .ZN(n83759) );
  NOR4_X1 U69348 ( .A1(n83763), .A2(n83764), .A3(n83765), .A4(n83766), .ZN(
        n83762) );
  OAI21_X1 U69349 ( .B1(n103552), .B2(n105864), .A(n83767), .ZN(n83766) );
  AOI22_X1 U69350 ( .A1(n105883), .A2(n108542), .B1(n83239), .B2(n108555), 
        .ZN(n83767) );
  NAND2_X1 U69351 ( .A1(n83768), .A2(n83769), .ZN(n83765) );
  AOI22_X1 U69352 ( .A1(n105881), .A2(n71234), .B1(n83128), .B2(n108585), .ZN(
        n83769) );
  AOI22_X1 U69353 ( .A1(n105879), .A2(n71222), .B1(n105884), .B2(n108537), 
        .ZN(n83768) );
  NAND2_X1 U69354 ( .A1(n83770), .A2(n83771), .ZN(n83764) );
  AOI22_X1 U69355 ( .A1(n71266), .A2(n105878), .B1(n83132), .B2(n108558), .ZN(
        n83771) );
  AOI22_X1 U69356 ( .A1(n83244), .A2(n108561), .B1(n83126), .B2(n108546), .ZN(
        n83770) );
  NAND2_X1 U69357 ( .A1(n83772), .A2(n83773), .ZN(n83763) );
  AOI22_X1 U69358 ( .A1(n105876), .A2(n108582), .B1(n83136), .B2(n71274), .ZN(
        n83773) );
  AOI22_X1 U69359 ( .A1(n83137), .A2(n108566), .B1(n83138), .B2(n71262), .ZN(
        n83772) );
  NOR4_X1 U69360 ( .A1(n83774), .A2(n83775), .A3(n83776), .A4(n83777), .ZN(
        n83761) );
  OAI21_X1 U69361 ( .B1(n103562), .B2(n83143), .A(n83778), .ZN(n83777) );
  NAND2_X1 U69363 ( .A1(n83779), .A2(n83780), .ZN(n83776) );
  AOI22_X1 U69364 ( .A1(n105870), .A2(n108595), .B1(n71182), .B2(n105869), 
        .ZN(n83780) );
  AOI22_X1 U69365 ( .A1(n105868), .A2(n108598), .B1(n105867), .B2(n108535), 
        .ZN(n83779) );
  OAI21_X1 U69366 ( .B1(n83254), .B2(n104615), .A(n83781), .ZN(n83775) );
  AOI22_X1 U69367 ( .A1(n105865), .A2(n71186), .B1(n83256), .B2(n108590), .ZN(
        n83781) );
  NAND2_X1 U69368 ( .A1(n83782), .A2(n83783), .ZN(n83774) );
  AOI22_X1 U69369 ( .A1(n105862), .A2(n108532), .B1(n105861), .B2(n108527), 
        .ZN(n83783) );
  AOI22_X1 U69370 ( .A1(n105860), .A2(n108523), .B1(n71194), .B2(n83154), .ZN(
        n83782) );
  NOR2_X1 U69371 ( .A1(n103559), .A2(n105858), .ZN(n83758) );
  AOI22_X1 U69372 ( .A1(n105856), .A2(n108529), .B1(n83165), .B2(n108576), 
        .ZN(n83756) );
  AOI22_X1 U69373 ( .A1(n105854), .A2(n108606), .B1(n106289), .B2(n108552), 
        .ZN(n83755) );
  AOI22_X1 U69374 ( .A1(n71222), .A2(n80260), .B1(n71293), .B2(n83259), .ZN(
        n83754) );
  NAND4_X2 U69375 ( .A1(n83784), .A2(n83785), .A3(n83786), .A4(n83787), .ZN(
        n58842) );
  NOR3_X1 U69376 ( .A1(n83788), .A2(n83789), .A3(n83790), .ZN(n83787) );
  NOR2_X1 U69377 ( .A1(n103530), .A2(n105166), .ZN(n83790) );
  AOI21_X1 U69378 ( .B1(n83791), .B2(n83792), .A(n106323), .ZN(n83789) );
  NOR4_X1 U69379 ( .A1(n83793), .A2(n83794), .A3(n83795), .A4(n83796), .ZN(
        n83792) );
  OAI21_X1 U69380 ( .B1(n103533), .B2(n106739), .A(n83797), .ZN(n83796) );
  AOI22_X1 U69381 ( .A1(n83122), .A2(n109681), .B1(n83123), .B2(n109686), .ZN(
        n83797) );
  NAND2_X1 U69382 ( .A1(n83798), .A2(n83799), .ZN(n83795) );
  AOI22_X1 U69383 ( .A1(n105882), .A2(n109690), .B1(n72717), .B2(n83127), .ZN(
        n83799) );
  AOI22_X1 U69384 ( .A1(n105880), .A2(n109730), .B1(n72705), .B2(n105879), 
        .ZN(n83798) );
  OAI21_X1 U69385 ( .B1(n101012), .B2(n106738), .A(n83800), .ZN(n83794) );
  AOI22_X1 U69386 ( .A1(n83131), .A2(n109717), .B1(n83132), .B2(n109702), .ZN(
        n83800) );
  NAND2_X1 U69387 ( .A1(n83801), .A2(n83802), .ZN(n83793) );
  AOI22_X1 U69388 ( .A1(n105876), .A2(n109727), .B1(n72757), .B2(n105875), 
        .ZN(n83802) );
  AOI22_X1 U69389 ( .A1(n83137), .A2(n109710), .B1(n72745), .B2(n105873), .ZN(
        n83801) );
  NOR4_X1 U69390 ( .A1(n83803), .A2(n83804), .A3(n83805), .A4(n83806), .ZN(
        n83791) );
  OAI21_X1 U69391 ( .B1(n103544), .B2(n83143), .A(n83807), .ZN(n83806) );
  NAND2_X1 U69393 ( .A1(n83808), .A2(n83809), .ZN(n83805) );
  AOI22_X1 U69394 ( .A1(n105870), .A2(n109740), .B1(n72665), .B2(n105869), 
        .ZN(n83809) );
  AOI22_X1 U69395 ( .A1(n105868), .A2(n109743), .B1(n105867), .B2(n109679), 
        .ZN(n83808) );
  OAI21_X1 U69396 ( .B1(n103542), .B2(n105169), .A(n83810), .ZN(n83804) );
  AOI22_X1 U69397 ( .A1(n72677), .A2(n105866), .B1(n72669), .B2(n83155), .ZN(
        n83810) );
  NAND2_X1 U69398 ( .A1(n83811), .A2(n83812), .ZN(n83803) );
  AOI22_X1 U69399 ( .A1(n105863), .A2(n109696), .B1(n83159), .B2(n109676), 
        .ZN(n83812) );
  AOI22_X1 U69400 ( .A1(n105861), .A2(n109671), .B1(n83161), .B2(n109667), 
        .ZN(n83811) );
  AND2_X2 U69401 ( .A1(n83162), .A2(n72776), .ZN(n83788) );
  AOI22_X1 U69402 ( .A1(n105857), .A2(n109660), .B1(n83164), .B2(n109673), 
        .ZN(n83786) );
  AOI22_X1 U69403 ( .A1(n105855), .A2(n109721), .B1(n83166), .B2(n109751), 
        .ZN(n83785) );
  AOI22_X1 U69404 ( .A1(n106288), .A2(n109696), .B1(n72705), .B2(n106285), 
        .ZN(n83784) );
  NAND4_X2 U69405 ( .A1(n83813), .A2(n83814), .A3(n83815), .A4(n83816), .ZN(
        n58841) );
  NOR3_X1 U69406 ( .A1(n83817), .A2(n83818), .A3(n83819), .ZN(n83816) );
  NOR2_X1 U69407 ( .A1(n103511), .A2(n105166), .ZN(n83819) );
  AOI21_X1 U69408 ( .B1(n83820), .B2(n83821), .A(n106323), .ZN(n83818) );
  NOR4_X1 U69409 ( .A1(n83822), .A2(n83823), .A3(n83824), .A4(n83825), .ZN(
        n83821) );
  OAI21_X1 U69410 ( .B1(n103515), .B2(n106739), .A(n83826), .ZN(n83825) );
  AOI22_X1 U69411 ( .A1(n83122), .A2(n109465), .B1(n83123), .B2(n109470), .ZN(
        n83826) );
  NAND2_X1 U69412 ( .A1(n83827), .A2(n83828), .ZN(n83824) );
  AOI22_X1 U69413 ( .A1(n83126), .A2(n109474), .B1(n72427), .B2(n83127), .ZN(
        n83828) );
  AOI22_X1 U69414 ( .A1(n83128), .A2(n109515), .B1(n72415), .B2(n83129), .ZN(
        n83827) );
  OAI21_X1 U69415 ( .B1(n101013), .B2(n106738), .A(n83829), .ZN(n83823) );
  AOI22_X1 U69416 ( .A1(n83131), .A2(n109502), .B1(n83132), .B2(n109486), .ZN(
        n83829) );
  NAND2_X1 U69417 ( .A1(n83830), .A2(n83831), .ZN(n83822) );
  AOI22_X1 U69418 ( .A1(n105876), .A2(n109512), .B1(n72467), .B2(n83136), .ZN(
        n83831) );
  AOI22_X1 U69419 ( .A1(n83137), .A2(n109494), .B1(n83138), .B2(n109498), .ZN(
        n83830) );
  NOR4_X1 U69420 ( .A1(n83832), .A2(n83833), .A3(n83834), .A4(n83835), .ZN(
        n83820) );
  OAI21_X1 U69421 ( .B1(n103526), .B2(n83143), .A(n83836), .ZN(n83835) );
  NAND2_X1 U69423 ( .A1(n83837), .A2(n83838), .ZN(n83834) );
  AOI22_X1 U69424 ( .A1(n105870), .A2(n109525), .B1(n72375), .B2(n105869), 
        .ZN(n83838) );
  AOI22_X1 U69425 ( .A1(n105868), .A2(n109528), .B1(n105867), .B2(n109463), 
        .ZN(n83837) );
  OAI21_X1 U69426 ( .B1(n103524), .B2(n105169), .A(n83839), .ZN(n83833) );
  AOI22_X1 U69427 ( .A1(n72387), .A2(n83154), .B1(n72379), .B2(n83155), .ZN(
        n83839) );
  NAND2_X1 U69428 ( .A1(n83840), .A2(n83841), .ZN(n83832) );
  AOI22_X1 U69429 ( .A1(n105863), .A2(n109480), .B1(n83159), .B2(n109460), 
        .ZN(n83841) );
  AOI22_X1 U69430 ( .A1(n105861), .A2(n109455), .B1(n83161), .B2(n109451), 
        .ZN(n83840) );
  AND2_X2 U69431 ( .A1(n105859), .A2(n72486), .ZN(n83817) );
  AOI22_X1 U69432 ( .A1(n105857), .A2(n109444), .B1(n83164), .B2(n109457), 
        .ZN(n83815) );
  AOI22_X1 U69433 ( .A1(n83165), .A2(n109506), .B1(n83166), .B2(n109536), .ZN(
        n83814) );
  AOI22_X1 U69434 ( .A1(n106289), .A2(n109480), .B1(n72415), .B2(n106285), 
        .ZN(n83813) );
  NAND4_X2 U69435 ( .A1(n83842), .A2(n83843), .A3(n83844), .A4(n83845), .ZN(
        n58840) );
  NOR3_X1 U69436 ( .A1(n83846), .A2(n83847), .A3(n83848), .ZN(n83845) );
  NOR2_X1 U69437 ( .A1(n103492), .A2(n105166), .ZN(n83848) );
  AOI21_X1 U69438 ( .B1(n83849), .B2(n83850), .A(n106323), .ZN(n83847) );
  NOR4_X1 U69439 ( .A1(n83851), .A2(n83852), .A3(n83853), .A4(n83854), .ZN(
        n83850) );
  OAI21_X1 U69440 ( .B1(n103496), .B2(n106739), .A(n83855), .ZN(n83854) );
  AOI22_X1 U69441 ( .A1(n83122), .A2(n109002), .B1(n83123), .B2(n109007), .ZN(
        n83855) );
  NAND2_X1 U69442 ( .A1(n83856), .A2(n83857), .ZN(n83853) );
  AOI22_X1 U69443 ( .A1(n83126), .A2(n109011), .B1(n71827), .B2(n83127), .ZN(
        n83857) );
  AOI22_X1 U69444 ( .A1(n83128), .A2(n109052), .B1(n71815), .B2(n105879), .ZN(
        n83856) );
  OAI21_X1 U69445 ( .B1(n101014), .B2(n106738), .A(n83858), .ZN(n83852) );
  AOI22_X1 U69446 ( .A1(n83131), .A2(n109039), .B1(n83132), .B2(n109023), .ZN(
        n83858) );
  NAND2_X1 U69447 ( .A1(n83859), .A2(n83860), .ZN(n83851) );
  AOI22_X1 U69448 ( .A1(n105876), .A2(n109049), .B1(n71867), .B2(n83136), .ZN(
        n83860) );
  AOI22_X1 U69449 ( .A1(n83137), .A2(n109031), .B1(n83138), .B2(n109035), .ZN(
        n83859) );
  NOR4_X1 U69450 ( .A1(n83861), .A2(n83862), .A3(n83863), .A4(n83864), .ZN(
        n83849) );
  OAI21_X1 U69451 ( .B1(n103507), .B2(n83143), .A(n83865), .ZN(n83864) );
  NAND2_X1 U69453 ( .A1(n83866), .A2(n83867), .ZN(n83863) );
  AOI22_X1 U69454 ( .A1(n105870), .A2(n109063), .B1(n71775), .B2(n105869), 
        .ZN(n83867) );
  AOI22_X1 U69455 ( .A1(n105868), .A2(n109066), .B1(n105867), .B2(n109000), 
        .ZN(n83866) );
  OAI21_X1 U69456 ( .B1(n103505), .B2(n105169), .A(n83868), .ZN(n83862) );
  AOI22_X1 U69457 ( .A1(n71787), .A2(n83154), .B1(n71779), .B2(n83155), .ZN(
        n83868) );
  NAND2_X1 U69458 ( .A1(n83869), .A2(n83870), .ZN(n83861) );
  AOI22_X1 U69459 ( .A1(n105863), .A2(n109017), .B1(n83159), .B2(n108997), 
        .ZN(n83870) );
  AOI22_X1 U69460 ( .A1(n105861), .A2(n108992), .B1(n83161), .B2(n108988), 
        .ZN(n83869) );
  AND2_X2 U69461 ( .A1(n83162), .A2(n71886), .ZN(n83846) );
  AOI22_X1 U69462 ( .A1(n105857), .A2(n108981), .B1(n83164), .B2(n108994), 
        .ZN(n83844) );
  AOI22_X1 U69463 ( .A1(n83165), .A2(n109043), .B1(n83166), .B2(n109074), .ZN(
        n83843) );
  AOI22_X1 U69464 ( .A1(n106286), .A2(n109017), .B1(n71815), .B2(n106285), 
        .ZN(n83842) );
  NAND4_X2 U69465 ( .A1(n83871), .A2(n83872), .A3(n83873), .A4(n83874), .ZN(
        n58839) );
  NOR3_X1 U69466 ( .A1(n83875), .A2(n83876), .A3(n83877), .ZN(n83874) );
  NOR2_X1 U69467 ( .A1(n103473), .A2(n105166), .ZN(n83877) );
  AOI21_X1 U69468 ( .B1(n83878), .B2(n83879), .A(n106323), .ZN(n83876) );
  NOR4_X1 U69469 ( .A1(n83880), .A2(n83881), .A3(n83882), .A4(n83883), .ZN(
        n83879) );
  OAI21_X1 U69470 ( .B1(n103477), .B2(n106739), .A(n83884), .ZN(n83883) );
  AOI22_X1 U69471 ( .A1(n83122), .A2(n109350), .B1(n83123), .B2(n109355), .ZN(
        n83884) );
  NAND2_X1 U69472 ( .A1(n83885), .A2(n83886), .ZN(n83882) );
  AOI22_X1 U69473 ( .A1(n83126), .A2(n109359), .B1(n105881), .B2(n72276), .ZN(
        n83886) );
  AOI22_X1 U69474 ( .A1(n83128), .A2(n109400), .B1(n83129), .B2(n72264), .ZN(
        n83885) );
  OAI21_X1 U69475 ( .B1(n101015), .B2(n105167), .A(n83887), .ZN(n83881) );
  AOI22_X1 U69476 ( .A1(n83131), .A2(n109387), .B1(n83132), .B2(n109371), .ZN(
        n83887) );
  NAND2_X1 U69477 ( .A1(n83888), .A2(n83889), .ZN(n83880) );
  AOI22_X1 U69478 ( .A1(n105876), .A2(n109397), .B1(n83136), .B2(n72316), .ZN(
        n83889) );
  AOI22_X1 U69479 ( .A1(n83137), .A2(n109379), .B1(n83138), .B2(n109383), .ZN(
        n83888) );
  NOR4_X1 U69480 ( .A1(n83890), .A2(n83891), .A3(n83892), .A4(n83893), .ZN(
        n83878) );
  OAI21_X1 U69481 ( .B1(n103488), .B2(n83143), .A(n83894), .ZN(n83893) );
  NAND2_X1 U69483 ( .A1(n83895), .A2(n83896), .ZN(n83892) );
  AOI22_X1 U69484 ( .A1(n105870), .A2(n109410), .B1(n72224), .B2(n105869), 
        .ZN(n83896) );
  AOI22_X1 U69485 ( .A1(n105868), .A2(n109413), .B1(n105867), .B2(n109348), 
        .ZN(n83895) );
  OAI21_X1 U69486 ( .B1(n103486), .B2(n105169), .A(n83897), .ZN(n83891) );
  AOI22_X1 U69487 ( .A1(n72236), .A2(n83154), .B1(n105865), .B2(n72228), .ZN(
        n83897) );
  NAND2_X1 U69488 ( .A1(n83898), .A2(n83899), .ZN(n83890) );
  AOI22_X1 U69489 ( .A1(n105863), .A2(n109365), .B1(n83159), .B2(n109345), 
        .ZN(n83899) );
  AOI22_X1 U69490 ( .A1(n105861), .A2(n109340), .B1(n83161), .B2(n109336), 
        .ZN(n83898) );
  AND2_X2 U69491 ( .A1(n105859), .A2(n72335), .ZN(n83875) );
  AOI22_X1 U69492 ( .A1(n105857), .A2(n109329), .B1(n83164), .B2(n109342), 
        .ZN(n83873) );
  AOI22_X1 U69493 ( .A1(n83165), .A2(n109391), .B1(n83166), .B2(n109421), .ZN(
        n83872) );
  AOI22_X1 U69494 ( .A1(n106288), .A2(n109365), .B1(n72264), .B2(n106285), 
        .ZN(n83871) );
  NAND4_X2 U69495 ( .A1(n83900), .A2(n83901), .A3(n83902), .A4(n83903), .ZN(
        n58838) );
  NOR3_X1 U69496 ( .A1(n83904), .A2(n83905), .A3(n83906), .ZN(n83903) );
  NOR2_X1 U69497 ( .A1(n103454), .A2(n105166), .ZN(n83906) );
  AOI21_X1 U69498 ( .B1(n83907), .B2(n83908), .A(n106323), .ZN(n83905) );
  NOR4_X1 U69499 ( .A1(n83909), .A2(n83910), .A3(n83911), .A4(n83912), .ZN(
        n83908) );
  OAI21_X1 U69500 ( .B1(n103458), .B2(n106739), .A(n83913), .ZN(n83912) );
  AOI22_X1 U69501 ( .A1(n105884), .A2(n109232), .B1(n83123), .B2(n109237), 
        .ZN(n83913) );
  NAND2_X1 U69502 ( .A1(n83914), .A2(n83915), .ZN(n83911) );
  AOI22_X1 U69503 ( .A1(n83126), .A2(n109241), .B1(n72125), .B2(n83127), .ZN(
        n83915) );
  AOI22_X1 U69504 ( .A1(n83128), .A2(n109281), .B1(n72113), .B2(n105879), .ZN(
        n83914) );
  OAI21_X1 U69505 ( .B1(n101016), .B2(n105167), .A(n83916), .ZN(n83910) );
  AOI22_X1 U69506 ( .A1(n83131), .A2(n109269), .B1(n83132), .B2(n109253), .ZN(
        n83916) );
  NAND2_X1 U69507 ( .A1(n83917), .A2(n83918), .ZN(n83909) );
  AOI22_X1 U69508 ( .A1(n105876), .A2(n109279), .B1(n72165), .B2(n83136), .ZN(
        n83918) );
  AOI22_X1 U69509 ( .A1(n83137), .A2(n109261), .B1(n83138), .B2(n109265), .ZN(
        n83917) );
  NOR4_X1 U69510 ( .A1(n83919), .A2(n83920), .A3(n83921), .A4(n83922), .ZN(
        n83907) );
  OAI21_X1 U69511 ( .B1(n103469), .B2(n83143), .A(n83923), .ZN(n83922) );
  NAND2_X1 U69513 ( .A1(n83924), .A2(n83925), .ZN(n83921) );
  AOI22_X1 U69514 ( .A1(n105870), .A2(n109291), .B1(n72073), .B2(n105869), 
        .ZN(n83925) );
  AOI22_X1 U69515 ( .A1(n105868), .A2(n109294), .B1(n105867), .B2(n109230), 
        .ZN(n83924) );
  OAI21_X1 U69516 ( .B1(n103467), .B2(n105169), .A(n83926), .ZN(n83920) );
  AOI22_X1 U69517 ( .A1(n72085), .A2(n83154), .B1(n72077), .B2(n105865), .ZN(
        n83926) );
  NAND2_X1 U69518 ( .A1(n83927), .A2(n83928), .ZN(n83919) );
  AOI22_X1 U69519 ( .A1(n105863), .A2(n109247), .B1(n83159), .B2(n109227), 
        .ZN(n83928) );
  AOI22_X1 U69520 ( .A1(n105861), .A2(n109222), .B1(n83161), .B2(n109218), 
        .ZN(n83927) );
  AND2_X2 U69521 ( .A1(n105859), .A2(n72184), .ZN(n83904) );
  AOI22_X1 U69522 ( .A1(n105857), .A2(n109211), .B1(n83164), .B2(n109224), 
        .ZN(n83902) );
  AOI22_X1 U69523 ( .A1(n83165), .A2(n109273), .B1(n83166), .B2(n109302), .ZN(
        n83901) );
  AOI22_X1 U69524 ( .A1(n106287), .A2(n109247), .B1(n72113), .B2(n106285), 
        .ZN(n83900) );
  NAND4_X2 U69525 ( .A1(n83929), .A2(n83930), .A3(n83931), .A4(n83932), .ZN(
        n58837) );
  NOR3_X1 U69526 ( .A1(n83933), .A2(n83934), .A3(n83935), .ZN(n83932) );
  NOR2_X1 U69527 ( .A1(n103434), .A2(n105166), .ZN(n83935) );
  AOI21_X1 U69528 ( .B1(n83936), .B2(n83937), .A(n106323), .ZN(n83934) );
  NOR4_X1 U69529 ( .A1(n83938), .A2(n83939), .A3(n83940), .A4(n83941), .ZN(
        n83937) );
  OAI21_X1 U69530 ( .B1(n103438), .B2(n106739), .A(n83942), .ZN(n83941) );
  AOI22_X1 U69531 ( .A1(n105884), .A2(n109124), .B1(n83123), .B2(n109129), 
        .ZN(n83942) );
  NAND2_X1 U69532 ( .A1(n83943), .A2(n83944), .ZN(n83940) );
  AOI22_X1 U69533 ( .A1(n83126), .A2(n109133), .B1(n71981), .B2(n105881), .ZN(
        n83944) );
  AOI22_X1 U69534 ( .A1(n83128), .A2(n109173), .B1(n71969), .B2(n83129), .ZN(
        n83943) );
  OAI21_X1 U69535 ( .B1(n106738), .B2(n104649), .A(n83945), .ZN(n83939) );
  AOI22_X1 U69536 ( .A1(n83131), .A2(n109160), .B1(n83132), .B2(n109145), .ZN(
        n83945) );
  NAND2_X1 U69537 ( .A1(n83946), .A2(n83947), .ZN(n83938) );
  AOI22_X1 U69538 ( .A1(n105876), .A2(n109170), .B1(n72021), .B2(n83136), .ZN(
        n83947) );
  AOI22_X1 U69539 ( .A1(n83137), .A2(n109152), .B1(n83138), .B2(n109156), .ZN(
        n83946) );
  NOR4_X1 U69540 ( .A1(n83948), .A2(n83949), .A3(n83950), .A4(n83951), .ZN(
        n83936) );
  OAI21_X1 U69541 ( .B1(n103449), .B2(n83143), .A(n83952), .ZN(n83951) );
  NAND2_X1 U69543 ( .A1(n83953), .A2(n83954), .ZN(n83950) );
  AOI22_X1 U69544 ( .A1(n105870), .A2(n109183), .B1(n71929), .B2(n105869), 
        .ZN(n83954) );
  AOI22_X1 U69545 ( .A1(n105868), .A2(n109186), .B1(n105867), .B2(n109122), 
        .ZN(n83953) );
  OAI21_X1 U69546 ( .B1(n103447), .B2(n105169), .A(n83955), .ZN(n83949) );
  AOI22_X1 U69547 ( .A1(n71941), .A2(n83154), .B1(n71933), .B2(n105865), .ZN(
        n83955) );
  NAND2_X1 U69548 ( .A1(n83956), .A2(n83957), .ZN(n83948) );
  AOI22_X1 U69549 ( .A1(n105863), .A2(n109139), .B1(n83159), .B2(n109119), 
        .ZN(n83957) );
  AOI22_X1 U69550 ( .A1(n105861), .A2(n109114), .B1(n83161), .B2(n109110), 
        .ZN(n83956) );
  AND2_X2 U69551 ( .A1(n105859), .A2(n72040), .ZN(n83933) );
  AOI22_X1 U69552 ( .A1(n105857), .A2(n109103), .B1(n83164), .B2(n109116), 
        .ZN(n83931) );
  AOI22_X1 U69553 ( .A1(n83165), .A2(n109164), .B1(n83166), .B2(n109194), .ZN(
        n83930) );
  AOI22_X1 U69554 ( .A1(n106288), .A2(n109139), .B1(n71969), .B2(n106285), 
        .ZN(n83929) );
  NAND4_X2 U69555 ( .A1(n83958), .A2(n83959), .A3(n83960), .A4(n83961), .ZN(
        n58836) );
  NOR3_X1 U69556 ( .A1(n83962), .A2(n83963), .A3(n83964), .ZN(n83961) );
  NOR2_X1 U69557 ( .A1(n103414), .A2(n105166), .ZN(n83964) );
  AOI21_X1 U69558 ( .B1(n83965), .B2(n83966), .A(n106323), .ZN(n83963) );
  NOR4_X1 U69559 ( .A1(n83967), .A2(n83968), .A3(n83969), .A4(n83970), .ZN(
        n83966) );
  OAI21_X1 U69560 ( .B1(n103418), .B2(n106739), .A(n83971), .ZN(n83970) );
  AOI22_X1 U69561 ( .A1(n105884), .A2(n108659), .B1(n83123), .B2(n108664), 
        .ZN(n83971) );
  NAND2_X1 U69562 ( .A1(n83972), .A2(n83973), .ZN(n83969) );
  AOI22_X1 U69563 ( .A1(n83126), .A2(n108668), .B1(n71383), .B2(n83127), .ZN(
        n83973) );
  AOI22_X1 U69564 ( .A1(n83128), .A2(n108708), .B1(n71371), .B2(n83129), .ZN(
        n83972) );
  OAI21_X1 U69565 ( .B1(n101017), .B2(n105167), .A(n83974), .ZN(n83968) );
  AOI22_X1 U69566 ( .A1(n83131), .A2(n108696), .B1(n83132), .B2(n108680), .ZN(
        n83974) );
  NAND2_X1 U69567 ( .A1(n83975), .A2(n83976), .ZN(n83967) );
  AOI22_X1 U69568 ( .A1(n105876), .A2(n108706), .B1(n71423), .B2(n83136), .ZN(
        n83976) );
  AOI22_X1 U69569 ( .A1(n83137), .A2(n108688), .B1(n83138), .B2(n108692), .ZN(
        n83975) );
  NOR4_X1 U69570 ( .A1(n83977), .A2(n83978), .A3(n83979), .A4(n83980), .ZN(
        n83965) );
  OAI21_X1 U69571 ( .B1(n103429), .B2(n83143), .A(n83981), .ZN(n83980) );
  NAND2_X1 U69573 ( .A1(n83982), .A2(n83983), .ZN(n83979) );
  AOI22_X1 U69574 ( .A1(n105870), .A2(n108718), .B1(n71331), .B2(n105869), 
        .ZN(n83983) );
  AOI22_X1 U69575 ( .A1(n105868), .A2(n108721), .B1(n105867), .B2(n108657), 
        .ZN(n83982) );
  OAI21_X1 U69576 ( .B1(n103427), .B2(n105169), .A(n83984), .ZN(n83978) );
  AOI22_X1 U69577 ( .A1(n71343), .A2(n83154), .B1(n71335), .B2(n105865), .ZN(
        n83984) );
  NAND2_X1 U69578 ( .A1(n83985), .A2(n83986), .ZN(n83977) );
  AOI22_X1 U69579 ( .A1(n105863), .A2(n108674), .B1(n83159), .B2(n108654), 
        .ZN(n83986) );
  AOI22_X1 U69580 ( .A1(n105861), .A2(n108649), .B1(n83161), .B2(n108645), 
        .ZN(n83985) );
  AND2_X2 U69581 ( .A1(n105859), .A2(n71442), .ZN(n83962) );
  AOI22_X1 U69582 ( .A1(n105857), .A2(n108638), .B1(n83164), .B2(n108651), 
        .ZN(n83960) );
  AOI22_X1 U69583 ( .A1(n83165), .A2(n108700), .B1(n83166), .B2(n108729), .ZN(
        n83959) );
  AOI22_X1 U69584 ( .A1(n106289), .A2(n108674), .B1(n71371), .B2(n106285), 
        .ZN(n83958) );
  NAND4_X2 U69585 ( .A1(n83987), .A2(n83988), .A3(n83989), .A4(n83990), .ZN(
        n58835) );
  NOR3_X1 U69586 ( .A1(n83991), .A2(n83992), .A3(n83993), .ZN(n83990) );
  NOR2_X1 U69587 ( .A1(n103394), .A2(n105166), .ZN(n83993) );
  AOI21_X1 U69588 ( .B1(n83994), .B2(n83995), .A(n106323), .ZN(n83992) );
  NOR4_X1 U69589 ( .A1(n83996), .A2(n83997), .A3(n83998), .A4(n83999), .ZN(
        n83995) );
  OAI21_X1 U69590 ( .B1(n103398), .B2(n106739), .A(n84000), .ZN(n83999) );
  AOI22_X1 U69591 ( .A1(n105884), .A2(n108886), .B1(n83123), .B2(n108891), 
        .ZN(n84000) );
  NAND2_X1 U69592 ( .A1(n84001), .A2(n84002), .ZN(n83998) );
  AOI22_X1 U69593 ( .A1(n83126), .A2(n108895), .B1(n71678), .B2(n105881), .ZN(
        n84002) );
  AOI22_X1 U69594 ( .A1(n83128), .A2(n108936), .B1(n71666), .B2(n83129), .ZN(
        n84001) );
  OAI21_X1 U69595 ( .B1(n101018), .B2(n105167), .A(n84003), .ZN(n83997) );
  AOI22_X1 U69596 ( .A1(n83131), .A2(n108923), .B1(n83132), .B2(n108907), .ZN(
        n84003) );
  NAND2_X1 U69597 ( .A1(n84004), .A2(n84005), .ZN(n83996) );
  AOI22_X1 U69598 ( .A1(n105876), .A2(n108933), .B1(n71718), .B2(n83136), .ZN(
        n84005) );
  AOI22_X1 U69599 ( .A1(n83137), .A2(n108915), .B1(n83138), .B2(n108919), .ZN(
        n84004) );
  NOR4_X1 U69600 ( .A1(n84006), .A2(n84007), .A3(n84008), .A4(n84009), .ZN(
        n83994) );
  OAI21_X1 U69601 ( .B1(n103409), .B2(n83143), .A(n84010), .ZN(n84009) );
  NAND2_X1 U69603 ( .A1(n84011), .A2(n84012), .ZN(n84008) );
  AOI22_X1 U69604 ( .A1(n105870), .A2(n108946), .B1(n71626), .B2(n105869), 
        .ZN(n84012) );
  AOI22_X1 U69605 ( .A1(n105868), .A2(n108949), .B1(n105867), .B2(n108884), 
        .ZN(n84011) );
  OAI21_X1 U69606 ( .B1(n103407), .B2(n105169), .A(n84013), .ZN(n84007) );
  AOI22_X1 U69607 ( .A1(n71638), .A2(n83154), .B1(n71630), .B2(n105865), .ZN(
        n84013) );
  NAND2_X1 U69608 ( .A1(n84014), .A2(n84015), .ZN(n84006) );
  AOI22_X1 U69609 ( .A1(n105863), .A2(n108901), .B1(n83159), .B2(n108881), 
        .ZN(n84015) );
  AOI22_X1 U69610 ( .A1(n105861), .A2(n108876), .B1(n83161), .B2(n108872), 
        .ZN(n84014) );
  AND2_X2 U69611 ( .A1(n105859), .A2(n71737), .ZN(n83991) );
  AOI22_X1 U69612 ( .A1(n105857), .A2(n108865), .B1(n83164), .B2(n108878), 
        .ZN(n83989) );
  AOI22_X1 U69613 ( .A1(n83165), .A2(n108927), .B1(n83166), .B2(n108957), .ZN(
        n83988) );
  AOI22_X1 U69614 ( .A1(n106286), .A2(n108901), .B1(n71666), .B2(n106285), 
        .ZN(n83987) );
  NAND4_X2 U69615 ( .A1(n84016), .A2(n84017), .A3(n84018), .A4(n84019), .ZN(
        n58834) );
  NOR3_X1 U69616 ( .A1(n84020), .A2(n84021), .A3(n84022), .ZN(n84019) );
  NOR2_X1 U69617 ( .A1(n103374), .A2(n105166), .ZN(n84022) );
  AOI21_X1 U69618 ( .B1(n84023), .B2(n84024), .A(n106323), .ZN(n84021) );
  NOR4_X1 U69619 ( .A1(n84025), .A2(n84026), .A3(n84027), .A4(n84028), .ZN(
        n84024) );
  OAI21_X1 U69620 ( .B1(n103378), .B2(n106739), .A(n84029), .ZN(n84028) );
  AOI22_X1 U69621 ( .A1(n105884), .A2(n108774), .B1(n83123), .B2(n108779), 
        .ZN(n84029) );
  NAND2_X1 U69622 ( .A1(n84030), .A2(n84031), .ZN(n84027) );
  AOI22_X1 U69623 ( .A1(n83126), .A2(n108783), .B1(n105881), .B2(n71534), .ZN(
        n84031) );
  AOI22_X1 U69624 ( .A1(n83128), .A2(n108824), .B1(n83129), .B2(n71522), .ZN(
        n84030) );
  OAI21_X1 U69625 ( .B1(n101019), .B2(n105167), .A(n84032), .ZN(n84026) );
  AOI22_X1 U69626 ( .A1(n83131), .A2(n108811), .B1(n105877), .B2(n108795), 
        .ZN(n84032) );
  NAND2_X1 U69627 ( .A1(n84033), .A2(n84034), .ZN(n84025) );
  AOI22_X1 U69628 ( .A1(n105876), .A2(n108821), .B1(n83136), .B2(n71574), .ZN(
        n84034) );
  AOI22_X1 U69629 ( .A1(n105874), .A2(n108803), .B1(n83138), .B2(n108807), 
        .ZN(n84033) );
  NOR4_X1 U69630 ( .A1(n84035), .A2(n84036), .A3(n84037), .A4(n84038), .ZN(
        n84023) );
  OAI21_X1 U69631 ( .B1(n103389), .B2(n83143), .A(n84039), .ZN(n84038) );
  NAND2_X1 U69633 ( .A1(n84040), .A2(n84041), .ZN(n84037) );
  AOI22_X1 U69634 ( .A1(n105870), .A2(n108834), .B1(n71482), .B2(n105869), 
        .ZN(n84041) );
  AOI22_X1 U69635 ( .A1(n105868), .A2(n108837), .B1(n105867), .B2(n108772), 
        .ZN(n84040) );
  OAI21_X1 U69636 ( .B1(n103387), .B2(n105169), .A(n84042), .ZN(n84036) );
  AOI22_X1 U69637 ( .A1(n71494), .A2(n83154), .B1(n71486), .B2(n105865), .ZN(
        n84042) );
  NAND2_X1 U69638 ( .A1(n84043), .A2(n84044), .ZN(n84035) );
  AOI22_X1 U69639 ( .A1(n105863), .A2(n108789), .B1(n83159), .B2(n108769), 
        .ZN(n84044) );
  AOI22_X1 U69640 ( .A1(n105861), .A2(n108764), .B1(n83161), .B2(n108760), 
        .ZN(n84043) );
  AND2_X2 U69641 ( .A1(n105859), .A2(n71593), .ZN(n84020) );
  AOI22_X1 U69642 ( .A1(n105857), .A2(n108753), .B1(n83164), .B2(n108766), 
        .ZN(n84018) );
  AOI22_X1 U69643 ( .A1(n83165), .A2(n108815), .B1(n83166), .B2(n108845), .ZN(
        n84017) );
  AOI22_X1 U69644 ( .A1(n106289), .A2(n108789), .B1(n71522), .B2(n106285), 
        .ZN(n84016) );
  NAND4_X2 U69645 ( .A1(n84045), .A2(n84046), .A3(n84047), .A4(n84048), .ZN(
        n58833) );
  NOR3_X1 U69646 ( .A1(n84049), .A2(n84050), .A3(n84051), .ZN(n84048) );
  NOR2_X1 U69647 ( .A1(n103354), .A2(n105166), .ZN(n84051) );
  OAI21_X1 U69648 ( .B1(n84052), .B2(n84053), .A(n84054), .ZN(n83114) );
  AOI21_X1 U69649 ( .B1(n84055), .B2(n84056), .A(n106323), .ZN(n84050) );
  NOR4_X1 U69650 ( .A1(n84057), .A2(n84058), .A3(n84059), .A4(n84060), .ZN(
        n84056) );
  OAI21_X1 U69651 ( .B1(n103358), .B2(n106739), .A(n84061), .ZN(n84060) );
  AOI22_X1 U69652 ( .A1(n105884), .A2(n107314), .B1(n105883), .B2(n107319), 
        .ZN(n84061) );
  NOR2_X1 U69653 ( .A1(n84062), .A2(n107024), .ZN(n83123) );
  NOR2_X1 U69654 ( .A1(n84062), .A2(n81208), .ZN(n83122) );
  NOR2_X1 U69655 ( .A1(n84062), .A2(n107026), .ZN(n83239) );
  NAND2_X1 U69656 ( .A1(n84063), .A2(n84064), .ZN(n84059) );
  AOI22_X1 U69657 ( .A1(n105882), .A2(n107323), .B1(n69643), .B2(n105881), 
        .ZN(n84064) );
  NOR2_X1 U69658 ( .A1(n84062), .A2(n106278), .ZN(n83127) );
  NOR2_X1 U69661 ( .A1(n84066), .A2(n106278), .ZN(n83126) );
  AOI22_X1 U69662 ( .A1(n105880), .A2(n107363), .B1(n69631), .B2(n105879), 
        .ZN(n84063) );
  NOR2_X1 U69663 ( .A1(n84066), .A2(n107024), .ZN(n83129) );
  NOR2_X1 U69664 ( .A1(n84067), .A2(n62190), .ZN(n83128) );
  OAI21_X1 U69665 ( .B1(n101020), .B2(n106738), .A(n84068), .ZN(n84058) );
  AOI22_X1 U69666 ( .A1(n105878), .A2(n107351), .B1(n105877), .B2(n107335), 
        .ZN(n84068) );
  NOR2_X1 U69667 ( .A1(n84052), .A2(n81208), .ZN(n83132) );
  NOR2_X1 U69668 ( .A1(n84069), .A2(n106278), .ZN(n83131) );
  NOR2_X1 U69669 ( .A1(n84069), .A2(n81208), .ZN(n83244) );
  NAND2_X1 U69670 ( .A1(n84070), .A2(n84071), .ZN(n84057) );
  AOI22_X1 U69671 ( .A1(n105876), .A2(n107361), .B1(n83136), .B2(n69683), .ZN(
        n84071) );
  NOR2_X1 U69672 ( .A1(n84069), .A2(n107026), .ZN(n83136) );
  NOR2_X1 U69673 ( .A1(n84067), .A2(n104582), .ZN(n83135) );
  AOI22_X1 U69674 ( .A1(n105874), .A2(n107343), .B1(n105873), .B2(n107347), 
        .ZN(n84070) );
  NOR2_X1 U69675 ( .A1(n84052), .A2(n106278), .ZN(n83138) );
  NOR2_X1 U69676 ( .A1(n84069), .A2(n107024), .ZN(n83137) );
  NAND2_X1 U69677 ( .A1(n84072), .A2(n105057), .ZN(n84069) );
  NOR2_X1 U69678 ( .A1(n62190), .A2(n106697), .ZN(n84072) );
  NOR4_X1 U69679 ( .A1(n84073), .A2(n84074), .A3(n84075), .A4(n84076), .ZN(
        n84055) );
  OAI21_X1 U69680 ( .B1(n103369), .B2(n83143), .A(n84077), .ZN(n84076) );
  NOR2_X1 U69683 ( .A1(n84078), .A2(n62190), .ZN(n83145) );
  NAND2_X1 U69686 ( .A1(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ), 
        .A2(n81238), .ZN(n84067) );
  OR2_X1 U69687 ( .A1(n84080), .A2(n107024), .ZN(n83143) );
  NAND2_X1 U69688 ( .A1(n84081), .A2(n84082), .ZN(n84075) );
  AOI22_X1 U69689 ( .A1(n105870), .A2(n107199), .B1(n69591), .B2(n105869), 
        .ZN(n84082) );
  NOR2_X1 U69690 ( .A1(n84083), .A2(n81208), .ZN(n83150) );
  NOR2_X1 U69691 ( .A1(n84080), .A2(n106278), .ZN(n83149) );
  AOI22_X1 U69692 ( .A1(n105868), .A2(n107193), .B1(n105867), .B2(n107312), 
        .ZN(n84081) );
  NOR2_X1 U69693 ( .A1(n84066), .A2(n81208), .ZN(n83152) );
  NOR2_X1 U69694 ( .A1(n106740), .A2(n81228), .ZN(n83151) );
  OAI21_X1 U69695 ( .B1(n103367), .B2(n105169), .A(n84084), .ZN(n84074) );
  AOI22_X1 U69696 ( .A1(n69603), .A2(n105866), .B1(n69595), .B2(n105865), .ZN(
        n84084) );
  NOR2_X1 U69697 ( .A1(n84085), .A2(n81208), .ZN(n83155) );
  NOR2_X1 U69698 ( .A1(n84085), .A2(n107024), .ZN(n83154) );
  NOR2_X1 U69699 ( .A1(n84080), .A2(n107026), .ZN(n83256) );
  NAND2_X1 U69700 ( .A1(n84086), .A2(n104582), .ZN(n84080) );
  NAND2_X1 U69701 ( .A1(n84087), .A2(n84088), .ZN(n84073) );
  AOI22_X1 U69702 ( .A1(n105863), .A2(n107329), .B1(n105862), .B2(n107309), 
        .ZN(n84088) );
  NOR2_X1 U69703 ( .A1(n84085), .A2(n107026), .ZN(n83159) );
  NOR2_X1 U69704 ( .A1(n84066), .A2(n107026), .ZN(n83158) );
  AOI22_X1 U69707 ( .A1(n83160), .A2(n107304), .B1(n105860), .B2(n107300), 
        .ZN(n84087) );
  NOR2_X1 U69708 ( .A1(n84083), .A2(n81209), .ZN(n83161) );
  NOR2_X1 U69709 ( .A1(n84085), .A2(n81209), .ZN(n83160) );
  NAND2_X1 U69710 ( .A1(n84090), .A2(n105057), .ZN(n84085) );
  NOR2_X1 U69711 ( .A1(n62190), .A2(n84091), .ZN(n84090) );
  AND2_X2 U69712 ( .A1(n105859), .A2(n69470), .ZN(n84049) );
  OAI21_X1 U69713 ( .B1(n80203), .B2(n83254), .A(n106761), .ZN(n83162) );
  NAND2_X1 U69714 ( .A1(n84092), .A2(n84086), .ZN(n83254) );
  NOR2_X1 U69715 ( .A1(n104582), .A2(n107026), .ZN(n84092) );
  AOI22_X1 U69716 ( .A1(n105857), .A2(n107293), .B1(n105856), .B2(n107306), 
        .ZN(n84047) );
  OAI21_X1 U69717 ( .B1(n84083), .B2(n84093), .A(n106281), .ZN(n83164) );
  OAI21_X1 U69718 ( .B1(n84083), .B2(n84053), .A(n106277), .ZN(n83163) );
  NAND2_X1 U69719 ( .A1(n84094), .A2(n105057), .ZN(n84083) );
  NOR2_X1 U69720 ( .A1(n84091), .A2(n104582), .ZN(n84094) );
  AOI22_X1 U69721 ( .A1(n105855), .A2(n107355), .B1(n105854), .B2(n107177), 
        .ZN(n84046) );
  OAI21_X1 U69722 ( .B1(n81252), .B2(n106740), .A(n81253), .ZN(n83166) );
  NOR2_X1 U69723 ( .A1(n84091), .A2(n105057), .ZN(n84086) );
  OAI21_X1 U69724 ( .B1(n84052), .B2(n84093), .A(n84095), .ZN(n83165) );
  NAND2_X1 U69725 ( .A1(n81230), .A2(n106328), .ZN(n84093) );
  NAND2_X1 U69726 ( .A1(n84096), .A2(n105057), .ZN(n84052) );
  NOR2_X1 U69727 ( .A1(n104582), .A2(n106697), .ZN(n84096) );
  XOR2_X1 U69728 ( .A(n81238), .B(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ), 
        .Z(n84091) );
  AOI22_X1 U69729 ( .A1(n106287), .A2(n107329), .B1(n69631), .B2(n106283), 
        .ZN(n84045) );
  NOR4_X1 U69730 ( .A1(n84098), .A2(n84099), .A3(n84100), .A4(n84101), .ZN(
        n84097) );
  NAND2_X1 U69731 ( .A1(n84102), .A2(n84103), .ZN(n84101) );
  AOI22_X1 U69732 ( .A1(n105170), .A2(n107911), .B1(n70348), .B2(n106287), 
        .ZN(n84103) );
  AOI22_X1 U69733 ( .A1(n106284), .A2(n107880), .B1(n106275), .B2(n107861), 
        .ZN(n84102) );
  NAND2_X1 U69734 ( .A1(n84104), .A2(n84105), .ZN(n84100) );
  AOI22_X1 U69735 ( .A1(n105853), .A2(n107927), .B1(n84107), .B2(n107939), 
        .ZN(n84105) );
  AOI22_X1 U69736 ( .A1(n105099), .A2(n70316), .B1(n70364), .B2(n105175), .ZN(
        n84104) );
  NAND2_X1 U69737 ( .A1(n84108), .A2(n84109), .ZN(n84099) );
  AOI22_X1 U69738 ( .A1(n84110), .A2(n107931), .B1(n84111), .B2(n107923), .ZN(
        n84109) );
  AOI22_X1 U69739 ( .A1(n84112), .A2(n107935), .B1(n105850), .B2(n107855), 
        .ZN(n84108) );
  NAND2_X1 U69740 ( .A1(n84114), .A2(n84115), .ZN(n84098) );
  AOI21_X1 U69741 ( .B1(n70405), .B2(n84116), .A(n84117), .ZN(n84115) );
  AOI21_X1 U69742 ( .B1(n84118), .B2(n84119), .A(n106323), .ZN(n84117) );
  NOR4_X1 U69743 ( .A1(n84120), .A2(n84121), .A3(n84122), .A4(n84123), .ZN(
        n84119) );
  OAI21_X1 U69744 ( .B1(n103342), .B2(n84124), .A(n84125), .ZN(n84123) );
  AOI22_X1 U69745 ( .A1(n70348), .A2(n105848), .B1(n105847), .B2(n107889), 
        .ZN(n84125) );
  OAI21_X1 U69746 ( .B1(n103344), .B2(n84128), .A(n84129), .ZN(n84122) );
  AOI22_X1 U69747 ( .A1(n70376), .A2(n105845), .B1(n70360), .B2(n105844), .ZN(
        n84129) );
  OAI21_X1 U69748 ( .B1(n105843), .B2(n107904), .A(n84133), .ZN(n84121) );
  AOI22_X1 U69749 ( .A1(n70364), .A2(n105842), .B1(n105841), .B2(n107901), 
        .ZN(n84133) );
  NAND2_X1 U69750 ( .A1(n84136), .A2(n84137), .ZN(n84120) );
  AOI22_X1 U69751 ( .A1(n84138), .A2(n107919), .B1(n70388), .B2(n105839), .ZN(
        n84137) );
  AOI22_X1 U69752 ( .A1(n84140), .A2(n107911), .B1(n84141), .B2(n107913), .ZN(
        n84136) );
  NOR4_X1 U69753 ( .A1(n84142), .A2(n84143), .A3(n84144), .A4(n84145), .ZN(
        n84118) );
  OAI21_X1 U69754 ( .B1(n84146), .B2(n107867), .A(n84147), .ZN(n84145) );
  AOI22_X1 U69755 ( .A1(n84148), .A2(n107861), .B1(n70304), .B2(n105834), .ZN(
        n84147) );
  OAI21_X1 U69756 ( .B1(n101021), .B2(n84150), .A(n84151), .ZN(n84144) );
  AOI22_X1 U69757 ( .A1(n70312), .A2(n84152), .B1(n84153), .B2(n107858), .ZN(
        n84151) );
  OAI21_X1 U69758 ( .B1(n84154), .B2(n104583), .A(n84155), .ZN(n84143) );
  AOI22_X1 U69759 ( .A1(n70320), .A2(n84156), .B1(n70324), .B2(n84157), .ZN(
        n84155) );
  OAI21_X1 U69760 ( .B1(n101148), .B2(n105827), .A(n84159), .ZN(n84142) );
  AOI22_X1 U69761 ( .A1(n105826), .A2(n107883), .B1(n105825), .B2(n107880), 
        .ZN(n84159) );
  AOI22_X1 U69762 ( .A1(n84162), .A2(n107946), .B1(n84163), .B2(n107943), .ZN(
        n84114) );
  NOR4_X1 U69763 ( .A1(n84165), .A2(n84166), .A3(n84167), .A4(n84168), .ZN(
        n84164) );
  NAND2_X1 U69764 ( .A1(n84169), .A2(n84170), .ZN(n84168) );
  AOI22_X1 U69765 ( .A1(n106745), .A2(n108007), .B1(n70490), .B2(n106287), 
        .ZN(n84170) );
  AOI22_X1 U69766 ( .A1(n70474), .A2(n106282), .B1(n106275), .B2(n107958), 
        .ZN(n84169) );
  NAND2_X1 U69767 ( .A1(n84171), .A2(n84172), .ZN(n84167) );
  AOI22_X1 U69768 ( .A1(n105853), .A2(n108023), .B1(n84107), .B2(n108035), 
        .ZN(n84172) );
  AOI22_X1 U69769 ( .A1(n70458), .A2(n105099), .B1(n70506), .B2(n105173), .ZN(
        n84171) );
  NAND2_X1 U69770 ( .A1(n84173), .A2(n84174), .ZN(n84166) );
  AOI22_X1 U69771 ( .A1(n84110), .A2(n108027), .B1(n84111), .B2(n108019), .ZN(
        n84174) );
  AOI22_X1 U69772 ( .A1(n84112), .A2(n108031), .B1(n105850), .B2(n107952), 
        .ZN(n84173) );
  NAND2_X1 U69773 ( .A1(n84175), .A2(n84176), .ZN(n84165) );
  AOI21_X1 U69774 ( .B1(n70547), .B2(n84116), .A(n84177), .ZN(n84176) );
  AOI21_X1 U69775 ( .B1(n84178), .B2(n84179), .A(n106327), .ZN(n84177) );
  NOR4_X1 U69776 ( .A1(n84180), .A2(n84181), .A3(n84182), .A4(n84183), .ZN(
        n84179) );
  OAI21_X1 U69777 ( .B1(n105849), .B2(n104653), .A(n84184), .ZN(n84183) );
  AOI22_X1 U69778 ( .A1(n70490), .A2(n105848), .B1(n105847), .B2(n107984), 
        .ZN(n84184) );
  OAI21_X1 U69779 ( .B1(n103332), .B2(n84128), .A(n84185), .ZN(n84182) );
  AOI22_X1 U69780 ( .A1(n70518), .A2(n105845), .B1(n70502), .B2(n105844), .ZN(
        n84185) );
  OAI21_X1 U69781 ( .B1(n105843), .B2(n108000), .A(n84186), .ZN(n84181) );
  AOI22_X1 U69782 ( .A1(n70506), .A2(n105842), .B1(n105841), .B2(n107997), 
        .ZN(n84186) );
  NAND2_X1 U69783 ( .A1(n84187), .A2(n84188), .ZN(n84180) );
  AOI22_X1 U69784 ( .A1(n84138), .A2(n108016), .B1(n70530), .B2(n105839), .ZN(
        n84188) );
  AOI22_X1 U69785 ( .A1(n84140), .A2(n108007), .B1(n84141), .B2(n108009), .ZN(
        n84187) );
  NOR4_X1 U69786 ( .A1(n84189), .A2(n84190), .A3(n84191), .A4(n84192), .ZN(
        n84178) );
  OAI21_X1 U69787 ( .B1(n84146), .B2(n107964), .A(n84193), .ZN(n84192) );
  AOI22_X1 U69788 ( .A1(n84148), .A2(n107958), .B1(n70446), .B2(n105834), .ZN(
        n84193) );
  OAI21_X1 U69789 ( .B1(n101022), .B2(n84150), .A(n84194), .ZN(n84191) );
  AOI22_X1 U69790 ( .A1(n70454), .A2(n84152), .B1(n84153), .B2(n107955), .ZN(
        n84194) );
  OAI21_X1 U69791 ( .B1(n84154), .B2(n104614), .A(n84195), .ZN(n84190) );
  AOI22_X1 U69792 ( .A1(n70462), .A2(n84156), .B1(n70466), .B2(n84157), .ZN(
        n84195) );
  OAI21_X1 U69793 ( .B1(n84158), .B2(n104648), .A(n84196), .ZN(n84189) );
  AOI22_X1 U69794 ( .A1(n105826), .A2(n107978), .B1(n70474), .B2(n105825), 
        .ZN(n84196) );
  AOI22_X1 U69795 ( .A1(n84162), .A2(n108042), .B1(n84163), .B2(n108039), .ZN(
        n84175) );
  NOR4_X1 U69796 ( .A1(n84198), .A2(n84199), .A3(n84200), .A4(n84201), .ZN(
        n84197) );
  NAND2_X1 U69797 ( .A1(n84202), .A2(n84203), .ZN(n84201) );
  AOI22_X1 U69798 ( .A1(n106745), .A2(n107278), .B1(n69543), .B2(n106287), 
        .ZN(n84203) );
  AOI22_X1 U69799 ( .A1(n106284), .A2(n107242), .B1(n106275), .B2(n107220), 
        .ZN(n84202) );
  NAND2_X1 U69800 ( .A1(n84204), .A2(n84205), .ZN(n84200) );
  AOI22_X1 U69801 ( .A1(n105853), .A2(n107202), .B1(n84107), .B2(n107178), 
        .ZN(n84205) );
  AOI22_X1 U69802 ( .A1(n69511), .A2(n105101), .B1(n106746), .B2(n107266), 
        .ZN(n84204) );
  NAND2_X1 U69803 ( .A1(n84206), .A2(n84207), .ZN(n84199) );
  AOI22_X1 U69804 ( .A1(n84110), .A2(n107194), .B1(n84111), .B2(n107210), .ZN(
        n84207) );
  AOI22_X1 U69805 ( .A1(n84112), .A2(n107186), .B1(n105850), .B2(n107214), 
        .ZN(n84206) );
  NAND2_X1 U69806 ( .A1(n84208), .A2(n84209), .ZN(n84198) );
  AOI21_X1 U69807 ( .B1(n69463), .B2(n84116), .A(n84210), .ZN(n84209) );
  AOI21_X1 U69808 ( .B1(n84211), .B2(n84212), .A(n106323), .ZN(n84210) );
  NOR4_X1 U69809 ( .A1(n84213), .A2(n84214), .A3(n84215), .A4(n84216), .ZN(
        n84212) );
  OAI21_X1 U69810 ( .B1(n103316), .B2(n105849), .A(n84217), .ZN(n84216) );
  AOI22_X1 U69811 ( .A1(n69543), .A2(n105848), .B1(n105847), .B2(n107252), 
        .ZN(n84217) );
  OAI21_X1 U69812 ( .B1(n103318), .B2(n84128), .A(n84218), .ZN(n84215) );
  AOI22_X1 U69813 ( .A1(n69571), .A2(n105845), .B1(n69555), .B2(n105844), .ZN(
        n84218) );
  OAI21_X1 U69814 ( .B1(n105843), .B2(n107271), .A(n84219), .ZN(n84214) );
  AOI22_X1 U69815 ( .A1(n105842), .A2(n107266), .B1(n105841), .B2(n107268), 
        .ZN(n84219) );
  NAND2_X1 U69816 ( .A1(n84220), .A2(n84221), .ZN(n84213) );
  AOI22_X1 U69817 ( .A1(n84138), .A2(n107286), .B1(n69583), .B2(n105839), .ZN(
        n84221) );
  AOI22_X1 U69818 ( .A1(n84140), .A2(n107278), .B1(n84141), .B2(n107280), .ZN(
        n84220) );
  NOR4_X1 U69819 ( .A1(n84222), .A2(n84223), .A3(n84224), .A4(n84225), .ZN(
        n84211) );
  OAI21_X1 U69820 ( .B1(n84146), .B2(n107227), .A(n84226), .ZN(n84225) );
  AOI22_X1 U69821 ( .A1(n84148), .A2(n107220), .B1(n105834), .B2(n107223), 
        .ZN(n84226) );
  OAI21_X1 U69822 ( .B1(n101023), .B2(n84150), .A(n84227), .ZN(n84224) );
  AOI22_X1 U69823 ( .A1(n69507), .A2(n84152), .B1(n84153), .B2(n107217), .ZN(
        n84227) );
  OAI21_X1 U69824 ( .B1(n84154), .B2(n104613), .A(n84228), .ZN(n84223) );
  AOI22_X1 U69825 ( .A1(n69515), .A2(n84156), .B1(n69519), .B2(n84157), .ZN(
        n84228) );
  OAI21_X1 U69826 ( .B1(n103320), .B2(n105827), .A(n84229), .ZN(n84222) );
  AOI22_X1 U69827 ( .A1(n105826), .A2(n107245), .B1(n105825), .B2(n107242), 
        .ZN(n84229) );
  AOI22_X1 U69828 ( .A1(n84162), .A2(n106838), .B1(n84163), .B2(n107170), .ZN(
        n84208) );
  NOR4_X1 U69829 ( .A1(n84231), .A2(n84232), .A3(n84233), .A4(n84234), .ZN(
        n84230) );
  NAND2_X1 U69830 ( .A1(n84235), .A2(n84236), .ZN(n84234) );
  AOI22_X1 U69831 ( .A1(n105170), .A2(n107816), .B1(n70204), .B2(n106288), 
        .ZN(n84236) );
  AOI22_X1 U69832 ( .A1(n106284), .A2(n107781), .B1(n106275), .B2(n107758), 
        .ZN(n84235) );
  NAND2_X1 U69833 ( .A1(n84237), .A2(n84238), .ZN(n84233) );
  AOI22_X1 U69834 ( .A1(n105853), .A2(n107831), .B1(n84107), .B2(n107844), 
        .ZN(n84238) );
  AOI22_X1 U69835 ( .A1(n70172), .A2(n105099), .B1(n106746), .B2(n107803), 
        .ZN(n84237) );
  NAND2_X1 U69836 ( .A1(n84239), .A2(n84240), .ZN(n84232) );
  AOI22_X1 U69837 ( .A1(n84110), .A2(n107836), .B1(n84111), .B2(n107827), .ZN(
        n84240) );
  AOI22_X1 U69838 ( .A1(n84112), .A2(n107840), .B1(n105850), .B2(n107752), 
        .ZN(n84239) );
  NAND2_X1 U69839 ( .A1(n84241), .A2(n84242), .ZN(n84231) );
  AOI21_X1 U69840 ( .B1(n70261), .B2(n84116), .A(n84243), .ZN(n84242) );
  AOI21_X1 U69841 ( .B1(n84244), .B2(n84245), .A(n106326), .ZN(n84243) );
  NOR4_X1 U69842 ( .A1(n84246), .A2(n84247), .A3(n84248), .A4(n84249), .ZN(
        n84245) );
  OAI21_X1 U69843 ( .B1(n105849), .B2(n104652), .A(n84250), .ZN(n84249) );
  AOI22_X1 U69844 ( .A1(n70204), .A2(n105848), .B1(n105847), .B2(n107791), 
        .ZN(n84250) );
  OAI21_X1 U69845 ( .B1(n103301), .B2(n84128), .A(n84251), .ZN(n84248) );
  AOI22_X1 U69846 ( .A1(n105845), .A2(n107812), .B1(n70216), .B2(n105844), 
        .ZN(n84251) );
  OAI21_X1 U69847 ( .B1(n105843), .B2(n107808), .A(n84252), .ZN(n84247) );
  AOI22_X1 U69848 ( .A1(n105842), .A2(n107803), .B1(n105841), .B2(n107805), 
        .ZN(n84252) );
  NAND2_X1 U69849 ( .A1(n84253), .A2(n84254), .ZN(n84246) );
  AOI22_X1 U69850 ( .A1(n84138), .A2(n107824), .B1(n70244), .B2(n105839), .ZN(
        n84254) );
  AOI22_X1 U69851 ( .A1(n84140), .A2(n107816), .B1(n84141), .B2(n107818), .ZN(
        n84253) );
  NOR4_X1 U69852 ( .A1(n84255), .A2(n84256), .A3(n84257), .A4(n84258), .ZN(
        n84244) );
  OAI21_X1 U69853 ( .B1(n103307), .B2(n105836), .A(n84259), .ZN(n84258) );
  AOI22_X1 U69854 ( .A1(n84148), .A2(n107758), .B1(n105834), .B2(n107761), 
        .ZN(n84259) );
  OAI21_X1 U69855 ( .B1(n101024), .B2(n84150), .A(n84260), .ZN(n84257) );
  AOI22_X1 U69856 ( .A1(n70168), .A2(n84152), .B1(n84153), .B2(n107755), .ZN(
        n84260) );
  OAI21_X1 U69857 ( .B1(n84154), .B2(n104612), .A(n84261), .ZN(n84256) );
  AOI22_X1 U69858 ( .A1(n70176), .A2(n84156), .B1(n70180), .B2(n84157), .ZN(
        n84261) );
  OAI21_X1 U69859 ( .B1(n103303), .B2(n84158), .A(n84262), .ZN(n84255) );
  AOI22_X1 U69860 ( .A1(n105826), .A2(n107784), .B1(n105825), .B2(n107781), 
        .ZN(n84262) );
  AOI22_X1 U69861 ( .A1(n84162), .A2(n107851), .B1(n84163), .B2(n107848), .ZN(
        n84241) );
  NOR4_X1 U69862 ( .A1(n84264), .A2(n84265), .A3(n84266), .A4(n84267), .ZN(
        n84263) );
  NAND2_X1 U69863 ( .A1(n84268), .A2(n84269), .ZN(n84267) );
  AOI22_X1 U69864 ( .A1(n105170), .A2(n110712), .B1(n74050), .B2(n106289), 
        .ZN(n84269) );
  AOI22_X1 U69865 ( .A1(n106284), .A2(n110682), .B1(n106275), .B2(n110661), 
        .ZN(n84268) );
  NAND2_X1 U69866 ( .A1(n84270), .A2(n84271), .ZN(n84266) );
  AOI22_X1 U69867 ( .A1(n105853), .A2(n110727), .B1(n84107), .B2(n110739), 
        .ZN(n84271) );
  AOI22_X1 U69868 ( .A1(n74018), .A2(n105099), .B1(n105173), .B2(n110701), 
        .ZN(n84270) );
  NAND2_X1 U69869 ( .A1(n84272), .A2(n84273), .ZN(n84265) );
  AOI22_X1 U69870 ( .A1(n84110), .A2(n110731), .B1(n84111), .B2(n110723), .ZN(
        n84273) );
  AOI22_X1 U69871 ( .A1(n84112), .A2(n110735), .B1(n105850), .B2(n110655), 
        .ZN(n84272) );
  NAND2_X1 U69872 ( .A1(n84274), .A2(n84275), .ZN(n84264) );
  AOI21_X1 U69873 ( .B1(n74107), .B2(n84116), .A(n84276), .ZN(n84275) );
  AOI21_X1 U69874 ( .B1(n84277), .B2(n84278), .A(n106325), .ZN(n84276) );
  NOR4_X1 U69875 ( .A1(n84279), .A2(n84280), .A3(n84281), .A4(n84282), .ZN(
        n84278) );
  OAI21_X1 U69876 ( .B1(n103282), .B2(n105849), .A(n84283), .ZN(n84282) );
  AOI22_X1 U69877 ( .A1(n74050), .A2(n105848), .B1(n105847), .B2(n110691), 
        .ZN(n84283) );
  OAI21_X1 U69878 ( .B1(n103284), .B2(n84128), .A(n84284), .ZN(n84281) );
  AOI22_X1 U69879 ( .A1(n105845), .A2(n110708), .B1(n74062), .B2(n105844), 
        .ZN(n84284) );
  OAI21_X1 U69880 ( .B1(n103280), .B2(n105843), .A(n84285), .ZN(n84280) );
  AOI22_X1 U69881 ( .A1(n105842), .A2(n110701), .B1(n105841), .B2(n110702), 
        .ZN(n84285) );
  NAND2_X1 U69882 ( .A1(n84286), .A2(n84287), .ZN(n84279) );
  AOI22_X1 U69883 ( .A1(n84138), .A2(n110720), .B1(n74090), .B2(n105839), .ZN(
        n84287) );
  AOI22_X1 U69884 ( .A1(n84140), .A2(n110712), .B1(n84141), .B2(n110714), .ZN(
        n84286) );
  NOR4_X1 U69885 ( .A1(n84288), .A2(n84289), .A3(n84290), .A4(n84291), .ZN(
        n84277) );
  OAI21_X1 U69886 ( .B1(n103290), .B2(n84146), .A(n84292), .ZN(n84291) );
  AOI22_X1 U69887 ( .A1(n84148), .A2(n110661), .B1(n105834), .B2(n110664), 
        .ZN(n84292) );
  OAI21_X1 U69888 ( .B1(n101025), .B2(n84150), .A(n84293), .ZN(n84290) );
  AOI22_X1 U69889 ( .A1(n74014), .A2(n84152), .B1(n84153), .B2(n110658), .ZN(
        n84293) );
  OAI21_X1 U69890 ( .B1(n84154), .B2(n104611), .A(n84294), .ZN(n84289) );
  AOI22_X1 U69891 ( .A1(n74022), .A2(n84156), .B1(n74026), .B2(n84157), .ZN(
        n84294) );
  OAI21_X1 U69892 ( .B1(n103286), .B2(n105827), .A(n84295), .ZN(n84288) );
  AOI22_X1 U69893 ( .A1(n105826), .A2(n110685), .B1(n105825), .B2(n110682), 
        .ZN(n84295) );
  AOI22_X1 U69894 ( .A1(n84162), .A2(n110746), .B1(n84163), .B2(n110743), .ZN(
        n84274) );
  NOR4_X1 U69895 ( .A1(n84297), .A2(n84298), .A3(n84299), .A4(n84300), .ZN(
        n84296) );
  NAND2_X1 U69896 ( .A1(n84301), .A2(n84302), .ZN(n84300) );
  AOI22_X1 U69897 ( .A1(n105170), .A2(n108115), .B1(n70637), .B2(n106287), 
        .ZN(n84302) );
  AOI22_X1 U69898 ( .A1(n106284), .A2(n108082), .B1(n106275), .B2(n108060), 
        .ZN(n84301) );
  NAND2_X1 U69899 ( .A1(n84303), .A2(n84304), .ZN(n84299) );
  AOI22_X1 U69900 ( .A1(n105853), .A2(n108131), .B1(n84107), .B2(n108144), 
        .ZN(n84304) );
  AOI22_X1 U69901 ( .A1(n70605), .A2(n105099), .B1(n105174), .B2(n108104), 
        .ZN(n84303) );
  NAND2_X1 U69902 ( .A1(n84305), .A2(n84306), .ZN(n84298) );
  AOI22_X1 U69903 ( .A1(n84110), .A2(n108136), .B1(n84111), .B2(n108127), .ZN(
        n84306) );
  AOI22_X1 U69904 ( .A1(n84112), .A2(n108140), .B1(n105850), .B2(n108054), 
        .ZN(n84305) );
  NAND2_X1 U69905 ( .A1(n84307), .A2(n84308), .ZN(n84297) );
  AOI21_X1 U69906 ( .B1(n70694), .B2(n84116), .A(n84309), .ZN(n84308) );
  AOI21_X1 U69907 ( .B1(n84310), .B2(n84311), .A(n106324), .ZN(n84309) );
  NOR4_X1 U69908 ( .A1(n84312), .A2(n84313), .A3(n84314), .A4(n84315), .ZN(
        n84311) );
  OAI21_X1 U69909 ( .B1(n103263), .B2(n105849), .A(n84316), .ZN(n84315) );
  AOI22_X1 U69910 ( .A1(n70637), .A2(n105848), .B1(n105847), .B2(n108091), 
        .ZN(n84316) );
  OAI21_X1 U69911 ( .B1(n103265), .B2(n84128), .A(n84317), .ZN(n84314) );
  AOI22_X1 U69912 ( .A1(n105845), .A2(n108111), .B1(n70649), .B2(n105844), 
        .ZN(n84317) );
  OAI21_X1 U69913 ( .B1(n103261), .B2(n105843), .A(n84318), .ZN(n84313) );
  AOI22_X1 U69914 ( .A1(n105842), .A2(n108104), .B1(n105841), .B2(n108105), 
        .ZN(n84318) );
  NAND2_X1 U69915 ( .A1(n84319), .A2(n84320), .ZN(n84312) );
  AOI22_X1 U69916 ( .A1(n84138), .A2(n108123), .B1(n70677), .B2(n105839), .ZN(
        n84320) );
  AOI22_X1 U69917 ( .A1(n84140), .A2(n108115), .B1(n84141), .B2(n108117), .ZN(
        n84319) );
  NOR4_X1 U69918 ( .A1(n84321), .A2(n84322), .A3(n84323), .A4(n84324), .ZN(
        n84310) );
  OAI21_X1 U69919 ( .B1(n103271), .B2(n105836), .A(n84325), .ZN(n84324) );
  AOI22_X1 U69920 ( .A1(n84148), .A2(n108060), .B1(n105834), .B2(n108063), 
        .ZN(n84325) );
  OAI21_X1 U69921 ( .B1(n101026), .B2(n84150), .A(n84326), .ZN(n84323) );
  AOI22_X1 U69922 ( .A1(n70601), .A2(n84152), .B1(n84153), .B2(n108057), .ZN(
        n84326) );
  OAI21_X1 U69923 ( .B1(n84154), .B2(n104610), .A(n84327), .ZN(n84322) );
  AOI22_X1 U69924 ( .A1(n70609), .A2(n84156), .B1(n70613), .B2(n84157), .ZN(
        n84327) );
  OAI21_X1 U69925 ( .B1(n103267), .B2(n84158), .A(n84328), .ZN(n84321) );
  AOI22_X1 U69926 ( .A1(n105826), .A2(n108085), .B1(n105825), .B2(n108082), 
        .ZN(n84328) );
  AOI22_X1 U69927 ( .A1(n84162), .A2(n108151), .B1(n84163), .B2(n108148), .ZN(
        n84307) );
  NOR4_X1 U69928 ( .A1(n84330), .A2(n84331), .A3(n84332), .A4(n84333), .ZN(
        n84329) );
  NAND2_X1 U69929 ( .A1(n84334), .A2(n84335), .ZN(n84333) );
  AOI22_X1 U69930 ( .A1(n105170), .A2(n110814), .B1(n74191), .B2(n106286), 
        .ZN(n84335) );
  AOI22_X1 U69931 ( .A1(n106283), .A2(n110780), .B1(n106275), .B2(n110758), 
        .ZN(n84334) );
  NAND2_X1 U69932 ( .A1(n84336), .A2(n84337), .ZN(n84332) );
  AOI22_X1 U69933 ( .A1(n105853), .A2(n110830), .B1(n84107), .B2(n110842), 
        .ZN(n84337) );
  AOI22_X1 U69934 ( .A1(n74159), .A2(n105101), .B1(n105173), .B2(n110803), 
        .ZN(n84336) );
  NAND2_X1 U69935 ( .A1(n84338), .A2(n84339), .ZN(n84331) );
  AOI22_X1 U69936 ( .A1(n84110), .A2(n110834), .B1(n84111), .B2(n110826), .ZN(
        n84339) );
  AOI22_X1 U69937 ( .A1(n84112), .A2(n110838), .B1(n105850), .B2(n110752), 
        .ZN(n84338) );
  NAND2_X1 U69938 ( .A1(n84340), .A2(n84341), .ZN(n84330) );
  AOI21_X1 U69939 ( .B1(n74248), .B2(n84116), .A(n84342), .ZN(n84341) );
  AOI21_X1 U69940 ( .B1(n84343), .B2(n84344), .A(n106324), .ZN(n84342) );
  NOR4_X1 U69941 ( .A1(n84345), .A2(n84346), .A3(n84347), .A4(n84348), .ZN(
        n84344) );
  OAI21_X1 U69942 ( .B1(n103244), .B2(n105849), .A(n84349), .ZN(n84348) );
  AOI22_X1 U69943 ( .A1(n74191), .A2(n105848), .B1(n105847), .B2(n110790), 
        .ZN(n84349) );
  OAI21_X1 U69944 ( .B1(n103246), .B2(n84128), .A(n84350), .ZN(n84347) );
  AOI22_X1 U69945 ( .A1(n105845), .A2(n110810), .B1(n74203), .B2(n105844), 
        .ZN(n84350) );
  OAI21_X1 U69946 ( .B1(n103242), .B2(n105843), .A(n84351), .ZN(n84346) );
  AOI22_X1 U69947 ( .A1(n105842), .A2(n110803), .B1(n105841), .B2(n110804), 
        .ZN(n84351) );
  NAND2_X1 U69948 ( .A1(n84352), .A2(n84353), .ZN(n84345) );
  AOI22_X1 U69949 ( .A1(n84138), .A2(n110822), .B1(n74231), .B2(n105839), .ZN(
        n84353) );
  AOI22_X1 U69950 ( .A1(n84140), .A2(n110814), .B1(n84141), .B2(n110816), .ZN(
        n84352) );
  NOR4_X1 U69951 ( .A1(n84354), .A2(n84355), .A3(n84356), .A4(n84357), .ZN(
        n84343) );
  OAI21_X1 U69952 ( .B1(n103252), .B2(n84146), .A(n84358), .ZN(n84357) );
  AOI22_X1 U69953 ( .A1(n84148), .A2(n110758), .B1(n105834), .B2(n110761), 
        .ZN(n84358) );
  OAI21_X1 U69954 ( .B1(n101027), .B2(n84150), .A(n84359), .ZN(n84356) );
  AOI22_X1 U69955 ( .A1(n74155), .A2(n84152), .B1(n84153), .B2(n110755), .ZN(
        n84359) );
  OAI21_X1 U69956 ( .B1(n84154), .B2(n104609), .A(n84360), .ZN(n84355) );
  AOI22_X1 U69957 ( .A1(n74163), .A2(n84156), .B1(n74167), .B2(n84157), .ZN(
        n84360) );
  OAI21_X1 U69958 ( .B1(n103248), .B2(n105827), .A(n84361), .ZN(n84354) );
  AOI22_X1 U69959 ( .A1(n105826), .A2(n110783), .B1(n105825), .B2(n110780), 
        .ZN(n84361) );
  AOI22_X1 U69960 ( .A1(n84162), .A2(n110849), .B1(n84163), .B2(n110846), .ZN(
        n84340) );
  NOR4_X1 U69961 ( .A1(n84363), .A2(n84364), .A3(n84365), .A4(n84366), .ZN(
        n84362) );
  NAND2_X1 U69962 ( .A1(n84367), .A2(n84368), .ZN(n84366) );
  AOI22_X1 U69963 ( .A1(n105171), .A2(n110914), .B1(n74331), .B2(n80259), .ZN(
        n84368) );
  AOI22_X1 U69964 ( .A1(n106284), .A2(n110881), .B1(n106275), .B2(n110859), 
        .ZN(n84367) );
  NAND2_X1 U69965 ( .A1(n84369), .A2(n84370), .ZN(n84365) );
  AOI22_X1 U69966 ( .A1(n105853), .A2(n110931), .B1(n84107), .B2(n110943), 
        .ZN(n84370) );
  AOI22_X1 U69967 ( .A1(n74299), .A2(n105099), .B1(n106746), .B2(n110900), 
        .ZN(n84369) );
  NAND2_X1 U69968 ( .A1(n84371), .A2(n84372), .ZN(n84364) );
  AOI22_X1 U69969 ( .A1(n84110), .A2(n110935), .B1(n84111), .B2(n110927), .ZN(
        n84372) );
  AOI22_X1 U69970 ( .A1(n84112), .A2(n110939), .B1(n105850), .B2(n110853), 
        .ZN(n84371) );
  NAND2_X1 U69971 ( .A1(n84373), .A2(n84374), .ZN(n84363) );
  AOI21_X1 U69972 ( .B1(n74388), .B2(n84116), .A(n84375), .ZN(n84374) );
  AOI21_X1 U69973 ( .B1(n84376), .B2(n84377), .A(n106325), .ZN(n84375) );
  NOR4_X1 U69974 ( .A1(n84378), .A2(n84379), .A3(n84380), .A4(n84381), .ZN(
        n84377) );
  OAI21_X1 U69975 ( .B1(n103225), .B2(n105849), .A(n84382), .ZN(n84381) );
  AOI22_X1 U69976 ( .A1(n74331), .A2(n105848), .B1(n105847), .B2(n110890), 
        .ZN(n84382) );
  OAI21_X1 U69977 ( .B1(n103227), .B2(n84128), .A(n84383), .ZN(n84380) );
  AOI22_X1 U69978 ( .A1(n105845), .A2(n110910), .B1(n74343), .B2(n105844), 
        .ZN(n84383) );
  OAI21_X1 U69979 ( .B1(n103223), .B2(n105843), .A(n84384), .ZN(n84379) );
  AOI22_X1 U69980 ( .A1(n105842), .A2(n110900), .B1(n105841), .B2(n110902), 
        .ZN(n84384) );
  NAND2_X1 U69981 ( .A1(n84385), .A2(n84386), .ZN(n84378) );
  AOI22_X1 U69982 ( .A1(n84138), .A2(n110923), .B1(n74371), .B2(n105839), .ZN(
        n84386) );
  AOI22_X1 U69983 ( .A1(n84140), .A2(n110914), .B1(n84141), .B2(n110916), .ZN(
        n84385) );
  NOR4_X1 U69984 ( .A1(n84387), .A2(n84388), .A3(n84389), .A4(n84390), .ZN(
        n84376) );
  OAI21_X1 U69985 ( .B1(n103233), .B2(n105836), .A(n84391), .ZN(n84390) );
  AOI22_X1 U69986 ( .A1(n84148), .A2(n110859), .B1(n105834), .B2(n110862), 
        .ZN(n84391) );
  OAI21_X1 U69987 ( .B1(n101028), .B2(n84150), .A(n84392), .ZN(n84389) );
  AOI22_X1 U69988 ( .A1(n74295), .A2(n84152), .B1(n84153), .B2(n110856), .ZN(
        n84392) );
  OAI21_X1 U69989 ( .B1(n84154), .B2(n104608), .A(n84393), .ZN(n84388) );
  AOI22_X1 U69990 ( .A1(n74303), .A2(n84156), .B1(n74307), .B2(n84157), .ZN(
        n84393) );
  OAI21_X1 U69991 ( .B1(n103229), .B2(n84158), .A(n84394), .ZN(n84387) );
  AOI22_X1 U69992 ( .A1(n74319), .A2(n105826), .B1(n105825), .B2(n110881), 
        .ZN(n84394) );
  AOI22_X1 U69993 ( .A1(n84162), .A2(n110950), .B1(n84163), .B2(n110947), .ZN(
        n84373) );
  NOR4_X1 U69994 ( .A1(n84396), .A2(n84397), .A3(n84398), .A4(n84399), .ZN(
        n84395) );
  NAND2_X1 U69995 ( .A1(n84400), .A2(n84401), .ZN(n84399) );
  AOI22_X1 U69996 ( .A1(n105172), .A2(n110509), .B1(n73767), .B2(n106288), 
        .ZN(n84401) );
  AOI22_X1 U69997 ( .A1(n106284), .A2(n110475), .B1(n106275), .B2(n110454), 
        .ZN(n84400) );
  NAND2_X1 U69998 ( .A1(n84402), .A2(n84403), .ZN(n84398) );
  AOI22_X1 U69999 ( .A1(n105853), .A2(n110524), .B1(n84107), .B2(n110536), 
        .ZN(n84403) );
  AOI22_X1 U70000 ( .A1(n73735), .A2(n105099), .B1(n105173), .B2(n110495), 
        .ZN(n84402) );
  NAND2_X1 U70001 ( .A1(n84404), .A2(n84405), .ZN(n84397) );
  AOI22_X1 U70002 ( .A1(n84110), .A2(n110528), .B1(n84111), .B2(n110520), .ZN(
        n84405) );
  AOI22_X1 U70003 ( .A1(n84112), .A2(n110532), .B1(n84113), .B2(n110448), .ZN(
        n84404) );
  NAND2_X1 U70004 ( .A1(n84406), .A2(n84407), .ZN(n84396) );
  AOI21_X1 U70005 ( .B1(n73824), .B2(n84116), .A(n84408), .ZN(n84407) );
  AOI21_X1 U70006 ( .B1(n84409), .B2(n84410), .A(n106326), .ZN(n84408) );
  NOR4_X1 U70007 ( .A1(n84411), .A2(n84412), .A3(n84413), .A4(n84414), .ZN(
        n84410) );
  OAI21_X1 U70008 ( .B1(n103207), .B2(n105849), .A(n84415), .ZN(n84414) );
  AOI22_X1 U70009 ( .A1(n73767), .A2(n84126), .B1(n105847), .B2(n110484), .ZN(
        n84415) );
  OAI21_X1 U70010 ( .B1(n103209), .B2(n84128), .A(n84416), .ZN(n84413) );
  AOI22_X1 U70011 ( .A1(n105845), .A2(n110505), .B1(n73779), .B2(n105844), 
        .ZN(n84416) );
  OAI21_X1 U70012 ( .B1(n103205), .B2(n105843), .A(n84417), .ZN(n84412) );
  AOI22_X1 U70013 ( .A1(n105842), .A2(n110495), .B1(n105841), .B2(n110497), 
        .ZN(n84417) );
  NAND2_X1 U70014 ( .A1(n84418), .A2(n84419), .ZN(n84411) );
  AOI22_X1 U70015 ( .A1(n84138), .A2(n110517), .B1(n73807), .B2(n105839), .ZN(
        n84419) );
  AOI22_X1 U70016 ( .A1(n84140), .A2(n110509), .B1(n84141), .B2(n110511), .ZN(
        n84418) );
  NOR4_X1 U70017 ( .A1(n84420), .A2(n84421), .A3(n84422), .A4(n84423), .ZN(
        n84409) );
  OAI21_X1 U70018 ( .B1(n103214), .B2(n84146), .A(n84424), .ZN(n84423) );
  AOI22_X1 U70019 ( .A1(n84148), .A2(n110454), .B1(n105834), .B2(n110457), 
        .ZN(n84424) );
  OAI21_X1 U70020 ( .B1(n101029), .B2(n84150), .A(n84425), .ZN(n84422) );
  AOI22_X1 U70021 ( .A1(n73731), .A2(n84152), .B1(n84153), .B2(n110451), .ZN(
        n84425) );
  OAI21_X1 U70022 ( .B1(n84154), .B2(n104607), .A(n84426), .ZN(n84421) );
  AOI22_X1 U70023 ( .A1(n73739), .A2(n84156), .B1(n73743), .B2(n84157), .ZN(
        n84426) );
  OAI21_X1 U70024 ( .B1(n103211), .B2(n105827), .A(n84427), .ZN(n84420) );
  AOI22_X1 U70025 ( .A1(n105826), .A2(n110478), .B1(n105825), .B2(n110475), 
        .ZN(n84427) );
  AOI22_X1 U70026 ( .A1(n84162), .A2(n110543), .B1(n84163), .B2(n110540), .ZN(
        n84406) );
  NOR4_X1 U70027 ( .A1(n84429), .A2(n84430), .A3(n84431), .A4(n84432), .ZN(
        n84428) );
  NAND2_X1 U70028 ( .A1(n84433), .A2(n84434), .ZN(n84432) );
  AOI22_X1 U70029 ( .A1(n106745), .A2(n110292), .B1(n73471), .B2(n106286), 
        .ZN(n84434) );
  AOI22_X1 U70030 ( .A1(n106284), .A2(n110257), .B1(n106275), .B2(n110236), 
        .ZN(n84433) );
  NAND2_X1 U70031 ( .A1(n84435), .A2(n84436), .ZN(n84431) );
  AOI22_X1 U70032 ( .A1(n105853), .A2(n110309), .B1(n84107), .B2(n110321), 
        .ZN(n84436) );
  AOI22_X1 U70033 ( .A1(n73439), .A2(n105099), .B1(n105173), .B2(n110279), 
        .ZN(n84435) );
  NAND2_X1 U70034 ( .A1(n84437), .A2(n84438), .ZN(n84430) );
  AOI22_X1 U70035 ( .A1(n84110), .A2(n110313), .B1(n84111), .B2(n110305), .ZN(
        n84438) );
  AOI22_X1 U70036 ( .A1(n84112), .A2(n110317), .B1(n84113), .B2(n110231), .ZN(
        n84437) );
  NAND2_X1 U70037 ( .A1(n84439), .A2(n84440), .ZN(n84429) );
  AOI21_X1 U70038 ( .B1(n73528), .B2(n84116), .A(n84441), .ZN(n84440) );
  AOI21_X1 U70039 ( .B1(n84442), .B2(n84443), .A(n106326), .ZN(n84441) );
  NOR4_X1 U70040 ( .A1(n84444), .A2(n84445), .A3(n84446), .A4(n84447), .ZN(
        n84443) );
  OAI21_X1 U70041 ( .B1(n103188), .B2(n105849), .A(n84448), .ZN(n84447) );
  AOI22_X1 U70042 ( .A1(n73471), .A2(n84126), .B1(n105847), .B2(n110266), .ZN(
        n84448) );
  OAI21_X1 U70043 ( .B1(n103190), .B2(n84128), .A(n84449), .ZN(n84446) );
  AOI22_X1 U70044 ( .A1(n105845), .A2(n110288), .B1(n73483), .B2(n105844), 
        .ZN(n84449) );
  OAI21_X1 U70045 ( .B1(n103186), .B2(n105843), .A(n84450), .ZN(n84445) );
  AOI22_X1 U70046 ( .A1(n105842), .A2(n110279), .B1(n105841), .B2(n110280), 
        .ZN(n84450) );
  NAND2_X1 U70047 ( .A1(n84451), .A2(n84452), .ZN(n84444) );
  AOI22_X1 U70048 ( .A1(n84138), .A2(n110301), .B1(n73511), .B2(n105839), .ZN(
        n84452) );
  AOI22_X1 U70049 ( .A1(n84140), .A2(n110292), .B1(n84141), .B2(n110294), .ZN(
        n84451) );
  NOR4_X1 U70050 ( .A1(n84453), .A2(n84454), .A3(n84455), .A4(n84456), .ZN(
        n84442) );
  OAI21_X1 U70051 ( .B1(n103196), .B2(n84146), .A(n84457), .ZN(n84456) );
  AOI22_X1 U70052 ( .A1(n84148), .A2(n110236), .B1(n105834), .B2(n110239), 
        .ZN(n84457) );
  OAI21_X1 U70053 ( .B1(n101030), .B2(n84150), .A(n84458), .ZN(n84455) );
  AOI22_X1 U70054 ( .A1(n73435), .A2(n84152), .B1(n84153), .B2(n110233), .ZN(
        n84458) );
  OAI21_X1 U70055 ( .B1(n84154), .B2(n104606), .A(n84459), .ZN(n84454) );
  AOI22_X1 U70056 ( .A1(n73443), .A2(n84156), .B1(n73447), .B2(n84157), .ZN(
        n84459) );
  OAI21_X1 U70057 ( .B1(n103192), .B2(n84158), .A(n84460), .ZN(n84453) );
  AOI22_X1 U70058 ( .A1(n105826), .A2(n110260), .B1(n105825), .B2(n110257), 
        .ZN(n84460) );
  AOI22_X1 U70059 ( .A1(n84162), .A2(n110328), .B1(n84163), .B2(n110325), .ZN(
        n84439) );
  NOR4_X1 U70060 ( .A1(n84462), .A2(n84463), .A3(n84464), .A4(n84465), .ZN(
        n84461) );
  NAND2_X1 U70061 ( .A1(n84466), .A2(n84467), .ZN(n84465) );
  AOI22_X1 U70062 ( .A1(n105171), .A2(n110612), .B1(n73908), .B2(n106289), 
        .ZN(n84467) );
  AOI22_X1 U70063 ( .A1(n106283), .A2(n110574), .B1(n106275), .B2(n110553), 
        .ZN(n84466) );
  NAND2_X1 U70064 ( .A1(n84468), .A2(n84469), .ZN(n84464) );
  AOI22_X1 U70065 ( .A1(n105853), .A2(n110629), .B1(n84107), .B2(n110641), 
        .ZN(n84469) );
  AOI22_X1 U70066 ( .A1(n73876), .A2(n105100), .B1(n105174), .B2(n110598), 
        .ZN(n84468) );
  NAND2_X1 U70067 ( .A1(n84470), .A2(n84471), .ZN(n84463) );
  AOI22_X1 U70068 ( .A1(n84110), .A2(n110633), .B1(n84111), .B2(n110625), .ZN(
        n84471) );
  AOI22_X1 U70069 ( .A1(n84112), .A2(n110637), .B1(n84113), .B2(n110548), .ZN(
        n84470) );
  NAND2_X1 U70070 ( .A1(n84472), .A2(n84473), .ZN(n84462) );
  AOI21_X1 U70071 ( .B1(n73965), .B2(n84116), .A(n84474), .ZN(n84473) );
  AOI21_X1 U70072 ( .B1(n84475), .B2(n84476), .A(n106327), .ZN(n84474) );
  NOR4_X1 U70073 ( .A1(n84477), .A2(n84478), .A3(n84479), .A4(n84480), .ZN(
        n84476) );
  OAI21_X1 U70074 ( .B1(n103169), .B2(n105849), .A(n84481), .ZN(n84480) );
  AOI22_X1 U70075 ( .A1(n73908), .A2(n84126), .B1(n105847), .B2(n110584), .ZN(
        n84481) );
  OAI21_X1 U70076 ( .B1(n103171), .B2(n84128), .A(n84482), .ZN(n84479) );
  AOI22_X1 U70077 ( .A1(n105845), .A2(n110608), .B1(n73920), .B2(n105844), 
        .ZN(n84482) );
  OAI21_X1 U70078 ( .B1(n103167), .B2(n105843), .A(n84483), .ZN(n84478) );
  AOI22_X1 U70079 ( .A1(n105842), .A2(n110598), .B1(n105841), .B2(n110600), 
        .ZN(n84483) );
  NAND2_X1 U70080 ( .A1(n84484), .A2(n84485), .ZN(n84477) );
  AOI22_X1 U70081 ( .A1(n84138), .A2(n110622), .B1(n84139), .B2(n110618), .ZN(
        n84485) );
  AOI22_X1 U70082 ( .A1(n84140), .A2(n110612), .B1(n84141), .B2(n110614), .ZN(
        n84484) );
  NOR4_X1 U70083 ( .A1(n84486), .A2(n84487), .A3(n84488), .A4(n84489), .ZN(
        n84475) );
  OAI21_X1 U70084 ( .B1(n103177), .B2(n84146), .A(n84490), .ZN(n84489) );
  AOI22_X1 U70085 ( .A1(n84148), .A2(n110553), .B1(n105834), .B2(n110556), 
        .ZN(n84490) );
  OAI21_X1 U70086 ( .B1(n101031), .B2(n84150), .A(n84491), .ZN(n84488) );
  AOI22_X1 U70087 ( .A1(n73872), .A2(n84152), .B1(n84153), .B2(n110550), .ZN(
        n84491) );
  OAI21_X1 U70088 ( .B1(n84154), .B2(n104605), .A(n84492), .ZN(n84487) );
  AOI22_X1 U70089 ( .A1(n73880), .A2(n84156), .B1(n73884), .B2(n84157), .ZN(
        n84492) );
  OAI21_X1 U70090 ( .B1(n103173), .B2(n105827), .A(n84493), .ZN(n84486) );
  AOI22_X1 U70091 ( .A1(n105826), .A2(n110577), .B1(n105825), .B2(n110574), 
        .ZN(n84493) );
  AOI22_X1 U70092 ( .A1(n84162), .A2(n110648), .B1(n84163), .B2(n110645), .ZN(
        n84472) );
  NOR4_X1 U70093 ( .A1(n84495), .A2(n84496), .A3(n84497), .A4(n84498), .ZN(
        n84494) );
  NAND2_X1 U70094 ( .A1(n84499), .A2(n84500), .ZN(n84498) );
  AOI22_X1 U70095 ( .A1(n105170), .A2(n110401), .B1(n73620), .B2(n106288), 
        .ZN(n84500) );
  AOI22_X1 U70096 ( .A1(n106284), .A2(n110365), .B1(n106276), .B2(n110344), 
        .ZN(n84499) );
  NAND2_X1 U70097 ( .A1(n84501), .A2(n84502), .ZN(n84497) );
  AOI22_X1 U70098 ( .A1(n105853), .A2(n110418), .B1(n105852), .B2(n110430), 
        .ZN(n84502) );
  AOI22_X1 U70099 ( .A1(n73588), .A2(n105099), .B1(n106746), .B2(n110388), 
        .ZN(n84501) );
  NAND2_X1 U70100 ( .A1(n84503), .A2(n84504), .ZN(n84496) );
  AOI22_X1 U70101 ( .A1(n105851), .A2(n110422), .B1(n84111), .B2(n110414), 
        .ZN(n84504) );
  AOI22_X1 U70102 ( .A1(n84112), .A2(n110426), .B1(n84113), .B2(n110339), .ZN(
        n84503) );
  NAND2_X1 U70103 ( .A1(n84505), .A2(n84506), .ZN(n84495) );
  AOI21_X1 U70104 ( .B1(n73677), .B2(n84116), .A(n84507), .ZN(n84506) );
  AOI21_X1 U70105 ( .B1(n84508), .B2(n84509), .A(n106323), .ZN(n84507) );
  NOR4_X1 U70106 ( .A1(n84510), .A2(n84511), .A3(n84512), .A4(n84513), .ZN(
        n84509) );
  OAI21_X1 U70107 ( .B1(n103149), .B2(n105849), .A(n84514), .ZN(n84513) );
  AOI22_X1 U70108 ( .A1(n73620), .A2(n84126), .B1(n105847), .B2(n110375), .ZN(
        n84514) );
  OAI21_X1 U70109 ( .B1(n103151), .B2(n84128), .A(n84515), .ZN(n84512) );
  AOI22_X1 U70110 ( .A1(n105845), .A2(n110397), .B1(n73632), .B2(n105844), 
        .ZN(n84515) );
  OAI21_X1 U70111 ( .B1(n103147), .B2(n105843), .A(n84516), .ZN(n84511) );
  AOI22_X1 U70112 ( .A1(n105842), .A2(n110388), .B1(n105841), .B2(n110389), 
        .ZN(n84516) );
  NAND2_X1 U70113 ( .A1(n84517), .A2(n84518), .ZN(n84510) );
  AOI22_X1 U70114 ( .A1(n105840), .A2(n110410), .B1(n73660), .B2(n105839), 
        .ZN(n84518) );
  AOI22_X1 U70115 ( .A1(n105838), .A2(n110401), .B1(n84141), .B2(n110403), 
        .ZN(n84517) );
  NOR4_X1 U70116 ( .A1(n84519), .A2(n84520), .A3(n84521), .A4(n84522), .ZN(
        n84508) );
  OAI21_X1 U70117 ( .B1(n103158), .B2(n84146), .A(n84523), .ZN(n84522) );
  AOI22_X1 U70118 ( .A1(n105835), .A2(n110344), .B1(n105834), .B2(n110347), 
        .ZN(n84523) );
  OAI21_X1 U70119 ( .B1(n101032), .B2(n84150), .A(n84524), .ZN(n84521) );
  AOI22_X1 U70120 ( .A1(n73584), .A2(n105832), .B1(n84153), .B2(n110341), .ZN(
        n84524) );
  OAI21_X1 U70121 ( .B1(n84154), .B2(n104604), .A(n84525), .ZN(n84520) );
  AOI22_X1 U70122 ( .A1(n73592), .A2(n105829), .B1(n73596), .B2(n105828), .ZN(
        n84525) );
  OAI21_X1 U70123 ( .B1(n103154), .B2(n84158), .A(n84526), .ZN(n84519) );
  AOI22_X1 U70124 ( .A1(n105826), .A2(n110368), .B1(n105825), .B2(n110365), 
        .ZN(n84526) );
  AOI22_X1 U70125 ( .A1(n84162), .A2(n110437), .B1(n84163), .B2(n110434), .ZN(
        n84505) );
  NOR4_X1 U70126 ( .A1(n84528), .A2(n84529), .A3(n84530), .A4(n84531), .ZN(
        n84527) );
  NAND2_X1 U70127 ( .A1(n84532), .A2(n84533), .ZN(n84531) );
  AOI22_X1 U70128 ( .A1(n105171), .A2(n110079), .B1(n73182), .B2(n106288), 
        .ZN(n84533) );
  AOI22_X1 U70129 ( .A1(n106283), .A2(n110041), .B1(n106276), .B2(n110019), 
        .ZN(n84532) );
  NAND2_X1 U70130 ( .A1(n84534), .A2(n84535), .ZN(n84530) );
  AOI22_X1 U70131 ( .A1(n105853), .A2(n110096), .B1(n105852), .B2(n110108), 
        .ZN(n84535) );
  AOI22_X1 U70132 ( .A1(n73150), .A2(n105100), .B1(n105173), .B2(n110066), 
        .ZN(n84534) );
  NAND2_X1 U70133 ( .A1(n84536), .A2(n84537), .ZN(n84529) );
  AOI22_X1 U70134 ( .A1(n105851), .A2(n110100), .B1(n84111), .B2(n110092), 
        .ZN(n84537) );
  AOI22_X1 U70135 ( .A1(n84112), .A2(n110104), .B1(n84113), .B2(n110013), .ZN(
        n84536) );
  NAND2_X1 U70136 ( .A1(n84538), .A2(n84539), .ZN(n84528) );
  AOI21_X1 U70137 ( .B1(n73239), .B2(n84116), .A(n84540), .ZN(n84539) );
  AOI21_X1 U70138 ( .B1(n84541), .B2(n84542), .A(n106324), .ZN(n84540) );
  NOR4_X1 U70139 ( .A1(n84543), .A2(n84544), .A3(n84545), .A4(n84546), .ZN(
        n84542) );
  OAI21_X1 U70140 ( .B1(n103131), .B2(n84124), .A(n84547), .ZN(n84546) );
  AOI22_X1 U70141 ( .A1(n73182), .A2(n84126), .B1(n105847), .B2(n110051), .ZN(
        n84547) );
  OAI21_X1 U70142 ( .B1(n103133), .B2(n105846), .A(n84548), .ZN(n84545) );
  AOI22_X1 U70143 ( .A1(n105845), .A2(n110075), .B1(n73194), .B2(n105844), 
        .ZN(n84548) );
  OAI21_X1 U70144 ( .B1(n103129), .B2(n84132), .A(n84549), .ZN(n84544) );
  AOI22_X1 U70145 ( .A1(n105842), .A2(n110066), .B1(n105841), .B2(n110067), 
        .ZN(n84549) );
  NAND2_X1 U70146 ( .A1(n84550), .A2(n84551), .ZN(n84543) );
  AOI22_X1 U70147 ( .A1(n105840), .A2(n110088), .B1(n73222), .B2(n105839), 
        .ZN(n84551) );
  AOI22_X1 U70148 ( .A1(n105838), .A2(n110079), .B1(n105837), .B2(n110081), 
        .ZN(n84550) );
  NOR4_X1 U70149 ( .A1(n84552), .A2(n84553), .A3(n84554), .A4(n84555), .ZN(
        n84541) );
  OAI21_X1 U70150 ( .B1(n103138), .B2(n84146), .A(n84556), .ZN(n84555) );
  AOI22_X1 U70151 ( .A1(n105835), .A2(n110019), .B1(n105834), .B2(n110022), 
        .ZN(n84556) );
  OAI21_X1 U70152 ( .B1(n101033), .B2(n105833), .A(n84557), .ZN(n84554) );
  AOI22_X1 U70153 ( .A1(n73146), .A2(n105832), .B1(n105831), .B2(n110016), 
        .ZN(n84557) );
  OAI21_X1 U70154 ( .B1(n105830), .B2(n104603), .A(n84558), .ZN(n84553) );
  AOI22_X1 U70155 ( .A1(n73154), .A2(n105829), .B1(n73158), .B2(n105828), .ZN(
        n84558) );
  OAI21_X1 U70156 ( .B1(n101149), .B2(n105827), .A(n84559), .ZN(n84552) );
  AOI22_X1 U70157 ( .A1(n105826), .A2(n110044), .B1(n105825), .B2(n110041), 
        .ZN(n84559) );
  AOI22_X1 U70158 ( .A1(n84162), .A2(n110115), .B1(n84163), .B2(n110112), .ZN(
        n84538) );
  NOR4_X1 U70159 ( .A1(n84561), .A2(n84562), .A3(n84563), .A4(n84564), .ZN(
        n84560) );
  NAND2_X1 U70160 ( .A1(n84565), .A2(n84566), .ZN(n84564) );
  AOI22_X1 U70161 ( .A1(n105172), .A2(n110186), .B1(n73324), .B2(n106288), 
        .ZN(n84566) );
  AOI22_X1 U70162 ( .A1(n106284), .A2(n110148), .B1(n106276), .B2(n110126), 
        .ZN(n84565) );
  NAND2_X1 U70163 ( .A1(n84567), .A2(n84568), .ZN(n84563) );
  AOI22_X1 U70164 ( .A1(n105853), .A2(n110203), .B1(n105852), .B2(n110215), 
        .ZN(n84568) );
  AOI22_X1 U70165 ( .A1(n73292), .A2(n105100), .B1(n106746), .B2(n110173), 
        .ZN(n84567) );
  NAND2_X1 U70166 ( .A1(n84569), .A2(n84570), .ZN(n84562) );
  AOI22_X1 U70167 ( .A1(n105851), .A2(n110207), .B1(n84111), .B2(n110199), 
        .ZN(n84570) );
  AOI22_X1 U70168 ( .A1(n84112), .A2(n110211), .B1(n84113), .B2(n110121), .ZN(
        n84569) );
  NAND2_X1 U70169 ( .A1(n84571), .A2(n84572), .ZN(n84561) );
  AOI21_X1 U70170 ( .B1(n73381), .B2(n84116), .A(n84573), .ZN(n84572) );
  AOI21_X1 U70171 ( .B1(n84574), .B2(n84575), .A(n106325), .ZN(n84573) );
  NOR4_X1 U70172 ( .A1(n84576), .A2(n84577), .A3(n84578), .A4(n84579), .ZN(
        n84575) );
  OAI21_X1 U70173 ( .B1(n103111), .B2(n105849), .A(n84580), .ZN(n84579) );
  AOI22_X1 U70174 ( .A1(n73324), .A2(n84126), .B1(n105847), .B2(n110158), .ZN(
        n84580) );
  OAI21_X1 U70175 ( .B1(n103113), .B2(n84128), .A(n84581), .ZN(n84578) );
  AOI22_X1 U70176 ( .A1(n105845), .A2(n110182), .B1(n73336), .B2(n105844), 
        .ZN(n84581) );
  OAI21_X1 U70177 ( .B1(n103109), .B2(n105843), .A(n84582), .ZN(n84577) );
  AOI22_X1 U70178 ( .A1(n105842), .A2(n110173), .B1(n105841), .B2(n110174), 
        .ZN(n84582) );
  NAND2_X1 U70179 ( .A1(n84583), .A2(n84584), .ZN(n84576) );
  AOI22_X1 U70180 ( .A1(n105840), .A2(n110195), .B1(n73364), .B2(n105839), 
        .ZN(n84584) );
  AOI22_X1 U70181 ( .A1(n105838), .A2(n110186), .B1(n105837), .B2(n110188), 
        .ZN(n84583) );
  NOR4_X1 U70182 ( .A1(n84585), .A2(n84586), .A3(n84587), .A4(n84588), .ZN(
        n84574) );
  OAI21_X1 U70183 ( .B1(n103120), .B2(n84146), .A(n84589), .ZN(n84588) );
  AOI22_X1 U70184 ( .A1(n105835), .A2(n110126), .B1(n105834), .B2(n110129), 
        .ZN(n84589) );
  OAI21_X1 U70185 ( .B1(n101034), .B2(n84150), .A(n84590), .ZN(n84587) );
  AOI22_X1 U70186 ( .A1(n73288), .A2(n105832), .B1(n105831), .B2(n110123), 
        .ZN(n84590) );
  OAI21_X1 U70187 ( .B1(n84154), .B2(n104602), .A(n84591), .ZN(n84586) );
  AOI22_X1 U70188 ( .A1(n73296), .A2(n105829), .B1(n73300), .B2(n105828), .ZN(
        n84591) );
  OAI21_X1 U70189 ( .B1(n103116), .B2(n84158), .A(n84592), .ZN(n84585) );
  AOI22_X1 U70190 ( .A1(n105826), .A2(n110151), .B1(n105825), .B2(n110148), 
        .ZN(n84592) );
  AOI22_X1 U70191 ( .A1(n84162), .A2(n110222), .B1(n84163), .B2(n110219), .ZN(
        n84571) );
  NOR4_X1 U70192 ( .A1(n84594), .A2(n84595), .A3(n84596), .A4(n84597), .ZN(
        n84593) );
  NAND2_X1 U70193 ( .A1(n84598), .A2(n84599), .ZN(n84597) );
  AOI22_X1 U70194 ( .A1(n106745), .A2(n109971), .B1(n73040), .B2(n106288), 
        .ZN(n84599) );
  AOI22_X1 U70195 ( .A1(n106283), .A2(n109932), .B1(n106276), .B2(n109910), 
        .ZN(n84598) );
  NAND2_X1 U70196 ( .A1(n84600), .A2(n84601), .ZN(n84596) );
  AOI22_X1 U70197 ( .A1(n105853), .A2(n109988), .B1(n105852), .B2(n110000), 
        .ZN(n84601) );
  AOI22_X1 U70198 ( .A1(n73008), .A2(n81199), .B1(n105173), .B2(n109957), .ZN(
        n84600) );
  NAND2_X1 U70199 ( .A1(n84602), .A2(n84603), .ZN(n84595) );
  AOI22_X1 U70200 ( .A1(n105851), .A2(n109992), .B1(n84111), .B2(n109984), 
        .ZN(n84603) );
  AOI22_X1 U70201 ( .A1(n84112), .A2(n109996), .B1(n84113), .B2(n109904), .ZN(
        n84602) );
  NAND2_X1 U70202 ( .A1(n84604), .A2(n84605), .ZN(n84594) );
  AOI21_X1 U70203 ( .B1(n73097), .B2(n84116), .A(n84606), .ZN(n84605) );
  AOI21_X1 U70204 ( .B1(n84607), .B2(n84608), .A(n106324), .ZN(n84606) );
  NOR4_X1 U70205 ( .A1(n84609), .A2(n84610), .A3(n84611), .A4(n84612), .ZN(
        n84608) );
  OAI21_X1 U70206 ( .B1(n103091), .B2(n84124), .A(n84613), .ZN(n84612) );
  AOI22_X1 U70207 ( .A1(n73040), .A2(n84126), .B1(n105847), .B2(n109942), .ZN(
        n84613) );
  OAI21_X1 U70208 ( .B1(n103093), .B2(n105846), .A(n84614), .ZN(n84611) );
  AOI22_X1 U70209 ( .A1(n105845), .A2(n109967), .B1(n73052), .B2(n105844), 
        .ZN(n84614) );
  OAI21_X1 U70210 ( .B1(n103089), .B2(n84132), .A(n84615), .ZN(n84610) );
  AOI22_X1 U70211 ( .A1(n105842), .A2(n109957), .B1(n105841), .B2(n109959), 
        .ZN(n84615) );
  NAND2_X1 U70212 ( .A1(n84616), .A2(n84617), .ZN(n84609) );
  AOI22_X1 U70213 ( .A1(n105840), .A2(n109980), .B1(n73080), .B2(n105839), 
        .ZN(n84617) );
  AOI22_X1 U70214 ( .A1(n105838), .A2(n109971), .B1(n105837), .B2(n109973), 
        .ZN(n84616) );
  NOR4_X1 U70215 ( .A1(n84618), .A2(n84619), .A3(n84620), .A4(n84621), .ZN(
        n84607) );
  OAI21_X1 U70216 ( .B1(n103100), .B2(n105836), .A(n84622), .ZN(n84621) );
  AOI22_X1 U70217 ( .A1(n105835), .A2(n109910), .B1(n105834), .B2(n109913), 
        .ZN(n84622) );
  OAI21_X1 U70218 ( .B1(n101035), .B2(n105833), .A(n84623), .ZN(n84620) );
  AOI22_X1 U70219 ( .A1(n73004), .A2(n105832), .B1(n105831), .B2(n109907), 
        .ZN(n84623) );
  OAI21_X1 U70220 ( .B1(n105830), .B2(n104601), .A(n84624), .ZN(n84619) );
  AOI22_X1 U70221 ( .A1(n73012), .A2(n105829), .B1(n73016), .B2(n105828), .ZN(
        n84624) );
  OAI21_X1 U70222 ( .B1(n103096), .B2(n105827), .A(n84625), .ZN(n84618) );
  AOI22_X1 U70223 ( .A1(n105826), .A2(n109935), .B1(n105825), .B2(n109932), 
        .ZN(n84625) );
  AOI22_X1 U70224 ( .A1(n84162), .A2(n110007), .B1(n84163), .B2(n110004), .ZN(
        n84604) );
  NOR4_X1 U70225 ( .A1(n84627), .A2(n84628), .A3(n84629), .A4(n84630), .ZN(
        n84626) );
  NAND2_X1 U70226 ( .A1(n84631), .A2(n84632), .ZN(n84630) );
  AOI22_X1 U70227 ( .A1(n105172), .A2(n109854), .B1(n72890), .B2(n106288), 
        .ZN(n84632) );
  AOI22_X1 U70228 ( .A1(n106284), .A2(n109815), .B1(n106276), .B2(n109792), 
        .ZN(n84631) );
  NAND2_X1 U70229 ( .A1(n84633), .A2(n84634), .ZN(n84629) );
  AOI22_X1 U70230 ( .A1(n105853), .A2(n109871), .B1(n105852), .B2(n109883), 
        .ZN(n84634) );
  AOI22_X1 U70231 ( .A1(n72858), .A2(n105100), .B1(n106746), .B2(n109840), 
        .ZN(n84633) );
  NAND2_X1 U70232 ( .A1(n84635), .A2(n84636), .ZN(n84628) );
  AOI22_X1 U70233 ( .A1(n105851), .A2(n109875), .B1(n84111), .B2(n109867), 
        .ZN(n84636) );
  AOI22_X1 U70234 ( .A1(n84112), .A2(n109879), .B1(n105850), .B2(n109786), 
        .ZN(n84635) );
  NAND2_X1 U70235 ( .A1(n84637), .A2(n84638), .ZN(n84627) );
  AOI21_X1 U70236 ( .B1(n72947), .B2(n84116), .A(n84639), .ZN(n84638) );
  AOI21_X1 U70237 ( .B1(n84640), .B2(n84641), .A(n106325), .ZN(n84639) );
  NOR4_X1 U70238 ( .A1(n84642), .A2(n84643), .A3(n84644), .A4(n84645), .ZN(
        n84641) );
  OAI21_X1 U70239 ( .B1(n103071), .B2(n105849), .A(n84646), .ZN(n84645) );
  AOI22_X1 U70240 ( .A1(n72890), .A2(n105848), .B1(n105847), .B2(n109825), 
        .ZN(n84646) );
  OAI21_X1 U70241 ( .B1(n103073), .B2(n84128), .A(n84647), .ZN(n84644) );
  AOI22_X1 U70242 ( .A1(n105845), .A2(n109850), .B1(n72902), .B2(n105844), 
        .ZN(n84647) );
  OAI21_X1 U70243 ( .B1(n103069), .B2(n105843), .A(n84648), .ZN(n84643) );
  AOI22_X1 U70244 ( .A1(n105842), .A2(n109840), .B1(n105841), .B2(n109842), 
        .ZN(n84648) );
  NAND2_X1 U70245 ( .A1(n84649), .A2(n84650), .ZN(n84642) );
  AOI22_X1 U70246 ( .A1(n105840), .A2(n109863), .B1(n72930), .B2(n105839), 
        .ZN(n84650) );
  AOI22_X1 U70247 ( .A1(n105838), .A2(n109854), .B1(n105837), .B2(n109856), 
        .ZN(n84649) );
  NOR4_X1 U70248 ( .A1(n84651), .A2(n84652), .A3(n84653), .A4(n84654), .ZN(
        n84640) );
  OAI21_X1 U70249 ( .B1(n103080), .B2(n84146), .A(n84655), .ZN(n84654) );
  AOI22_X1 U70250 ( .A1(n105835), .A2(n109792), .B1(n105834), .B2(n109795), 
        .ZN(n84655) );
  OAI21_X1 U70251 ( .B1(n101036), .B2(n84150), .A(n84656), .ZN(n84653) );
  AOI22_X1 U70252 ( .A1(n72854), .A2(n105832), .B1(n105831), .B2(n109789), 
        .ZN(n84656) );
  OAI21_X1 U70253 ( .B1(n84154), .B2(n104600), .A(n84657), .ZN(n84652) );
  AOI22_X1 U70254 ( .A1(n72862), .A2(n105829), .B1(n72866), .B2(n105828), .ZN(
        n84657) );
  OAI21_X1 U70255 ( .B1(n103076), .B2(n84158), .A(n84658), .ZN(n84651) );
  AOI22_X1 U70256 ( .A1(n105826), .A2(n109818), .B1(n105825), .B2(n109815), 
        .ZN(n84658) );
  AOI22_X1 U70257 ( .A1(n84162), .A2(n109890), .B1(n84163), .B2(n109887), .ZN(
        n84637) );
  NOR4_X1 U70258 ( .A1(n84660), .A2(n84661), .A3(n84662), .A4(n84663), .ZN(
        n84659) );
  NAND2_X1 U70259 ( .A1(n84664), .A2(n84665), .ZN(n84663) );
  AOI22_X1 U70260 ( .A1(n105170), .A2(n108228), .B1(n70786), .B2(n106288), 
        .ZN(n84665) );
  AOI22_X1 U70261 ( .A1(n106283), .A2(n108189), .B1(n106276), .B2(n108166), 
        .ZN(n84664) );
  NAND2_X1 U70262 ( .A1(n84666), .A2(n84667), .ZN(n84662) );
  AOI22_X1 U70263 ( .A1(n105853), .A2(n108245), .B1(n105852), .B2(n108257), 
        .ZN(n84667) );
  AOI22_X1 U70264 ( .A1(n70754), .A2(n105101), .B1(n106746), .B2(n108214), 
        .ZN(n84666) );
  NAND2_X1 U70265 ( .A1(n84668), .A2(n84669), .ZN(n84661) );
  AOI22_X1 U70266 ( .A1(n105851), .A2(n108249), .B1(n84111), .B2(n108241), 
        .ZN(n84669) );
  AOI22_X1 U70267 ( .A1(n84112), .A2(n108253), .B1(n84113), .B2(n108160), .ZN(
        n84668) );
  NAND2_X1 U70268 ( .A1(n84670), .A2(n84671), .ZN(n84660) );
  AOI21_X1 U70269 ( .B1(n70843), .B2(n84116), .A(n84672), .ZN(n84671) );
  AOI21_X1 U70270 ( .B1(n84673), .B2(n84674), .A(n106326), .ZN(n84672) );
  NOR4_X1 U70271 ( .A1(n84675), .A2(n84676), .A3(n84677), .A4(n84678), .ZN(
        n84674) );
  OAI21_X1 U70272 ( .B1(n103051), .B2(n105849), .A(n84679), .ZN(n84678) );
  AOI22_X1 U70273 ( .A1(n70786), .A2(n84126), .B1(n84127), .B2(n108199), .ZN(
        n84679) );
  OAI21_X1 U70274 ( .B1(n103053), .B2(n105846), .A(n84680), .ZN(n84677) );
  AOI22_X1 U70275 ( .A1(n105845), .A2(n108224), .B1(n70798), .B2(n105844), 
        .ZN(n84680) );
  OAI21_X1 U70276 ( .B1(n103049), .B2(n84132), .A(n84681), .ZN(n84676) );
  AOI22_X1 U70277 ( .A1(n105842), .A2(n108214), .B1(n105841), .B2(n108216), 
        .ZN(n84681) );
  NAND2_X1 U70278 ( .A1(n84682), .A2(n84683), .ZN(n84675) );
  AOI22_X1 U70279 ( .A1(n105840), .A2(n108237), .B1(n70826), .B2(n105839), 
        .ZN(n84683) );
  AOI22_X1 U70280 ( .A1(n105838), .A2(n108228), .B1(n105837), .B2(n108230), 
        .ZN(n84682) );
  NOR4_X1 U70281 ( .A1(n84684), .A2(n84685), .A3(n84686), .A4(n84687), .ZN(
        n84673) );
  OAI21_X1 U70282 ( .B1(n103060), .B2(n105836), .A(n84688), .ZN(n84687) );
  AOI22_X1 U70283 ( .A1(n105835), .A2(n108166), .B1(n105834), .B2(n108169), 
        .ZN(n84688) );
  OAI21_X1 U70284 ( .B1(n101037), .B2(n105833), .A(n84689), .ZN(n84686) );
  AOI22_X1 U70285 ( .A1(n70750), .A2(n105832), .B1(n105831), .B2(n108163), 
        .ZN(n84689) );
  OAI21_X1 U70286 ( .B1(n105830), .B2(n104599), .A(n84690), .ZN(n84685) );
  AOI22_X1 U70287 ( .A1(n70758), .A2(n105829), .B1(n70762), .B2(n105828), .ZN(
        n84690) );
  OAI21_X1 U70288 ( .B1(n103056), .B2(n84158), .A(n84691), .ZN(n84684) );
  AOI22_X1 U70289 ( .A1(n105826), .A2(n108192), .B1(n105825), .B2(n108189), 
        .ZN(n84691) );
  AOI22_X1 U70290 ( .A1(n84162), .A2(n108264), .B1(n84163), .B2(n108261), .ZN(
        n84670) );
  NOR4_X1 U70291 ( .A1(n84693), .A2(n84694), .A3(n84695), .A4(n84696), .ZN(
        n84692) );
  NAND2_X1 U70292 ( .A1(n84697), .A2(n84698), .ZN(n84696) );
  AOI22_X1 U70293 ( .A1(n105171), .A2(n108351), .B1(n70945), .B2(n106288), 
        .ZN(n84698) );
  AOI22_X1 U70294 ( .A1(n106283), .A2(n108312), .B1(n106276), .B2(n108289), 
        .ZN(n84697) );
  NAND2_X1 U70295 ( .A1(n84699), .A2(n84700), .ZN(n84695) );
  AOI22_X1 U70296 ( .A1(n105853), .A2(n108368), .B1(n105852), .B2(n108380), 
        .ZN(n84700) );
  AOI22_X1 U70297 ( .A1(n70913), .A2(n105100), .B1(n105174), .B2(n108337), 
        .ZN(n84699) );
  NAND2_X1 U70298 ( .A1(n84701), .A2(n84702), .ZN(n84694) );
  AOI22_X1 U70299 ( .A1(n105851), .A2(n108372), .B1(n84111), .B2(n108364), 
        .ZN(n84702) );
  AOI22_X1 U70300 ( .A1(n84112), .A2(n108376), .B1(n105850), .B2(n108283), 
        .ZN(n84701) );
  NAND2_X1 U70301 ( .A1(n84703), .A2(n84704), .ZN(n84693) );
  AOI21_X1 U70302 ( .B1(n71002), .B2(n84116), .A(n84705), .ZN(n84704) );
  AOI21_X1 U70303 ( .B1(n84706), .B2(n84707), .A(n106323), .ZN(n84705) );
  NOR4_X1 U70304 ( .A1(n84708), .A2(n84709), .A3(n84710), .A4(n84711), .ZN(
        n84707) );
  OAI21_X1 U70305 ( .B1(n103031), .B2(n84124), .A(n84712), .ZN(n84711) );
  AOI22_X1 U70306 ( .A1(n70945), .A2(n105848), .B1(n105847), .B2(n108322), 
        .ZN(n84712) );
  OAI21_X1 U70307 ( .B1(n103033), .B2(n84128), .A(n84713), .ZN(n84710) );
  AOI22_X1 U70308 ( .A1(n105845), .A2(n108347), .B1(n70957), .B2(n105844), 
        .ZN(n84713) );
  OAI21_X1 U70309 ( .B1(n103029), .B2(n105843), .A(n84714), .ZN(n84709) );
  AOI22_X1 U70310 ( .A1(n105842), .A2(n108337), .B1(n105841), .B2(n108339), 
        .ZN(n84714) );
  NAND2_X1 U70311 ( .A1(n84715), .A2(n84716), .ZN(n84708) );
  AOI22_X1 U70312 ( .A1(n105840), .A2(n108360), .B1(n70985), .B2(n105839), 
        .ZN(n84716) );
  AOI22_X1 U70313 ( .A1(n105838), .A2(n108351), .B1(n105837), .B2(n108353), 
        .ZN(n84715) );
  NOR4_X1 U70314 ( .A1(n84717), .A2(n84718), .A3(n84719), .A4(n84720), .ZN(
        n84706) );
  OAI21_X1 U70315 ( .B1(n103040), .B2(n84146), .A(n84721), .ZN(n84720) );
  AOI22_X1 U70316 ( .A1(n105835), .A2(n108289), .B1(n105834), .B2(n108292), 
        .ZN(n84721) );
  OAI21_X1 U70317 ( .B1(n101038), .B2(n84150), .A(n84722), .ZN(n84719) );
  AOI22_X1 U70318 ( .A1(n70909), .A2(n105832), .B1(n105831), .B2(n108286), 
        .ZN(n84722) );
  OAI21_X1 U70319 ( .B1(n84154), .B2(n104598), .A(n84723), .ZN(n84718) );
  AOI22_X1 U70320 ( .A1(n70917), .A2(n105829), .B1(n70921), .B2(n105828), .ZN(
        n84723) );
  OAI21_X1 U70321 ( .B1(n103036), .B2(n84158), .A(n84724), .ZN(n84717) );
  AOI22_X1 U70322 ( .A1(n105826), .A2(n108315), .B1(n105825), .B2(n108312), 
        .ZN(n84724) );
  AOI22_X1 U70323 ( .A1(n84162), .A2(n108387), .B1(n84163), .B2(n108384), .ZN(
        n84703) );
  NOR4_X1 U70324 ( .A1(n84726), .A2(n84727), .A3(n84728), .A4(n84729), .ZN(
        n84725) );
  NAND2_X1 U70325 ( .A1(n84730), .A2(n84731), .ZN(n84729) );
  AOI22_X1 U70326 ( .A1(n105172), .A2(n108462), .B1(n71090), .B2(n106288), 
        .ZN(n84731) );
  AOI22_X1 U70327 ( .A1(n106283), .A2(n108423), .B1(n106276), .B2(n108400), 
        .ZN(n84730) );
  NAND2_X1 U70328 ( .A1(n84732), .A2(n84733), .ZN(n84728) );
  AOI22_X1 U70329 ( .A1(n105853), .A2(n108479), .B1(n105852), .B2(n108491), 
        .ZN(n84733) );
  AOI22_X1 U70330 ( .A1(n71058), .A2(n105100), .B1(n106746), .B2(n108448), 
        .ZN(n84732) );
  NAND2_X1 U70331 ( .A1(n84734), .A2(n84735), .ZN(n84727) );
  AOI22_X1 U70332 ( .A1(n105851), .A2(n108483), .B1(n84111), .B2(n108475), 
        .ZN(n84735) );
  AOI22_X1 U70333 ( .A1(n84112), .A2(n108487), .B1(n84113), .B2(n108394), .ZN(
        n84734) );
  NAND2_X1 U70334 ( .A1(n84736), .A2(n84737), .ZN(n84726) );
  AOI21_X1 U70335 ( .B1(n71147), .B2(n84116), .A(n84738), .ZN(n84737) );
  AOI21_X1 U70336 ( .B1(n84739), .B2(n84740), .A(n106327), .ZN(n84738) );
  NOR4_X1 U70337 ( .A1(n84741), .A2(n84742), .A3(n84743), .A4(n84744), .ZN(
        n84740) );
  OAI21_X1 U70338 ( .B1(n103011), .B2(n105849), .A(n84745), .ZN(n84744) );
  AOI22_X1 U70339 ( .A1(n71090), .A2(n84126), .B1(n84127), .B2(n108433), .ZN(
        n84745) );
  OAI21_X1 U70340 ( .B1(n103013), .B2(n105846), .A(n84746), .ZN(n84743) );
  AOI22_X1 U70341 ( .A1(n105845), .A2(n108458), .B1(n71102), .B2(n105844), 
        .ZN(n84746) );
  OAI21_X1 U70342 ( .B1(n103009), .B2(n84132), .A(n84747), .ZN(n84742) );
  AOI22_X1 U70343 ( .A1(n105842), .A2(n108448), .B1(n84135), .B2(n108450), 
        .ZN(n84747) );
  NAND2_X1 U70344 ( .A1(n84748), .A2(n84749), .ZN(n84741) );
  AOI22_X1 U70345 ( .A1(n105840), .A2(n108471), .B1(n71130), .B2(n105839), 
        .ZN(n84749) );
  AOI22_X1 U70346 ( .A1(n105838), .A2(n108462), .B1(n105837), .B2(n108464), 
        .ZN(n84748) );
  NOR4_X1 U70347 ( .A1(n84750), .A2(n84751), .A3(n84752), .A4(n84753), .ZN(
        n84739) );
  OAI21_X1 U70348 ( .B1(n103020), .B2(n105836), .A(n84754), .ZN(n84753) );
  AOI22_X1 U70349 ( .A1(n105835), .A2(n108400), .B1(n105834), .B2(n108403), 
        .ZN(n84754) );
  OAI21_X1 U70350 ( .B1(n101039), .B2(n105833), .A(n84755), .ZN(n84752) );
  AOI22_X1 U70351 ( .A1(n71054), .A2(n105832), .B1(n105831), .B2(n108397), 
        .ZN(n84755) );
  OAI21_X1 U70352 ( .B1(n105830), .B2(n104597), .A(n84756), .ZN(n84751) );
  AOI22_X1 U70353 ( .A1(n71062), .A2(n105829), .B1(n71066), .B2(n105828), .ZN(
        n84756) );
  OAI21_X1 U70354 ( .B1(n103016), .B2(n84158), .A(n84757), .ZN(n84750) );
  AOI22_X1 U70355 ( .A1(n105826), .A2(n108426), .B1(n105825), .B2(n108423), 
        .ZN(n84757) );
  AOI22_X1 U70356 ( .A1(n84162), .A2(n108498), .B1(n84163), .B2(n108495), .ZN(
        n84736) );
  NOR4_X1 U70357 ( .A1(n84759), .A2(n84760), .A3(n84761), .A4(n84762), .ZN(
        n84758) );
  NAND2_X1 U70358 ( .A1(n84763), .A2(n84764), .ZN(n84762) );
  AOI22_X1 U70359 ( .A1(n106745), .A2(n107700), .B1(n70051), .B2(n106288), 
        .ZN(n84764) );
  AOI22_X1 U70360 ( .A1(n106282), .A2(n107661), .B1(n106276), .B2(n107638), 
        .ZN(n84763) );
  NAND2_X1 U70361 ( .A1(n84765), .A2(n84766), .ZN(n84761) );
  AOI22_X1 U70362 ( .A1(n105853), .A2(n107716), .B1(n105852), .B2(n107728), 
        .ZN(n84766) );
  AOI22_X1 U70363 ( .A1(n70019), .A2(n105100), .B1(n106746), .B2(n107686), 
        .ZN(n84765) );
  NAND2_X1 U70364 ( .A1(n84767), .A2(n84768), .ZN(n84760) );
  AOI22_X1 U70365 ( .A1(n105851), .A2(n107720), .B1(n84111), .B2(n107712), 
        .ZN(n84768) );
  AOI22_X1 U70366 ( .A1(n84112), .A2(n107724), .B1(n105850), .B2(n107632), 
        .ZN(n84767) );
  NAND2_X1 U70367 ( .A1(n84769), .A2(n84770), .ZN(n84759) );
  AOI21_X1 U70368 ( .B1(n70108), .B2(n84116), .A(n84771), .ZN(n84770) );
  AOI21_X1 U70369 ( .B1(n84772), .B2(n84773), .A(n106323), .ZN(n84771) );
  NOR4_X1 U70370 ( .A1(n84774), .A2(n84775), .A3(n84776), .A4(n84777), .ZN(
        n84773) );
  OAI21_X1 U70371 ( .B1(n102991), .B2(n84124), .A(n84778), .ZN(n84777) );
  AOI22_X1 U70372 ( .A1(n70051), .A2(n105848), .B1(n84127), .B2(n107671), .ZN(
        n84778) );
  OAI21_X1 U70373 ( .B1(n102993), .B2(n84128), .A(n84779), .ZN(n84776) );
  AOI22_X1 U70374 ( .A1(n105845), .A2(n107696), .B1(n70063), .B2(n105844), 
        .ZN(n84779) );
  OAI21_X1 U70375 ( .B1(n102989), .B2(n105843), .A(n84780), .ZN(n84775) );
  AOI22_X1 U70376 ( .A1(n105842), .A2(n107686), .B1(n84135), .B2(n107688), 
        .ZN(n84780) );
  NAND2_X1 U70377 ( .A1(n84781), .A2(n84782), .ZN(n84774) );
  AOI22_X1 U70378 ( .A1(n105840), .A2(n107709), .B1(n70091), .B2(n105839), 
        .ZN(n84782) );
  AOI22_X1 U70379 ( .A1(n105838), .A2(n107700), .B1(n105837), .B2(n107702), 
        .ZN(n84781) );
  NOR4_X1 U70380 ( .A1(n84783), .A2(n84784), .A3(n84785), .A4(n84786), .ZN(
        n84772) );
  OAI21_X1 U70381 ( .B1(n103000), .B2(n84146), .A(n84787), .ZN(n84786) );
  AOI22_X1 U70382 ( .A1(n105835), .A2(n107638), .B1(n105834), .B2(n107641), 
        .ZN(n84787) );
  OAI21_X1 U70383 ( .B1(n101040), .B2(n84150), .A(n84788), .ZN(n84785) );
  AOI22_X1 U70384 ( .A1(n70015), .A2(n105832), .B1(n105831), .B2(n107635), 
        .ZN(n84788) );
  OAI21_X1 U70385 ( .B1(n84154), .B2(n104596), .A(n84789), .ZN(n84784) );
  AOI22_X1 U70386 ( .A1(n70023), .A2(n105829), .B1(n70027), .B2(n105828), .ZN(
        n84789) );
  OAI21_X1 U70387 ( .B1(n102996), .B2(n84158), .A(n84790), .ZN(n84783) );
  AOI22_X1 U70388 ( .A1(n105826), .A2(n107664), .B1(n84161), .B2(n107661), 
        .ZN(n84790) );
  AOI22_X1 U70389 ( .A1(n84162), .A2(n107735), .B1(n84163), .B2(n107732), .ZN(
        n84769) );
  NOR4_X1 U70390 ( .A1(n84792), .A2(n84793), .A3(n84794), .A4(n84795), .ZN(
        n84791) );
  NAND2_X1 U70391 ( .A1(n84796), .A2(n84797), .ZN(n84795) );
  AOI22_X1 U70392 ( .A1(n105170), .A2(n109615), .B1(n72580), .B2(n106288), 
        .ZN(n84797) );
  AOI22_X1 U70393 ( .A1(n106283), .A2(n109579), .B1(n106276), .B2(n109556), 
        .ZN(n84796) );
  NAND2_X1 U70394 ( .A1(n84798), .A2(n84799), .ZN(n84794) );
  AOI22_X1 U70395 ( .A1(n84106), .A2(n109631), .B1(n105852), .B2(n109643), 
        .ZN(n84799) );
  AOI22_X1 U70396 ( .A1(n72548), .A2(n105099), .B1(n105173), .B2(n109604), 
        .ZN(n84798) );
  NAND2_X1 U70397 ( .A1(n84800), .A2(n84801), .ZN(n84793) );
  AOI22_X1 U70398 ( .A1(n105851), .A2(n109635), .B1(n84111), .B2(n109627), 
        .ZN(n84801) );
  AOI22_X1 U70399 ( .A1(n84112), .A2(n109639), .B1(n84113), .B2(n109550), .ZN(
        n84800) );
  NAND2_X1 U70400 ( .A1(n84802), .A2(n84803), .ZN(n84792) );
  AOI21_X1 U70401 ( .B1(n72637), .B2(n84116), .A(n84804), .ZN(n84803) );
  AOI21_X1 U70402 ( .B1(n84805), .B2(n84806), .A(n106323), .ZN(n84804) );
  NOR4_X1 U70403 ( .A1(n84807), .A2(n84808), .A3(n84809), .A4(n84810), .ZN(
        n84806) );
  OAI21_X1 U70404 ( .B1(n102973), .B2(n84124), .A(n84811), .ZN(n84810) );
  AOI22_X1 U70405 ( .A1(n72580), .A2(n84126), .B1(n84127), .B2(n109589), .ZN(
        n84811) );
  OAI21_X1 U70406 ( .B1(n102975), .B2(n105846), .A(n84812), .ZN(n84809) );
  AOI22_X1 U70407 ( .A1(n105845), .A2(n109611), .B1(n72592), .B2(n84131), .ZN(
        n84812) );
  OAI21_X1 U70408 ( .B1(n102971), .B2(n84132), .A(n84813), .ZN(n84808) );
  AOI22_X1 U70409 ( .A1(n105842), .A2(n109604), .B1(n72600), .B2(n105841), 
        .ZN(n84813) );
  NAND2_X1 U70410 ( .A1(n84814), .A2(n84815), .ZN(n84807) );
  AOI22_X1 U70411 ( .A1(n105840), .A2(n109624), .B1(n72620), .B2(n105839), 
        .ZN(n84815) );
  AOI22_X1 U70412 ( .A1(n105838), .A2(n109615), .B1(n105837), .B2(n109617), 
        .ZN(n84814) );
  NOR4_X1 U70413 ( .A1(n84816), .A2(n84817), .A3(n84818), .A4(n84819), .ZN(
        n84805) );
  OAI21_X1 U70414 ( .B1(n102980), .B2(n105836), .A(n84820), .ZN(n84819) );
  AOI22_X1 U70415 ( .A1(n105835), .A2(n109556), .B1(n84149), .B2(n109559), 
        .ZN(n84820) );
  OAI21_X1 U70416 ( .B1(n101041), .B2(n105833), .A(n84821), .ZN(n84818) );
  AOI22_X1 U70417 ( .A1(n72544), .A2(n105832), .B1(n105831), .B2(n109553), 
        .ZN(n84821) );
  OAI21_X1 U70418 ( .B1(n105830), .B2(n104595), .A(n84822), .ZN(n84817) );
  AOI22_X1 U70419 ( .A1(n72552), .A2(n105829), .B1(n72556), .B2(n105828), .ZN(
        n84822) );
  OAI21_X1 U70420 ( .B1(n101150), .B2(n84158), .A(n84823), .ZN(n84816) );
  AOI22_X1 U70421 ( .A1(n84160), .A2(n109582), .B1(n84161), .B2(n109579), .ZN(
        n84823) );
  AOI22_X1 U70422 ( .A1(n84162), .A2(n109650), .B1(n84163), .B2(n109647), .ZN(
        n84802) );
  NOR4_X1 U70423 ( .A1(n84825), .A2(n84826), .A3(n84827), .A4(n84828), .ZN(
        n84824) );
  NAND2_X1 U70424 ( .A1(n84829), .A2(n84830), .ZN(n84828) );
  AOI22_X1 U70425 ( .A1(n105171), .A2(n108577), .B1(n71239), .B2(n106288), 
        .ZN(n84830) );
  AOI22_X1 U70426 ( .A1(n106283), .A2(n108540), .B1(n106276), .B2(n108517), 
        .ZN(n84829) );
  NAND2_X1 U70427 ( .A1(n84831), .A2(n84832), .ZN(n84827) );
  AOI22_X1 U70428 ( .A1(n84106), .A2(n108593), .B1(n105852), .B2(n108605), 
        .ZN(n84832) );
  AOI22_X1 U70429 ( .A1(n71207), .A2(n105100), .B1(n105175), .B2(n108565), 
        .ZN(n84831) );
  NAND2_X1 U70430 ( .A1(n84833), .A2(n84834), .ZN(n84826) );
  AOI22_X1 U70431 ( .A1(n105851), .A2(n108597), .B1(n84111), .B2(n108589), 
        .ZN(n84834) );
  AOI22_X1 U70432 ( .A1(n84112), .A2(n108601), .B1(n84113), .B2(n108511), .ZN(
        n84833) );
  NAND2_X1 U70433 ( .A1(n84835), .A2(n84836), .ZN(n84825) );
  AOI21_X1 U70434 ( .B1(n71296), .B2(n84116), .A(n84837), .ZN(n84836) );
  AOI21_X1 U70435 ( .B1(n84838), .B2(n84839), .A(n106326), .ZN(n84837) );
  NOR4_X1 U70436 ( .A1(n84840), .A2(n84841), .A3(n84842), .A4(n84843), .ZN(
        n84839) );
  OAI21_X1 U70437 ( .B1(n102954), .B2(n84124), .A(n84844), .ZN(n84843) );
  AOI22_X1 U70438 ( .A1(n71239), .A2(n84126), .B1(n84127), .B2(n108550), .ZN(
        n84844) );
  OAI21_X1 U70439 ( .B1(n102956), .B2(n105846), .A(n84845), .ZN(n84842) );
  AOI22_X1 U70440 ( .A1(n84130), .A2(n108573), .B1(n71251), .B2(n84131), .ZN(
        n84845) );
  OAI21_X1 U70441 ( .B1(n102952), .B2(n84132), .A(n84846), .ZN(n84841) );
  AOI22_X1 U70442 ( .A1(n84134), .A2(n108565), .B1(n84135), .B2(n108567), .ZN(
        n84846) );
  NAND2_X1 U70443 ( .A1(n84847), .A2(n84848), .ZN(n84840) );
  AOI22_X1 U70444 ( .A1(n105840), .A2(n108586), .B1(n71279), .B2(n84139), .ZN(
        n84848) );
  AOI22_X1 U70445 ( .A1(n105838), .A2(n108577), .B1(n105837), .B2(n108579), 
        .ZN(n84847) );
  NOR4_X1 U70446 ( .A1(n84849), .A2(n84850), .A3(n84851), .A4(n84852), .ZN(
        n84838) );
  OAI21_X1 U70447 ( .B1(n102963), .B2(n84146), .A(n84853), .ZN(n84852) );
  AOI22_X1 U70448 ( .A1(n105835), .A2(n108517), .B1(n84149), .B2(n108520), 
        .ZN(n84853) );
  OAI21_X1 U70449 ( .B1(n101042), .B2(n105833), .A(n84854), .ZN(n84851) );
  AOI22_X1 U70450 ( .A1(n71203), .A2(n105832), .B1(n105831), .B2(n108514), 
        .ZN(n84854) );
  OAI21_X1 U70451 ( .B1(n105830), .B2(n104594), .A(n84855), .ZN(n84850) );
  AOI22_X1 U70452 ( .A1(n71211), .A2(n105829), .B1(n71215), .B2(n105828), .ZN(
        n84855) );
  OAI21_X1 U70453 ( .B1(n102959), .B2(n84158), .A(n84856), .ZN(n84849) );
  AOI22_X1 U70454 ( .A1(n84160), .A2(n108543), .B1(n84161), .B2(n108540), .ZN(
        n84856) );
  AOI22_X1 U70455 ( .A1(n84162), .A2(n108612), .B1(n84163), .B2(n108609), .ZN(
        n84835) );
  NOR4_X1 U70456 ( .A1(n84858), .A2(n84859), .A3(n84860), .A4(n84861), .ZN(
        n84857) );
  NAND2_X1 U70457 ( .A1(n84862), .A2(n84863), .ZN(n84861) );
  AOI22_X1 U70458 ( .A1(n105172), .A2(n109722), .B1(n72722), .B2(n106288), 
        .ZN(n84863) );
  AOI22_X1 U70459 ( .A1(n80260), .A2(n109684), .B1(n106276), .B2(n109661), 
        .ZN(n84862) );
  NAND2_X1 U70460 ( .A1(n84864), .A2(n84865), .ZN(n84860) );
  AOI22_X1 U70461 ( .A1(n84106), .A2(n109738), .B1(n105852), .B2(n109750), 
        .ZN(n84865) );
  AOI22_X1 U70462 ( .A1(n72690), .A2(n105101), .B1(n105173), .B2(n109709), 
        .ZN(n84864) );
  NAND2_X1 U70463 ( .A1(n84866), .A2(n84867), .ZN(n84859) );
  AOI22_X1 U70464 ( .A1(n105851), .A2(n109742), .B1(n84111), .B2(n109734), 
        .ZN(n84867) );
  AOI22_X1 U70465 ( .A1(n84112), .A2(n109746), .B1(n105850), .B2(n109655), 
        .ZN(n84866) );
  NAND2_X1 U70466 ( .A1(n84868), .A2(n84869), .ZN(n84858) );
  AOI21_X1 U70467 ( .B1(n72779), .B2(n84116), .A(n84870), .ZN(n84869) );
  AOI21_X1 U70468 ( .B1(n84871), .B2(n84872), .A(n106324), .ZN(n84870) );
  NOR4_X1 U70469 ( .A1(n84873), .A2(n84874), .A3(n84875), .A4(n84876), .ZN(
        n84872) );
  OAI21_X1 U70470 ( .B1(n102934), .B2(n84124), .A(n84877), .ZN(n84876) );
  AOI22_X1 U70471 ( .A1(n72722), .A2(n105848), .B1(n84127), .B2(n109694), .ZN(
        n84877) );
  OAI21_X1 U70472 ( .B1(n102936), .B2(n105846), .A(n84878), .ZN(n84875) );
  AOI22_X1 U70473 ( .A1(n84130), .A2(n109718), .B1(n72734), .B2(n84131), .ZN(
        n84878) );
  OAI21_X1 U70474 ( .B1(n102932), .B2(n84132), .A(n84879), .ZN(n84874) );
  AOI22_X1 U70475 ( .A1(n84134), .A2(n109709), .B1(n84135), .B2(n109711), .ZN(
        n84879) );
  NAND2_X1 U70476 ( .A1(n84880), .A2(n84881), .ZN(n84873) );
  AOI22_X1 U70477 ( .A1(n105840), .A2(n109731), .B1(n72762), .B2(n84139), .ZN(
        n84881) );
  AOI22_X1 U70478 ( .A1(n105838), .A2(n109722), .B1(n105837), .B2(n109724), 
        .ZN(n84880) );
  NOR4_X1 U70479 ( .A1(n84882), .A2(n84883), .A3(n84884), .A4(n84885), .ZN(
        n84871) );
  OAI21_X1 U70480 ( .B1(n102943), .B2(n105836), .A(n84886), .ZN(n84885) );
  AOI22_X1 U70481 ( .A1(n105835), .A2(n109661), .B1(n84149), .B2(n109664), 
        .ZN(n84886) );
  OAI21_X1 U70482 ( .B1(n101043), .B2(n105833), .A(n84887), .ZN(n84884) );
  AOI22_X1 U70483 ( .A1(n72686), .A2(n105832), .B1(n105831), .B2(n109658), 
        .ZN(n84887) );
  OAI21_X1 U70484 ( .B1(n105830), .B2(n104593), .A(n84888), .ZN(n84883) );
  AOI22_X1 U70485 ( .A1(n72694), .A2(n105829), .B1(n72698), .B2(n105828), .ZN(
        n84888) );
  OAI21_X1 U70486 ( .B1(n102939), .B2(n84158), .A(n84889), .ZN(n84882) );
  AOI22_X1 U70487 ( .A1(n84160), .A2(n109687), .B1(n84161), .B2(n109684), .ZN(
        n84889) );
  AOI22_X1 U70488 ( .A1(n84162), .A2(n109757), .B1(n84163), .B2(n109754), .ZN(
        n84868) );
  NOR4_X1 U70489 ( .A1(n84891), .A2(n84892), .A3(n84893), .A4(n84894), .ZN(
        n84890) );
  NAND2_X1 U70490 ( .A1(n84895), .A2(n84896), .ZN(n84894) );
  AOI22_X1 U70491 ( .A1(n106745), .A2(n109507), .B1(n72432), .B2(n106289), 
        .ZN(n84896) );
  AOI22_X1 U70492 ( .A1(n106283), .A2(n109468), .B1(n106276), .B2(n109445), 
        .ZN(n84895) );
  NAND2_X1 U70493 ( .A1(n84897), .A2(n84898), .ZN(n84893) );
  AOI22_X1 U70494 ( .A1(n84106), .A2(n109523), .B1(n105852), .B2(n109535), 
        .ZN(n84898) );
  AOI22_X1 U70495 ( .A1(n72400), .A2(n105100), .B1(n105173), .B2(n109493), 
        .ZN(n84897) );
  NAND2_X1 U70496 ( .A1(n84899), .A2(n84900), .ZN(n84892) );
  AOI22_X1 U70497 ( .A1(n105851), .A2(n109527), .B1(n84111), .B2(n109519), 
        .ZN(n84900) );
  AOI22_X1 U70498 ( .A1(n84112), .A2(n109531), .B1(n84113), .B2(n109439), .ZN(
        n84899) );
  NAND2_X1 U70499 ( .A1(n84901), .A2(n84902), .ZN(n84891) );
  AOI21_X1 U70500 ( .B1(n72489), .B2(n84116), .A(n84903), .ZN(n84902) );
  AOI21_X1 U70501 ( .B1(n84904), .B2(n84905), .A(n106325), .ZN(n84903) );
  NOR4_X1 U70502 ( .A1(n84906), .A2(n84907), .A3(n84908), .A4(n84909), .ZN(
        n84905) );
  OAI21_X1 U70503 ( .B1(n102914), .B2(n84124), .A(n84910), .ZN(n84909) );
  AOI22_X1 U70504 ( .A1(n72432), .A2(n105848), .B1(n84127), .B2(n109478), .ZN(
        n84910) );
  OAI21_X1 U70505 ( .B1(n102916), .B2(n105846), .A(n84911), .ZN(n84908) );
  AOI22_X1 U70506 ( .A1(n84130), .A2(n109503), .B1(n72444), .B2(n84131), .ZN(
        n84911) );
  OAI21_X1 U70507 ( .B1(n102912), .B2(n84132), .A(n84912), .ZN(n84907) );
  AOI22_X1 U70508 ( .A1(n84134), .A2(n109493), .B1(n84135), .B2(n109495), .ZN(
        n84912) );
  NAND2_X1 U70509 ( .A1(n84913), .A2(n84914), .ZN(n84906) );
  AOI22_X1 U70510 ( .A1(n105840), .A2(n109516), .B1(n72472), .B2(n84139), .ZN(
        n84914) );
  AOI22_X1 U70511 ( .A1(n105838), .A2(n109507), .B1(n105837), .B2(n109509), 
        .ZN(n84913) );
  NOR4_X1 U70512 ( .A1(n84915), .A2(n84916), .A3(n84917), .A4(n84918), .ZN(
        n84904) );
  OAI21_X1 U70513 ( .B1(n102923), .B2(n84146), .A(n84919), .ZN(n84918) );
  AOI22_X1 U70514 ( .A1(n105835), .A2(n109445), .B1(n84149), .B2(n109448), 
        .ZN(n84919) );
  OAI21_X1 U70515 ( .B1(n101044), .B2(n105833), .A(n84920), .ZN(n84917) );
  AOI22_X1 U70516 ( .A1(n72396), .A2(n105832), .B1(n105831), .B2(n109442), 
        .ZN(n84920) );
  OAI21_X1 U70517 ( .B1(n105830), .B2(n104592), .A(n84921), .ZN(n84916) );
  AOI22_X1 U70518 ( .A1(n72404), .A2(n105829), .B1(n72408), .B2(n105828), .ZN(
        n84921) );
  OAI21_X1 U70519 ( .B1(n102919), .B2(n105827), .A(n84922), .ZN(n84915) );
  AOI22_X1 U70520 ( .A1(n84160), .A2(n109471), .B1(n84161), .B2(n109468), .ZN(
        n84922) );
  AOI22_X1 U70521 ( .A1(n84162), .A2(n109542), .B1(n84163), .B2(n109539), .ZN(
        n84901) );
  NOR4_X1 U70522 ( .A1(n84924), .A2(n84925), .A3(n84926), .A4(n84927), .ZN(
        n84923) );
  NAND2_X1 U70523 ( .A1(n84928), .A2(n84929), .ZN(n84927) );
  AOI22_X1 U70524 ( .A1(n105170), .A2(n109044), .B1(n71832), .B2(n106289), 
        .ZN(n84929) );
  AOI22_X1 U70525 ( .A1(n106282), .A2(n109005), .B1(n106275), .B2(n108982), 
        .ZN(n84928) );
  NAND2_X1 U70526 ( .A1(n84930), .A2(n84931), .ZN(n84926) );
  AOI22_X1 U70527 ( .A1(n84106), .A2(n109061), .B1(n105852), .B2(n109073), 
        .ZN(n84931) );
  AOI22_X1 U70528 ( .A1(n71800), .A2(n105100), .B1(n106746), .B2(n109030), 
        .ZN(n84930) );
  NAND2_X1 U70529 ( .A1(n84932), .A2(n84933), .ZN(n84925) );
  AOI22_X1 U70530 ( .A1(n105851), .A2(n109065), .B1(n84111), .B2(n109057), 
        .ZN(n84933) );
  AOI22_X1 U70531 ( .A1(n84112), .A2(n109069), .B1(n105850), .B2(n108976), 
        .ZN(n84932) );
  NAND2_X1 U70532 ( .A1(n84934), .A2(n84935), .ZN(n84924) );
  AOI21_X1 U70533 ( .B1(n71889), .B2(n84116), .A(n84936), .ZN(n84935) );
  AOI21_X1 U70534 ( .B1(n84937), .B2(n84938), .A(n106324), .ZN(n84936) );
  NOR4_X1 U70535 ( .A1(n84939), .A2(n84940), .A3(n84941), .A4(n84942), .ZN(
        n84938) );
  OAI21_X1 U70536 ( .B1(n102894), .B2(n84124), .A(n84943), .ZN(n84942) );
  AOI22_X1 U70537 ( .A1(n71832), .A2(n105848), .B1(n84127), .B2(n109015), .ZN(
        n84943) );
  OAI21_X1 U70538 ( .B1(n102896), .B2(n105846), .A(n84944), .ZN(n84941) );
  AOI22_X1 U70539 ( .A1(n84130), .A2(n109040), .B1(n71844), .B2(n84131), .ZN(
        n84944) );
  OAI21_X1 U70540 ( .B1(n102892), .B2(n84132), .A(n84945), .ZN(n84940) );
  AOI22_X1 U70541 ( .A1(n84134), .A2(n109030), .B1(n84135), .B2(n109032), .ZN(
        n84945) );
  NAND2_X1 U70542 ( .A1(n84946), .A2(n84947), .ZN(n84939) );
  AOI22_X1 U70543 ( .A1(n105840), .A2(n109053), .B1(n71872), .B2(n84139), .ZN(
        n84947) );
  AOI22_X1 U70544 ( .A1(n105838), .A2(n109044), .B1(n105837), .B2(n109046), 
        .ZN(n84946) );
  NOR4_X1 U70545 ( .A1(n84948), .A2(n84949), .A3(n84950), .A4(n84951), .ZN(
        n84937) );
  OAI21_X1 U70546 ( .B1(n102903), .B2(n105836), .A(n84952), .ZN(n84951) );
  AOI22_X1 U70547 ( .A1(n105835), .A2(n108982), .B1(n84149), .B2(n108985), 
        .ZN(n84952) );
  OAI21_X1 U70548 ( .B1(n101045), .B2(n105833), .A(n84953), .ZN(n84950) );
  AOI22_X1 U70549 ( .A1(n71796), .A2(n105832), .B1(n105831), .B2(n108979), 
        .ZN(n84953) );
  OAI21_X1 U70550 ( .B1(n105830), .B2(n104591), .A(n84954), .ZN(n84949) );
  AOI22_X1 U70551 ( .A1(n71804), .A2(n105829), .B1(n71808), .B2(n105828), .ZN(
        n84954) );
  OAI21_X1 U70552 ( .B1(n102899), .B2(n105827), .A(n84955), .ZN(n84948) );
  AOI22_X1 U70553 ( .A1(n84160), .A2(n109008), .B1(n84161), .B2(n109005), .ZN(
        n84955) );
  AOI22_X1 U70554 ( .A1(n84162), .A2(n109080), .B1(n84163), .B2(n109077), .ZN(
        n84934) );
  NOR4_X1 U70555 ( .A1(n84957), .A2(n84958), .A3(n84959), .A4(n84960), .ZN(
        n84956) );
  NAND2_X1 U70556 ( .A1(n84961), .A2(n84962), .ZN(n84960) );
  AOI22_X1 U70557 ( .A1(n105171), .A2(n109392), .B1(n72281), .B2(n106289), 
        .ZN(n84962) );
  AOI22_X1 U70558 ( .A1(n106283), .A2(n109353), .B1(n106276), .B2(n109330), 
        .ZN(n84961) );
  NAND2_X1 U70559 ( .A1(n84963), .A2(n84964), .ZN(n84959) );
  AOI22_X1 U70560 ( .A1(n84106), .A2(n109408), .B1(n105852), .B2(n109420), 
        .ZN(n84964) );
  AOI22_X1 U70561 ( .A1(n72249), .A2(n105101), .B1(n105175), .B2(n109378), 
        .ZN(n84963) );
  NAND2_X1 U70562 ( .A1(n84965), .A2(n84966), .ZN(n84958) );
  AOI22_X1 U70563 ( .A1(n105851), .A2(n109412), .B1(n84111), .B2(n109404), 
        .ZN(n84966) );
  AOI22_X1 U70564 ( .A1(n84112), .A2(n109416), .B1(n105850), .B2(n109324), 
        .ZN(n84965) );
  NAND2_X1 U70565 ( .A1(n84967), .A2(n84968), .ZN(n84957) );
  AOI21_X1 U70566 ( .B1(n72338), .B2(n84116), .A(n84969), .ZN(n84968) );
  AOI21_X1 U70567 ( .B1(n84970), .B2(n84971), .A(n106324), .ZN(n84969) );
  NOR4_X1 U70568 ( .A1(n84972), .A2(n84973), .A3(n84974), .A4(n84975), .ZN(
        n84971) );
  OAI21_X1 U70569 ( .B1(n102874), .B2(n84124), .A(n84976), .ZN(n84975) );
  AOI22_X1 U70570 ( .A1(n72281), .A2(n105848), .B1(n84127), .B2(n109363), .ZN(
        n84976) );
  OAI21_X1 U70571 ( .B1(n102876), .B2(n105846), .A(n84977), .ZN(n84974) );
  AOI22_X1 U70572 ( .A1(n84130), .A2(n109388), .B1(n72293), .B2(n84131), .ZN(
        n84977) );
  OAI21_X1 U70573 ( .B1(n102872), .B2(n84132), .A(n84978), .ZN(n84973) );
  AOI22_X1 U70574 ( .A1(n84134), .A2(n109378), .B1(n84135), .B2(n109380), .ZN(
        n84978) );
  NAND2_X1 U70575 ( .A1(n84979), .A2(n84980), .ZN(n84972) );
  AOI22_X1 U70576 ( .A1(n105840), .A2(n109401), .B1(n72321), .B2(n84139), .ZN(
        n84980) );
  AOI22_X1 U70577 ( .A1(n105838), .A2(n109392), .B1(n105837), .B2(n109394), 
        .ZN(n84979) );
  NOR4_X1 U70578 ( .A1(n84981), .A2(n84982), .A3(n84983), .A4(n84984), .ZN(
        n84970) );
  OAI21_X1 U70579 ( .B1(n102883), .B2(n105836), .A(n84985), .ZN(n84984) );
  AOI22_X1 U70580 ( .A1(n105835), .A2(n109330), .B1(n84149), .B2(n109333), 
        .ZN(n84985) );
  OAI21_X1 U70581 ( .B1(n101046), .B2(n105833), .A(n84986), .ZN(n84983) );
  AOI22_X1 U70582 ( .A1(n72245), .A2(n105832), .B1(n105831), .B2(n109327), 
        .ZN(n84986) );
  OAI21_X1 U70583 ( .B1(n105830), .B2(n104590), .A(n84987), .ZN(n84982) );
  AOI22_X1 U70584 ( .A1(n72253), .A2(n105829), .B1(n72257), .B2(n105828), .ZN(
        n84987) );
  OAI21_X1 U70585 ( .B1(n102879), .B2(n105827), .A(n84988), .ZN(n84981) );
  AOI22_X1 U70586 ( .A1(n84160), .A2(n109356), .B1(n84161), .B2(n109353), .ZN(
        n84988) );
  AOI22_X1 U70587 ( .A1(n84162), .A2(n109427), .B1(n84163), .B2(n109424), .ZN(
        n84967) );
  NOR4_X1 U70588 ( .A1(n84990), .A2(n84991), .A3(n84992), .A4(n84993), .ZN(
        n84989) );
  NAND2_X1 U70589 ( .A1(n84994), .A2(n84995), .ZN(n84993) );
  AOI22_X1 U70590 ( .A1(n105172), .A2(n109274), .B1(n72130), .B2(n106289), 
        .ZN(n84995) );
  AOI22_X1 U70591 ( .A1(n106282), .A2(n109235), .B1(n106275), .B2(n109212), 
        .ZN(n84994) );
  NAND2_X1 U70592 ( .A1(n84996), .A2(n84997), .ZN(n84992) );
  AOI22_X1 U70593 ( .A1(n84106), .A2(n109289), .B1(n105852), .B2(n109301), 
        .ZN(n84997) );
  AOI22_X1 U70594 ( .A1(n72098), .A2(n81199), .B1(n105173), .B2(n109260), .ZN(
        n84996) );
  NAND2_X1 U70595 ( .A1(n84998), .A2(n84999), .ZN(n84991) );
  AOI22_X1 U70596 ( .A1(n105851), .A2(n109293), .B1(n84111), .B2(n109285), 
        .ZN(n84999) );
  AOI22_X1 U70597 ( .A1(n84112), .A2(n109297), .B1(n105850), .B2(n109206), 
        .ZN(n84998) );
  NAND2_X1 U70598 ( .A1(n85000), .A2(n85001), .ZN(n84990) );
  AOI21_X1 U70599 ( .B1(n72187), .B2(n84116), .A(n85002), .ZN(n85001) );
  AOI21_X1 U70600 ( .B1(n85003), .B2(n85004), .A(n106324), .ZN(n85002) );
  NOR4_X1 U70601 ( .A1(n85005), .A2(n85006), .A3(n85007), .A4(n85008), .ZN(
        n85004) );
  OAI21_X1 U70602 ( .B1(n102854), .B2(n84124), .A(n85009), .ZN(n85008) );
  AOI22_X1 U70603 ( .A1(n72130), .A2(n105848), .B1(n84127), .B2(n109245), .ZN(
        n85009) );
  OAI21_X1 U70604 ( .B1(n102856), .B2(n105846), .A(n85010), .ZN(n85007) );
  AOI22_X1 U70605 ( .A1(n84130), .A2(n109270), .B1(n72142), .B2(n84131), .ZN(
        n85010) );
  OAI21_X1 U70606 ( .B1(n102852), .B2(n84132), .A(n85011), .ZN(n85006) );
  AOI22_X1 U70607 ( .A1(n84134), .A2(n109260), .B1(n84135), .B2(n109262), .ZN(
        n85011) );
  NAND2_X1 U70608 ( .A1(n85012), .A2(n85013), .ZN(n85005) );
  AOI22_X1 U70609 ( .A1(n105840), .A2(n109282), .B1(n72170), .B2(n84139), .ZN(
        n85013) );
  AOI22_X1 U70610 ( .A1(n105838), .A2(n109274), .B1(n105837), .B2(n109276), 
        .ZN(n85012) );
  NOR4_X1 U70611 ( .A1(n85014), .A2(n85015), .A3(n85016), .A4(n85017), .ZN(
        n85003) );
  OAI21_X1 U70612 ( .B1(n102863), .B2(n105836), .A(n85018), .ZN(n85017) );
  AOI22_X1 U70613 ( .A1(n105835), .A2(n109212), .B1(n84149), .B2(n109215), 
        .ZN(n85018) );
  OAI21_X1 U70614 ( .B1(n101047), .B2(n105833), .A(n85019), .ZN(n85016) );
  AOI22_X1 U70615 ( .A1(n72094), .A2(n105832), .B1(n105831), .B2(n109209), 
        .ZN(n85019) );
  OAI21_X1 U70616 ( .B1(n105830), .B2(n104589), .A(n85020), .ZN(n85015) );
  AOI22_X1 U70617 ( .A1(n72102), .A2(n105829), .B1(n72106), .B2(n105828), .ZN(
        n85020) );
  OAI21_X1 U70618 ( .B1(n102859), .B2(n105827), .A(n85021), .ZN(n85014) );
  AOI22_X1 U70619 ( .A1(n84160), .A2(n109238), .B1(n84161), .B2(n109235), .ZN(
        n85021) );
  AOI22_X1 U70620 ( .A1(n84162), .A2(n109308), .B1(n84163), .B2(n109305), .ZN(
        n85000) );
  NOR4_X1 U70621 ( .A1(n85023), .A2(n85024), .A3(n85025), .A4(n85026), .ZN(
        n85022) );
  NAND2_X1 U70622 ( .A1(n85027), .A2(n85028), .ZN(n85026) );
  AOI22_X1 U70623 ( .A1(n106745), .A2(n109165), .B1(n71986), .B2(n106289), 
        .ZN(n85028) );
  AOI22_X1 U70624 ( .A1(n106283), .A2(n109127), .B1(n106276), .B2(n109104), 
        .ZN(n85027) );
  NAND2_X1 U70625 ( .A1(n85029), .A2(n85030), .ZN(n85025) );
  AOI22_X1 U70626 ( .A1(n84106), .A2(n109181), .B1(n105852), .B2(n109193), 
        .ZN(n85030) );
  AOI22_X1 U70627 ( .A1(n71954), .A2(n105101), .B1(n106746), .B2(n109151), 
        .ZN(n85029) );
  NAND2_X1 U70628 ( .A1(n85031), .A2(n85032), .ZN(n85024) );
  AOI22_X1 U70629 ( .A1(n105851), .A2(n109185), .B1(n84111), .B2(n109177), 
        .ZN(n85032) );
  AOI22_X1 U70630 ( .A1(n84112), .A2(n109189), .B1(n105850), .B2(n109098), 
        .ZN(n85031) );
  NAND2_X1 U70631 ( .A1(n85033), .A2(n85034), .ZN(n85023) );
  AOI21_X1 U70632 ( .B1(n72043), .B2(n84116), .A(n85035), .ZN(n85034) );
  AOI21_X1 U70633 ( .B1(n85036), .B2(n85037), .A(n106324), .ZN(n85035) );
  NOR4_X1 U70634 ( .A1(n85038), .A2(n85039), .A3(n85040), .A4(n85041), .ZN(
        n85037) );
  OAI21_X1 U70635 ( .B1(n102834), .B2(n84124), .A(n85042), .ZN(n85041) );
  AOI22_X1 U70636 ( .A1(n71986), .A2(n105848), .B1(n105847), .B2(n109137), 
        .ZN(n85042) );
  OAI21_X1 U70637 ( .B1(n102836), .B2(n105846), .A(n85043), .ZN(n85040) );
  AOI22_X1 U70638 ( .A1(n84130), .A2(n109161), .B1(n71998), .B2(n84131), .ZN(
        n85043) );
  OAI21_X1 U70639 ( .B1(n102832), .B2(n84132), .A(n85044), .ZN(n85039) );
  AOI22_X1 U70640 ( .A1(n84134), .A2(n109151), .B1(n84135), .B2(n109153), .ZN(
        n85044) );
  NAND2_X1 U70641 ( .A1(n85045), .A2(n85046), .ZN(n85038) );
  AOI22_X1 U70642 ( .A1(n105840), .A2(n109174), .B1(n72026), .B2(n84139), .ZN(
        n85046) );
  AOI22_X1 U70643 ( .A1(n105838), .A2(n109165), .B1(n105837), .B2(n109167), 
        .ZN(n85045) );
  NOR4_X1 U70644 ( .A1(n85047), .A2(n85048), .A3(n85049), .A4(n85050), .ZN(
        n85036) );
  OAI21_X1 U70645 ( .B1(n102843), .B2(n105836), .A(n85051), .ZN(n85050) );
  AOI22_X1 U70646 ( .A1(n105835), .A2(n109104), .B1(n84149), .B2(n109107), 
        .ZN(n85051) );
  OAI21_X1 U70647 ( .B1(n101048), .B2(n105833), .A(n85052), .ZN(n85049) );
  AOI22_X1 U70648 ( .A1(n71950), .A2(n105832), .B1(n105831), .B2(n109101), 
        .ZN(n85052) );
  OAI21_X1 U70649 ( .B1(n105830), .B2(n104588), .A(n85053), .ZN(n85048) );
  AOI22_X1 U70650 ( .A1(n71958), .A2(n105829), .B1(n71962), .B2(n105828), .ZN(
        n85053) );
  OAI21_X1 U70651 ( .B1(n102839), .B2(n105827), .A(n85054), .ZN(n85047) );
  AOI22_X1 U70652 ( .A1(n84160), .A2(n109130), .B1(n84161), .B2(n109127), .ZN(
        n85054) );
  AOI22_X1 U70653 ( .A1(n84162), .A2(n109200), .B1(n84163), .B2(n109197), .ZN(
        n85033) );
  NOR4_X1 U70654 ( .A1(n85056), .A2(n85057), .A3(n85058), .A4(n85059), .ZN(
        n85055) );
  NAND2_X1 U70655 ( .A1(n85060), .A2(n85061), .ZN(n85059) );
  AOI22_X1 U70656 ( .A1(n105170), .A2(n108701), .B1(n71388), .B2(n106289), 
        .ZN(n85061) );
  AOI22_X1 U70657 ( .A1(n80260), .A2(n108662), .B1(n81250), .B2(n108639), .ZN(
        n85060) );
  NAND2_X1 U70658 ( .A1(n85062), .A2(n85063), .ZN(n85058) );
  AOI22_X1 U70659 ( .A1(n84106), .A2(n108716), .B1(n105852), .B2(n108728), 
        .ZN(n85063) );
  AOI22_X1 U70660 ( .A1(n71356), .A2(n105099), .B1(n105174), .B2(n108687), 
        .ZN(n85062) );
  NAND2_X1 U70661 ( .A1(n85064), .A2(n85065), .ZN(n85057) );
  AOI22_X1 U70662 ( .A1(n105851), .A2(n108720), .B1(n84111), .B2(n108712), 
        .ZN(n85065) );
  AOI22_X1 U70663 ( .A1(n84112), .A2(n108724), .B1(n105850), .B2(n108633), 
        .ZN(n85064) );
  NAND2_X1 U70664 ( .A1(n85066), .A2(n85067), .ZN(n85056) );
  AOI21_X1 U70665 ( .B1(n71445), .B2(n84116), .A(n85068), .ZN(n85067) );
  AOI21_X1 U70666 ( .B1(n85069), .B2(n85070), .A(n106324), .ZN(n85068) );
  NOR4_X1 U70667 ( .A1(n85071), .A2(n85072), .A3(n85073), .A4(n85074), .ZN(
        n85070) );
  OAI21_X1 U70668 ( .B1(n102814), .B2(n84124), .A(n85075), .ZN(n85074) );
  AOI22_X1 U70669 ( .A1(n71388), .A2(n105848), .B1(n84127), .B2(n108672), .ZN(
        n85075) );
  OAI21_X1 U70670 ( .B1(n102816), .B2(n105846), .A(n85076), .ZN(n85073) );
  AOI22_X1 U70671 ( .A1(n84130), .A2(n108697), .B1(n71400), .B2(n105844), .ZN(
        n85076) );
  OAI21_X1 U70672 ( .B1(n102812), .B2(n84132), .A(n85077), .ZN(n85072) );
  AOI22_X1 U70673 ( .A1(n84134), .A2(n108687), .B1(n84135), .B2(n108689), .ZN(
        n85077) );
  NAND2_X1 U70674 ( .A1(n85078), .A2(n85079), .ZN(n85071) );
  AOI22_X1 U70675 ( .A1(n105840), .A2(n108709), .B1(n71428), .B2(n84139), .ZN(
        n85079) );
  AOI22_X1 U70676 ( .A1(n105838), .A2(n108701), .B1(n105837), .B2(n108703), 
        .ZN(n85078) );
  NOR4_X1 U70677 ( .A1(n85080), .A2(n85081), .A3(n85082), .A4(n85083), .ZN(
        n85069) );
  OAI21_X1 U70678 ( .B1(n102823), .B2(n105836), .A(n85084), .ZN(n85083) );
  AOI22_X1 U70679 ( .A1(n105835), .A2(n108639), .B1(n84149), .B2(n108642), 
        .ZN(n85084) );
  OAI21_X1 U70680 ( .B1(n101049), .B2(n105833), .A(n85085), .ZN(n85082) );
  AOI22_X1 U70681 ( .A1(n71352), .A2(n105832), .B1(n105831), .B2(n108636), 
        .ZN(n85085) );
  OAI21_X1 U70682 ( .B1(n105830), .B2(n104587), .A(n85086), .ZN(n85081) );
  AOI22_X1 U70683 ( .A1(n71360), .A2(n105829), .B1(n71364), .B2(n105828), .ZN(
        n85086) );
  OAI21_X1 U70684 ( .B1(n102819), .B2(n105827), .A(n85087), .ZN(n85080) );
  AOI22_X1 U70685 ( .A1(n84160), .A2(n108665), .B1(n84161), .B2(n108662), .ZN(
        n85087) );
  AOI22_X1 U70686 ( .A1(n84162), .A2(n108735), .B1(n84163), .B2(n108732), .ZN(
        n85066) );
  NOR4_X1 U70687 ( .A1(n85089), .A2(n85090), .A3(n85091), .A4(n85092), .ZN(
        n85088) );
  NAND2_X1 U70688 ( .A1(n85093), .A2(n85094), .ZN(n85092) );
  AOI22_X1 U70689 ( .A1(n105170), .A2(n108928), .B1(n71683), .B2(n106289), 
        .ZN(n85094) );
  AOI22_X1 U70690 ( .A1(n106282), .A2(n108889), .B1(n81250), .B2(n108866), 
        .ZN(n85093) );
  NAND2_X1 U70691 ( .A1(n85095), .A2(n85096), .ZN(n85091) );
  AOI22_X1 U70692 ( .A1(n84106), .A2(n108944), .B1(n105852), .B2(n108956), 
        .ZN(n85096) );
  AOI22_X1 U70693 ( .A1(n71651), .A2(n105101), .B1(n105173), .B2(n108914), 
        .ZN(n85095) );
  NAND2_X1 U70694 ( .A1(n85097), .A2(n85098), .ZN(n85090) );
  AOI22_X1 U70695 ( .A1(n105851), .A2(n108948), .B1(n84111), .B2(n108940), 
        .ZN(n85098) );
  AOI22_X1 U70696 ( .A1(n84112), .A2(n108952), .B1(n105850), .B2(n108860), 
        .ZN(n85097) );
  NAND2_X1 U70697 ( .A1(n85099), .A2(n85100), .ZN(n85089) );
  AOI21_X1 U70698 ( .B1(n71740), .B2(n84116), .A(n85101), .ZN(n85100) );
  AOI21_X1 U70699 ( .B1(n85102), .B2(n85103), .A(n106324), .ZN(n85101) );
  NOR4_X1 U70700 ( .A1(n85104), .A2(n85105), .A3(n85106), .A4(n85107), .ZN(
        n85103) );
  OAI21_X1 U70701 ( .B1(n102794), .B2(n84124), .A(n85108), .ZN(n85107) );
  AOI22_X1 U70702 ( .A1(n71683), .A2(n105848), .B1(n105847), .B2(n108899), 
        .ZN(n85108) );
  OAI21_X1 U70703 ( .B1(n102796), .B2(n105846), .A(n85109), .ZN(n85106) );
  AOI22_X1 U70704 ( .A1(n84130), .A2(n108924), .B1(n71695), .B2(n84131), .ZN(
        n85109) );
  OAI21_X1 U70705 ( .B1(n102792), .B2(n84132), .A(n85110), .ZN(n85105) );
  AOI22_X1 U70706 ( .A1(n84134), .A2(n108914), .B1(n84135), .B2(n108916), .ZN(
        n85110) );
  NAND2_X1 U70707 ( .A1(n85111), .A2(n85112), .ZN(n85104) );
  AOI22_X1 U70708 ( .A1(n105840), .A2(n108937), .B1(n71723), .B2(n84139), .ZN(
        n85112) );
  AOI22_X1 U70709 ( .A1(n105838), .A2(n108928), .B1(n105837), .B2(n108930), 
        .ZN(n85111) );
  NOR4_X1 U70710 ( .A1(n85113), .A2(n85114), .A3(n85115), .A4(n85116), .ZN(
        n85102) );
  OAI21_X1 U70711 ( .B1(n102803), .B2(n105836), .A(n85117), .ZN(n85116) );
  AOI22_X1 U70712 ( .A1(n105835), .A2(n108866), .B1(n84149), .B2(n108869), 
        .ZN(n85117) );
  OAI21_X1 U70713 ( .B1(n101050), .B2(n105833), .A(n85118), .ZN(n85115) );
  AOI22_X1 U70714 ( .A1(n71647), .A2(n105832), .B1(n105831), .B2(n108863), 
        .ZN(n85118) );
  OAI21_X1 U70715 ( .B1(n105830), .B2(n104586), .A(n85119), .ZN(n85114) );
  AOI22_X1 U70716 ( .A1(n71655), .A2(n105829), .B1(n71659), .B2(n105828), .ZN(
        n85119) );
  OAI21_X1 U70717 ( .B1(n102799), .B2(n105827), .A(n85120), .ZN(n85113) );
  AOI22_X1 U70718 ( .A1(n84160), .A2(n108892), .B1(n84161), .B2(n108889), .ZN(
        n85120) );
  AOI22_X1 U70719 ( .A1(n84162), .A2(n108963), .B1(n84163), .B2(n108960), .ZN(
        n85099) );
  NOR4_X1 U70720 ( .A1(n85122), .A2(n85123), .A3(n85124), .A4(n85125), .ZN(
        n85121) );
  NAND2_X1 U70721 ( .A1(n85126), .A2(n85127), .ZN(n85125) );
  AOI22_X1 U70722 ( .A1(n105171), .A2(n108816), .B1(n71539), .B2(n106289), 
        .ZN(n85127) );
  AOI22_X1 U70723 ( .A1(n106284), .A2(n108777), .B1(n81250), .B2(n108754), 
        .ZN(n85126) );
  NAND2_X1 U70724 ( .A1(n85128), .A2(n85129), .ZN(n85124) );
  AOI22_X1 U70725 ( .A1(n84106), .A2(n108832), .B1(n105852), .B2(n108844), 
        .ZN(n85129) );
  AOI22_X1 U70726 ( .A1(n71507), .A2(n105101), .B1(n105173), .B2(n108802), 
        .ZN(n85128) );
  NAND2_X1 U70727 ( .A1(n85130), .A2(n85131), .ZN(n85123) );
  AOI22_X1 U70728 ( .A1(n105851), .A2(n108836), .B1(n84111), .B2(n108828), 
        .ZN(n85131) );
  AOI22_X1 U70729 ( .A1(n84112), .A2(n108840), .B1(n105850), .B2(n108748), 
        .ZN(n85130) );
  NAND2_X1 U70730 ( .A1(n85132), .A2(n85133), .ZN(n85122) );
  AOI21_X1 U70731 ( .B1(n71596), .B2(n84116), .A(n85134), .ZN(n85133) );
  AOI21_X1 U70732 ( .B1(n85135), .B2(n85136), .A(n106324), .ZN(n85134) );
  NOR4_X1 U70733 ( .A1(n85137), .A2(n85138), .A3(n85139), .A4(n85140), .ZN(
        n85136) );
  OAI21_X1 U70734 ( .B1(n102774), .B2(n84124), .A(n85141), .ZN(n85140) );
  AOI22_X1 U70735 ( .A1(n71539), .A2(n105848), .B1(n84127), .B2(n108787), .ZN(
        n85141) );
  OAI21_X1 U70736 ( .B1(n102776), .B2(n105846), .A(n85142), .ZN(n85139) );
  AOI22_X1 U70737 ( .A1(n84130), .A2(n108812), .B1(n71551), .B2(n84131), .ZN(
        n85142) );
  OAI21_X1 U70738 ( .B1(n102772), .B2(n84132), .A(n85143), .ZN(n85138) );
  AOI22_X1 U70739 ( .A1(n84134), .A2(n108802), .B1(n84135), .B2(n108804), .ZN(
        n85143) );
  NAND2_X1 U70740 ( .A1(n85144), .A2(n85145), .ZN(n85137) );
  AOI22_X1 U70741 ( .A1(n105840), .A2(n108825), .B1(n71579), .B2(n84139), .ZN(
        n85145) );
  AOI22_X1 U70742 ( .A1(n105838), .A2(n108816), .B1(n105837), .B2(n108818), 
        .ZN(n85144) );
  NOR4_X1 U70743 ( .A1(n85146), .A2(n85147), .A3(n85148), .A4(n85149), .ZN(
        n85135) );
  OAI21_X1 U70744 ( .B1(n102783), .B2(n105836), .A(n85150), .ZN(n85149) );
  AOI22_X1 U70745 ( .A1(n105835), .A2(n108754), .B1(n84149), .B2(n108757), 
        .ZN(n85150) );
  OAI21_X1 U70746 ( .B1(n101051), .B2(n105833), .A(n85151), .ZN(n85148) );
  AOI22_X1 U70747 ( .A1(n71503), .A2(n105832), .B1(n105831), .B2(n108751), 
        .ZN(n85151) );
  OAI21_X1 U70748 ( .B1(n105830), .B2(n104585), .A(n85152), .ZN(n85147) );
  AOI22_X1 U70749 ( .A1(n71511), .A2(n105829), .B1(n71515), .B2(n105828), .ZN(
        n85152) );
  OAI21_X1 U70750 ( .B1(n102779), .B2(n105827), .A(n85153), .ZN(n85146) );
  AOI22_X1 U70751 ( .A1(n84160), .A2(n108780), .B1(n84161), .B2(n108777), .ZN(
        n85153) );
  AOI22_X1 U70752 ( .A1(n84162), .A2(n108851), .B1(n84163), .B2(n108848), .ZN(
        n85132) );
  NOR4_X1 U70753 ( .A1(n85155), .A2(n85156), .A3(n85157), .A4(n85158), .ZN(
        n85154) );
  NAND2_X1 U70754 ( .A1(n85159), .A2(n85160), .ZN(n85158) );
  AOI22_X1 U70755 ( .A1(n106745), .A2(n107356), .B1(n69648), .B2(n106289), 
        .ZN(n85160) );
  AOI22_X1 U70756 ( .A1(n106285), .A2(n107317), .B1(n81250), .B2(n107294), 
        .ZN(n85159) );
  NAND2_X1 U70757 ( .A1(n85161), .A2(n85162), .ZN(n85157) );
  AOI22_X1 U70758 ( .A1(n105853), .A2(n107203), .B1(n105852), .B2(n107179), 
        .ZN(n85162) );
  OAI21_X1 U70759 ( .B1(n81252), .B2(n85163), .A(n81253), .ZN(n84107) );
  OAI21_X1 U70760 ( .B1(n81254), .B2(n85163), .A(n106761), .ZN(n84106) );
  AOI22_X1 U70761 ( .A1(n69616), .A2(n105101), .B1(n105175), .B2(n107342), 
        .ZN(n85161) );
  NAND2_X1 U70762 ( .A1(n85164), .A2(n85165), .ZN(n85156) );
  AOI22_X1 U70763 ( .A1(n105851), .A2(n107195), .B1(n84111), .B2(n107211), 
        .ZN(n85165) );
  AND2_X2 U70764 ( .A1(n81198), .A2(n85166), .ZN(n84111) );
  NOR2_X1 U70765 ( .A1(n85167), .A2(n85163), .ZN(n84110) );
  OR2_X1 U70766 ( .A1(n106327), .A2(n81228), .ZN(n85167) );
  AOI22_X1 U70767 ( .A1(n84112), .A2(n107187), .B1(n105850), .B2(n107288), 
        .ZN(n85164) );
  NOR2_X1 U70768 ( .A1(n85168), .A2(n85169), .ZN(n84113) );
  NAND2_X1 U70769 ( .A1(n106328), .A2(n106280), .ZN(n85168) );
  AND2_X2 U70770 ( .A1(n81249), .A2(n85166), .ZN(n84112) );
  NAND2_X1 U70771 ( .A1(n85170), .A2(n85171), .ZN(n85155) );
  AOI21_X1 U70772 ( .B1(n69464), .B2(n84116), .A(n85172), .ZN(n85171) );
  AOI21_X1 U70773 ( .B1(n85173), .B2(n85174), .A(n106324), .ZN(n85172) );
  NOR4_X1 U70774 ( .A1(n85175), .A2(n85176), .A3(n85177), .A4(n85178), .ZN(
        n85174) );
  OAI21_X1 U70775 ( .B1(n102754), .B2(n105849), .A(n85179), .ZN(n85178) );
  AOI22_X1 U70776 ( .A1(n69648), .A2(n105848), .B1(n105847), .B2(n107327), 
        .ZN(n85179) );
  NOR2_X1 U70777 ( .A1(n106733), .A2(n81209), .ZN(n84127) );
  NOR2_X1 U70778 ( .A1(n106734), .A2(n107026), .ZN(n84126) );
  NAND2_X1 U70779 ( .A1(n85180), .A2(n81230), .ZN(n84124) );
  OAI21_X1 U70780 ( .B1(n102756), .B2(n105846), .A(n85181), .ZN(n85177) );
  AOI22_X1 U70781 ( .A1(n84130), .A2(n107352), .B1(n69660), .B2(n84131), .ZN(
        n85181) );
  NOR2_X1 U70782 ( .A1(n85182), .A2(n81208), .ZN(n84131) );
  NOR2_X1 U70783 ( .A1(n85182), .A2(n81209), .ZN(n84130) );
  NAND2_X1 U70784 ( .A1(n85183), .A2(n106279), .ZN(n84128) );
  OAI21_X1 U70785 ( .B1(n102752), .B2(n84132), .A(n85184), .ZN(n85176) );
  AOI22_X1 U70786 ( .A1(n84134), .A2(n107342), .B1(n105841), .B2(n107344), 
        .ZN(n85184) );
  NOR2_X1 U70787 ( .A1(n85182), .A2(n107024), .ZN(n84135) );
  NOR2_X1 U70788 ( .A1(n85185), .A2(n107024), .ZN(n84134) );
  NAND2_X1 U70789 ( .A1(n106735), .A2(n106279), .ZN(n84132) );
  NAND2_X1 U70790 ( .A1(n85186), .A2(n85187), .ZN(n85175) );
  AOI22_X1 U70791 ( .A1(n105840), .A2(n107364), .B1(n69688), .B2(n105839), 
        .ZN(n85187) );
  NOR2_X1 U70792 ( .A1(n85188), .A2(n104582), .ZN(n84139) );
  NOR2_X1 U70793 ( .A1(n85188), .A2(n62190), .ZN(n84138) );
  AOI22_X1 U70794 ( .A1(n105838), .A2(n107356), .B1(n105837), .B2(n107358), 
        .ZN(n85186) );
  NOR2_X1 U70795 ( .A1(n85182), .A2(n107026), .ZN(n84141) );
  NAND2_X1 U70796 ( .A1(n85189), .A2(n105058), .ZN(n85182) );
  NOR2_X1 U70797 ( .A1(n62190), .A2(n106697), .ZN(n85189) );
  NOR2_X1 U70798 ( .A1(n85185), .A2(n107026), .ZN(n84140) );
  NOR4_X1 U70799 ( .A1(n85190), .A2(n85191), .A3(n85192), .A4(n85193), .ZN(
        n85173) );
  OAI21_X1 U70800 ( .B1(n102763), .B2(n105836), .A(n85194), .ZN(n85193) );
  AOI22_X1 U70801 ( .A1(n105835), .A2(n107294), .B1(n84149), .B2(n107297), 
        .ZN(n85194) );
  NOR2_X1 U70802 ( .A1(n85195), .A2(n107024), .ZN(n84149) );
  NOR2_X1 U70803 ( .A1(n85169), .A2(n107024), .ZN(n84148) );
  NAND2_X1 U70804 ( .A1(n106736), .A2(n106279), .ZN(n84146) );
  OAI21_X1 U70805 ( .B1(n101052), .B2(n105833), .A(n85196), .ZN(n85192) );
  AOI22_X1 U70806 ( .A1(n69612), .A2(n105832), .B1(n105831), .B2(n107291), 
        .ZN(n85196) );
  NOR2_X1 U70807 ( .A1(n85195), .A2(n81208), .ZN(n84153) );
  NOR2_X1 U70808 ( .A1(n85195), .A2(n81209), .ZN(n84152) );
  NAND2_X1 U70809 ( .A1(n106735), .A2(n106280), .ZN(n84150) );
  NAND2_X1 U70810 ( .A1(n85197), .A2(n105058), .ZN(n85185) );
  NOR2_X1 U70811 ( .A1(n104582), .A2(n106697), .ZN(n85197) );
  OAI21_X1 U70812 ( .B1(n105830), .B2(n104584), .A(n85198), .ZN(n85191) );
  AOI22_X1 U70813 ( .A1(n69620), .A2(n105829), .B1(n69624), .B2(n105828), .ZN(
        n85198) );
  NOR2_X1 U70814 ( .A1(n106734), .A2(n81208), .ZN(n84157) );
  NOR2_X1 U70815 ( .A1(n85195), .A2(n107026), .ZN(n84156) );
  NAND2_X1 U70816 ( .A1(n85199), .A2(n105058), .ZN(n85195) );
  NOR2_X1 U70817 ( .A1(n62190), .A2(n85200), .ZN(n85199) );
  NAND2_X1 U70818 ( .A1(n106736), .A2(n81230), .ZN(n84154) );
  NAND2_X1 U70819 ( .A1(n85201), .A2(n105058), .ZN(n85169) );
  NOR2_X1 U70820 ( .A1(n85200), .A2(n104582), .ZN(n85201) );
  OAI21_X1 U70821 ( .B1(n102759), .B2(n84158), .A(n85202), .ZN(n85190) );
  AOI22_X1 U70822 ( .A1(n105826), .A2(n107320), .B1(n105825), .B2(n107317), 
        .ZN(n85202) );
  NOR2_X1 U70823 ( .A1(n106734), .A2(n107024), .ZN(n84161) );
  NOR2_X1 U70826 ( .A1(n106733), .A2(n107024), .ZN(n84160) );
  NAND2_X1 U70827 ( .A1(n85180), .A2(n106280), .ZN(n84158) );
  AND2_X2 U70830 ( .A1(n85205), .A2(n85166), .ZN(n84116) );
  NOR2_X1 U70831 ( .A1(n85163), .A2(n62190), .ZN(n85166) );
  NOR2_X1 U70832 ( .A1(n80203), .A2(n81209), .ZN(n85205) );
  AOI22_X1 U70833 ( .A1(n84162), .A2(n106767), .B1(n84163), .B2(n107171), .ZN(
        n85170) );
  AND2_X2 U70834 ( .A1(n85206), .A2(n85207), .ZN(n84163) );
  NOR2_X1 U70835 ( .A1(n62190), .A2(n80203), .ZN(n85206) );
  AND2_X2 U70836 ( .A1(n85208), .A2(n85207), .ZN(n84162) );
  OR2_X1 U70838 ( .A1(n85200), .A2(n105058), .ZN(n85163) );
  XOR2_X1 U70839 ( .A(n81238), .B(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ), 
        .Z(n85200) );
  NAND2_X1 U70841 ( .A1(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ), 
        .A2(n81238), .ZN(n85188) );
  NAND4_X2 U70842 ( .A1(n85210), .A2(n85211), .A3(n85212), .A4(n85213), .ZN(
        n58800) );
  NOR3_X1 U70843 ( .A1(n85214), .A2(n85215), .A3(n85216), .ZN(n85213) );
  NOR2_X1 U70844 ( .A1(n102741), .A2(n85217), .ZN(n85216) );
  AOI21_X1 U70845 ( .B1(n85218), .B2(n85219), .A(n106324), .ZN(n85215) );
  NOR4_X1 U70846 ( .A1(n85220), .A2(n85221), .A3(n85222), .A4(n85223), .ZN(
        n85219) );
  OAI21_X1 U70847 ( .B1(n105823), .B2(n104655), .A(n85225), .ZN(n85223) );
  AOI22_X1 U70848 ( .A1(n85226), .A2(n107884), .B1(n85227), .B2(n107888), .ZN(
        n85225) );
  NAND2_X1 U70849 ( .A1(n85228), .A2(n85229), .ZN(n85222) );
  AOI22_X1 U70850 ( .A1(n85230), .A2(n107908), .B1(n105819), .B2(n107895), 
        .ZN(n85229) );
  AOI22_X1 U70851 ( .A1(n85232), .A2(n107890), .B1(n70329), .B2(n105817), .ZN(
        n85228) );
  NAND2_X1 U70852 ( .A1(n85234), .A2(n85235), .ZN(n85221) );
  AOI22_X1 U70853 ( .A1(n105816), .A2(n107899), .B1(n70365), .B2(n105815), 
        .ZN(n85235) );
  AOI22_X1 U70854 ( .A1(n70369), .A2(n85238), .B1(n105813), .B2(n107905), .ZN(
        n85234) );
  NAND2_X1 U70855 ( .A1(n85240), .A2(n85241), .ZN(n85220) );
  AOI22_X1 U70856 ( .A1(n105812), .A2(n107916), .B1(n85243), .B2(n107914), 
        .ZN(n85241) );
  AOI22_X1 U70857 ( .A1(n85244), .A2(n107912), .B1(n105809), .B2(n107920), 
        .ZN(n85240) );
  NOR4_X1 U70858 ( .A1(n85246), .A2(n85247), .A3(n85248), .A4(n85249), .ZN(
        n85218) );
  OAI21_X1 U70859 ( .B1(n102747), .B2(n85250), .A(n85251), .ZN(n85249) );
  AOI22_X1 U70860 ( .A1(n85252), .A2(n107934), .B1(n70424), .B2(n85253), .ZN(
        n85251) );
  NAND2_X1 U70861 ( .A1(n85254), .A2(n85255), .ZN(n85248) );
  AOI22_X1 U70862 ( .A1(n85256), .A2(n70297), .B1(n85257), .B2(n70404), .ZN(
        n85255) );
  AOI22_X1 U70863 ( .A1(n105802), .A2(n107930), .B1(n85259), .B2(n107922), 
        .ZN(n85254) );
  OAI21_X1 U70864 ( .B1(n102745), .B2(n85260), .A(n85261), .ZN(n85247) );
  AOI22_X1 U70865 ( .A1(n105799), .A2(n107856), .B1(n85263), .B2(n107897), 
        .ZN(n85261) );
  NAND2_X1 U70866 ( .A1(n85264), .A2(n85265), .ZN(n85246) );
  AOI22_X1 U70867 ( .A1(n105797), .A2(n107877), .B1(n85267), .B2(n70317), .ZN(
        n85265) );
  AOI22_X1 U70868 ( .A1(n85268), .A2(n107871), .B1(n85269), .B2(n107864), .ZN(
        n85264) );
  NOR2_X1 U70869 ( .A1(n102739), .A2(n85270), .ZN(n85214) );
  AOI22_X1 U70870 ( .A1(n105101), .A2(n70317), .B1(n70365), .B2(n105174), .ZN(
        n85212) );
  AOI22_X1 U70871 ( .A1(n105170), .A2(n107912), .B1(n105792), .B2(n107862), 
        .ZN(n85211) );
  AOI22_X1 U70872 ( .A1(n85272), .A2(n107926), .B1(n85273), .B2(n107938), .ZN(
        n85210) );
  NAND4_X2 U70873 ( .A1(n85274), .A2(n85275), .A3(n85276), .A4(n85277), .ZN(
        n58799) );
  NOR3_X1 U70874 ( .A1(n85278), .A2(n85279), .A3(n85280), .ZN(n85277) );
  NOR2_X1 U70875 ( .A1(n102727), .A2(n85217), .ZN(n85280) );
  AOI21_X1 U70876 ( .B1(n85281), .B2(n85282), .A(n106324), .ZN(n85279) );
  NOR4_X1 U70877 ( .A1(n85283), .A2(n85284), .A3(n85285), .A4(n85286), .ZN(
        n85282) );
  OAI21_X1 U70878 ( .B1(n105823), .B2(n104654), .A(n85287), .ZN(n85286) );
  AOI22_X1 U70879 ( .A1(n85226), .A2(n107979), .B1(n85227), .B2(n107983), .ZN(
        n85287) );
  NAND2_X1 U70880 ( .A1(n85288), .A2(n85289), .ZN(n85285) );
  AOI22_X1 U70881 ( .A1(n85230), .A2(n108004), .B1(n105819), .B2(n107989), 
        .ZN(n85289) );
  AOI22_X1 U70882 ( .A1(n85232), .A2(n107985), .B1(n70471), .B2(n105817), .ZN(
        n85288) );
  NAND2_X1 U70883 ( .A1(n85290), .A2(n85291), .ZN(n85284) );
  AOI22_X1 U70884 ( .A1(n105816), .A2(n107993), .B1(n70507), .B2(n105815), 
        .ZN(n85291) );
  AOI22_X1 U70885 ( .A1(n70511), .A2(n85238), .B1(n105813), .B2(n108001), .ZN(
        n85290) );
  NAND2_X1 U70886 ( .A1(n85292), .A2(n85293), .ZN(n85283) );
  AOI22_X1 U70887 ( .A1(n105812), .A2(n108013), .B1(n85243), .B2(n108010), 
        .ZN(n85293) );
  AOI22_X1 U70888 ( .A1(n85244), .A2(n108008), .B1(n70535), .B2(n105809), .ZN(
        n85292) );
  NOR4_X1 U70889 ( .A1(n85294), .A2(n85295), .A3(n85296), .A4(n85297), .ZN(
        n85281) );
  OAI21_X1 U70890 ( .B1(n102734), .B2(n85250), .A(n85298), .ZN(n85297) );
  AOI22_X1 U70891 ( .A1(n85252), .A2(n108030), .B1(n70566), .B2(n105805), .ZN(
        n85298) );
  NAND2_X1 U70892 ( .A1(n85299), .A2(n85300), .ZN(n85296) );
  AOI22_X1 U70893 ( .A1(n85256), .A2(n70439), .B1(n85257), .B2(n70546), .ZN(
        n85300) );
  AOI22_X1 U70894 ( .A1(n105802), .A2(n108026), .B1(n85259), .B2(n108018), 
        .ZN(n85299) );
  OAI21_X1 U70895 ( .B1(n102733), .B2(n85260), .A(n85301), .ZN(n85295) );
  AOI22_X1 U70896 ( .A1(n105799), .A2(n107953), .B1(n85263), .B2(n107991), 
        .ZN(n85301) );
  NAND2_X1 U70897 ( .A1(n85302), .A2(n85303), .ZN(n85294) );
  AOI22_X1 U70898 ( .A1(n105797), .A2(n107974), .B1(n85267), .B2(n107970), 
        .ZN(n85303) );
  AOI22_X1 U70899 ( .A1(n85268), .A2(n107968), .B1(n85269), .B2(n107961), .ZN(
        n85302) );
  NOR2_X1 U70900 ( .A1(n102725), .A2(n85270), .ZN(n85278) );
  AOI22_X1 U70901 ( .A1(n105100), .A2(n107970), .B1(n70507), .B2(n105175), 
        .ZN(n85276) );
  AOI22_X1 U70902 ( .A1(n105172), .A2(n108008), .B1(n105792), .B2(n107959), 
        .ZN(n85275) );
  AOI22_X1 U70903 ( .A1(n85272), .A2(n108022), .B1(n85273), .B2(n108034), .ZN(
        n85274) );
  NAND4_X2 U70904 ( .A1(n85304), .A2(n85305), .A3(n85306), .A4(n85307), .ZN(
        n58798) );
  NOR3_X1 U70905 ( .A1(n85308), .A2(n85309), .A3(n85310), .ZN(n85307) );
  NOR2_X1 U70906 ( .A1(n102710), .A2(n85217), .ZN(n85310) );
  AOI21_X1 U70907 ( .B1(n85311), .B2(n85312), .A(n106324), .ZN(n85309) );
  NOR4_X1 U70908 ( .A1(n85313), .A2(n85314), .A3(n85315), .A4(n85316), .ZN(
        n85312) );
  OAI21_X1 U70909 ( .B1(n101151), .B2(n105823), .A(n85317), .ZN(n85316) );
  AOI22_X1 U70910 ( .A1(n85226), .A2(n107246), .B1(n85227), .B2(n107250), .ZN(
        n85317) );
  NAND2_X1 U70911 ( .A1(n85318), .A2(n85319), .ZN(n85315) );
  AOI22_X1 U70912 ( .A1(n85230), .A2(n107275), .B1(n105819), .B2(n107258), 
        .ZN(n85319) );
  AOI22_X1 U70913 ( .A1(n85232), .A2(n107253), .B1(n69524), .B2(n105817), .ZN(
        n85318) );
  NAND2_X1 U70914 ( .A1(n85320), .A2(n85321), .ZN(n85314) );
  AOI22_X1 U70915 ( .A1(n105816), .A2(n107263), .B1(n69560), .B2(n105815), 
        .ZN(n85321) );
  AOI22_X1 U70916 ( .A1(n69564), .A2(n105814), .B1(n105813), .B2(n107272), 
        .ZN(n85320) );
  NAND2_X1 U70917 ( .A1(n85322), .A2(n85323), .ZN(n85313) );
  AOI22_X1 U70918 ( .A1(n105812), .A2(n107283), .B1(n85243), .B2(n107281), 
        .ZN(n85323) );
  AOI22_X1 U70919 ( .A1(n85244), .A2(n107279), .B1(n69588), .B2(n105809), .ZN(
        n85322) );
  NOR4_X1 U70920 ( .A1(n85324), .A2(n85325), .A3(n85326), .A4(n85327), .ZN(
        n85311) );
  OAI21_X1 U70921 ( .B1(n102718), .B2(n85250), .A(n85328), .ZN(n85327) );
  AOI22_X1 U70922 ( .A1(n85252), .A2(n107188), .B1(n69425), .B2(n85253), .ZN(
        n85328) );
  NAND2_X1 U70923 ( .A1(n85329), .A2(n85330), .ZN(n85326) );
  AOI22_X1 U70924 ( .A1(n85256), .A2(n69492), .B1(n85257), .B2(n69465), .ZN(
        n85330) );
  AOI22_X1 U70925 ( .A1(n105802), .A2(n107196), .B1(n85259), .B2(n107212), 
        .ZN(n85329) );
  OAI21_X1 U70926 ( .B1(n102716), .B2(n85260), .A(n85331), .ZN(n85325) );
  AOI22_X1 U70927 ( .A1(n105799), .A2(n107215), .B1(n85263), .B2(n107261), 
        .ZN(n85331) );
  NAND2_X1 U70928 ( .A1(n85332), .A2(n85333), .ZN(n85324) );
  AOI22_X1 U70929 ( .A1(n105797), .A2(n107238), .B1(n85267), .B2(n107233), 
        .ZN(n85333) );
  AOI22_X1 U70930 ( .A1(n85268), .A2(n107231), .B1(n85269), .B2(n107224), .ZN(
        n85332) );
  NOR2_X1 U70931 ( .A1(n102708), .A2(n85270), .ZN(n85308) );
  AOI22_X1 U70932 ( .A1(n105101), .A2(n107233), .B1(n69560), .B2(n105173), 
        .ZN(n85306) );
  AOI22_X1 U70933 ( .A1(n106745), .A2(n107279), .B1(n105792), .B2(n107221), 
        .ZN(n85305) );
  AOI22_X1 U70934 ( .A1(n85272), .A2(n107204), .B1(n85273), .B2(n107180), .ZN(
        n85304) );
  NAND4_X2 U70935 ( .A1(n85334), .A2(n85335), .A3(n85336), .A4(n85337), .ZN(
        n58797) );
  NOR3_X1 U70936 ( .A1(n85338), .A2(n85339), .A3(n85340), .ZN(n85337) );
  NOR2_X1 U70937 ( .A1(n102694), .A2(n85217), .ZN(n85340) );
  AOI21_X1 U70938 ( .B1(n85341), .B2(n85342), .A(n106325), .ZN(n85339) );
  NOR4_X1 U70939 ( .A1(n85343), .A2(n85344), .A3(n85345), .A4(n85346), .ZN(
        n85342) );
  OAI21_X1 U70940 ( .B1(n101152), .B2(n105823), .A(n85347), .ZN(n85346) );
  AOI22_X1 U70941 ( .A1(n85226), .A2(n107785), .B1(n85227), .B2(n107789), .ZN(
        n85347) );
  NAND2_X1 U70942 ( .A1(n85348), .A2(n85349), .ZN(n85345) );
  AOI22_X1 U70943 ( .A1(n85230), .A2(n107813), .B1(n70209), .B2(n105819), .ZN(
        n85349) );
  AOI22_X1 U70944 ( .A1(n85232), .A2(n107792), .B1(n70185), .B2(n105817), .ZN(
        n85348) );
  NAND2_X1 U70945 ( .A1(n85350), .A2(n85351), .ZN(n85344) );
  AOI22_X1 U70946 ( .A1(n105816), .A2(n107800), .B1(n85237), .B2(n70221), .ZN(
        n85351) );
  AOI22_X1 U70947 ( .A1(n70225), .A2(n105814), .B1(n105813), .B2(n107809), 
        .ZN(n85350) );
  NAND2_X1 U70948 ( .A1(n85352), .A2(n85353), .ZN(n85343) );
  AOI22_X1 U70949 ( .A1(n105812), .A2(n107821), .B1(n85243), .B2(n107819), 
        .ZN(n85353) );
  AOI22_X1 U70950 ( .A1(n85244), .A2(n107817), .B1(n70249), .B2(n105809), .ZN(
        n85352) );
  NOR4_X1 U70951 ( .A1(n85354), .A2(n85355), .A3(n85356), .A4(n85357), .ZN(
        n85341) );
  OAI21_X1 U70952 ( .B1(n102702), .B2(n85250), .A(n85358), .ZN(n85357) );
  AOI22_X1 U70953 ( .A1(n85252), .A2(n107839), .B1(n70280), .B2(n105805), .ZN(
        n85358) );
  NAND2_X1 U70954 ( .A1(n85359), .A2(n85360), .ZN(n85356) );
  AOI22_X1 U70955 ( .A1(n70153), .A2(n105804), .B1(n85257), .B2(n70260), .ZN(
        n85360) );
  AOI22_X1 U70956 ( .A1(n105802), .A2(n107835), .B1(n85259), .B2(n107826), 
        .ZN(n85359) );
  OAI21_X1 U70957 ( .B1(n102700), .B2(n85260), .A(n85361), .ZN(n85355) );
  AOI22_X1 U70958 ( .A1(n105799), .A2(n107753), .B1(n85263), .B2(n107798), 
        .ZN(n85361) );
  NAND2_X1 U70959 ( .A1(n85362), .A2(n85363), .ZN(n85354) );
  AOI22_X1 U70960 ( .A1(n105797), .A2(n107777), .B1(n85267), .B2(n107771), 
        .ZN(n85363) );
  AOI22_X1 U70961 ( .A1(n85268), .A2(n107769), .B1(n85269), .B2(n107762), .ZN(
        n85362) );
  NOR2_X1 U70962 ( .A1(n101054), .A2(n85270), .ZN(n85338) );
  AOI22_X1 U70963 ( .A1(n105099), .A2(n107771), .B1(n70221), .B2(n106746), 
        .ZN(n85336) );
  AOI22_X1 U70964 ( .A1(n105170), .A2(n107817), .B1(n105792), .B2(n107759), 
        .ZN(n85335) );
  AOI22_X1 U70965 ( .A1(n85272), .A2(n107830), .B1(n85273), .B2(n107843), .ZN(
        n85334) );
  NAND4_X2 U70966 ( .A1(n85364), .A2(n85365), .A3(n85366), .A4(n85367), .ZN(
        n58796) );
  NOR3_X1 U70967 ( .A1(n85368), .A2(n85369), .A3(n85370), .ZN(n85367) );
  NOR2_X1 U70968 ( .A1(n102679), .A2(n85217), .ZN(n85370) );
  AOI21_X1 U70969 ( .B1(n85371), .B2(n85372), .A(n106324), .ZN(n85369) );
  NOR4_X1 U70970 ( .A1(n85373), .A2(n85374), .A3(n85375), .A4(n85376), .ZN(
        n85372) );
  OAI21_X1 U70971 ( .B1(n101153), .B2(n105823), .A(n85377), .ZN(n85376) );
  AOI22_X1 U70972 ( .A1(n85226), .A2(n110686), .B1(n85227), .B2(n110690), .ZN(
        n85377) );
  NAND2_X1 U70973 ( .A1(n85378), .A2(n85379), .ZN(n85375) );
  AOI22_X1 U70974 ( .A1(n85230), .A2(n110709), .B1(n74055), .B2(n105819), .ZN(
        n85379) );
  AOI22_X1 U70975 ( .A1(n85232), .A2(n110692), .B1(n74031), .B2(n105817), .ZN(
        n85378) );
  NAND2_X1 U70976 ( .A1(n85380), .A2(n85381), .ZN(n85374) );
  AOI22_X1 U70977 ( .A1(n105816), .A2(n110699), .B1(n74067), .B2(n105815), 
        .ZN(n85381) );
  AOI22_X1 U70978 ( .A1(n105814), .A2(n74071), .B1(n105813), .B2(n110706), 
        .ZN(n85380) );
  NAND2_X1 U70979 ( .A1(n85382), .A2(n85383), .ZN(n85373) );
  AOI22_X1 U70980 ( .A1(n105812), .A2(n110717), .B1(n85243), .B2(n110715), 
        .ZN(n85383) );
  AOI22_X1 U70981 ( .A1(n85244), .A2(n110713), .B1(n74095), .B2(n105809), .ZN(
        n85382) );
  NOR4_X1 U70982 ( .A1(n85384), .A2(n85385), .A3(n85386), .A4(n85387), .ZN(
        n85371) );
  OAI21_X1 U70983 ( .B1(n102688), .B2(n85250), .A(n85388), .ZN(n85387) );
  AOI22_X1 U70984 ( .A1(n85252), .A2(n110734), .B1(n74126), .B2(n85253), .ZN(
        n85388) );
  NAND2_X1 U70985 ( .A1(n85389), .A2(n85390), .ZN(n85386) );
  AOI22_X1 U70986 ( .A1(n73999), .A2(n105804), .B1(n85257), .B2(n74106), .ZN(
        n85390) );
  AOI22_X1 U70987 ( .A1(n105802), .A2(n110730), .B1(n85259), .B2(n110722), 
        .ZN(n85389) );
  OAI21_X1 U70988 ( .B1(n102686), .B2(n85260), .A(n85391), .ZN(n85385) );
  AOI22_X1 U70989 ( .A1(n105799), .A2(n110656), .B1(n85263), .B2(n110698), 
        .ZN(n85391) );
  NAND2_X1 U70990 ( .A1(n85392), .A2(n85393), .ZN(n85384) );
  AOI22_X1 U70991 ( .A1(n105797), .A2(n110679), .B1(n85267), .B2(n110674), 
        .ZN(n85393) );
  AOI22_X1 U70992 ( .A1(n85268), .A2(n110672), .B1(n85269), .B2(n110665), .ZN(
        n85392) );
  NOR2_X1 U70993 ( .A1(n101055), .A2(n85270), .ZN(n85368) );
  AOI22_X1 U70994 ( .A1(n105101), .A2(n110674), .B1(n74067), .B2(n105175), 
        .ZN(n85366) );
  AOI22_X1 U70995 ( .A1(n105172), .A2(n110713), .B1(n105792), .B2(n110662), 
        .ZN(n85365) );
  AOI22_X1 U70996 ( .A1(n85272), .A2(n110726), .B1(n85273), .B2(n110738), .ZN(
        n85364) );
  NAND4_X2 U70997 ( .A1(n85394), .A2(n85395), .A3(n85396), .A4(n85397), .ZN(
        n58795) );
  NOR3_X1 U70998 ( .A1(n85398), .A2(n85399), .A3(n85400), .ZN(n85397) );
  NOR2_X1 U70999 ( .A1(n102665), .A2(n85217), .ZN(n85400) );
  AOI21_X1 U71000 ( .B1(n85401), .B2(n85402), .A(n106325), .ZN(n85399) );
  NOR4_X1 U71001 ( .A1(n85403), .A2(n85404), .A3(n85405), .A4(n85406), .ZN(
        n85402) );
  OAI21_X1 U71002 ( .B1(n101154), .B2(n105823), .A(n85407), .ZN(n85406) );
  AOI22_X1 U71003 ( .A1(n85226), .A2(n108086), .B1(n85227), .B2(n108090), .ZN(
        n85407) );
  NAND2_X1 U71004 ( .A1(n85408), .A2(n85409), .ZN(n85405) );
  AOI22_X1 U71005 ( .A1(n85230), .A2(n108112), .B1(n105819), .B2(n108097), 
        .ZN(n85409) );
  AOI22_X1 U71006 ( .A1(n85232), .A2(n108092), .B1(n70618), .B2(n105817), .ZN(
        n85408) );
  NAND2_X1 U71007 ( .A1(n85410), .A2(n85411), .ZN(n85404) );
  AOI22_X1 U71008 ( .A1(n105816), .A2(n108102), .B1(n85237), .B2(n70654), .ZN(
        n85411) );
  AOI22_X1 U71009 ( .A1(n70658), .A2(n105814), .B1(n105813), .B2(n108109), 
        .ZN(n85410) );
  NAND2_X1 U71010 ( .A1(n85412), .A2(n85413), .ZN(n85403) );
  AOI22_X1 U71011 ( .A1(n105812), .A2(n108120), .B1(n85243), .B2(n108118), 
        .ZN(n85413) );
  AOI22_X1 U71012 ( .A1(n85244), .A2(n108116), .B1(n105809), .B2(n108124), 
        .ZN(n85412) );
  NOR4_X1 U71013 ( .A1(n85414), .A2(n85415), .A3(n85416), .A4(n85417), .ZN(
        n85401) );
  OAI21_X1 U71014 ( .B1(n102673), .B2(n85250), .A(n85418), .ZN(n85417) );
  AOI22_X1 U71015 ( .A1(n85252), .A2(n108139), .B1(n70713), .B2(n105805), .ZN(
        n85418) );
  NAND2_X1 U71016 ( .A1(n85419), .A2(n85420), .ZN(n85416) );
  AOI22_X1 U71017 ( .A1(n70586), .A2(n105804), .B1(n85257), .B2(n70693), .ZN(
        n85420) );
  AOI22_X1 U71018 ( .A1(n105802), .A2(n108135), .B1(n85259), .B2(n108126), 
        .ZN(n85419) );
  OAI21_X1 U71019 ( .B1(n102672), .B2(n85260), .A(n85421), .ZN(n85415) );
  AOI22_X1 U71020 ( .A1(n105799), .A2(n108055), .B1(n85263), .B2(n108100), 
        .ZN(n85421) );
  NAND2_X1 U71021 ( .A1(n85422), .A2(n85423), .ZN(n85414) );
  AOI22_X1 U71022 ( .A1(n105797), .A2(n108079), .B1(n85267), .B2(n108073), 
        .ZN(n85423) );
  AOI22_X1 U71023 ( .A1(n85268), .A2(n108071), .B1(n85269), .B2(n108064), .ZN(
        n85422) );
  NOR2_X1 U71024 ( .A1(n102663), .A2(n85270), .ZN(n85398) );
  AOI22_X1 U71025 ( .A1(n105101), .A2(n108073), .B1(n70654), .B2(n105175), 
        .ZN(n85396) );
  AOI22_X1 U71026 ( .A1(n106745), .A2(n108116), .B1(n105792), .B2(n108061), 
        .ZN(n85395) );
  AOI22_X1 U71027 ( .A1(n85272), .A2(n108130), .B1(n85273), .B2(n108143), .ZN(
        n85394) );
  NAND4_X2 U71028 ( .A1(n85424), .A2(n85425), .A3(n85426), .A4(n85427), .ZN(
        n58794) );
  NOR3_X1 U71029 ( .A1(n85428), .A2(n85429), .A3(n85430), .ZN(n85427) );
  NOR2_X1 U71030 ( .A1(n102646), .A2(n85217), .ZN(n85430) );
  AOI21_X1 U71031 ( .B1(n85431), .B2(n85432), .A(n106325), .ZN(n85429) );
  NOR4_X1 U71032 ( .A1(n85433), .A2(n85434), .A3(n85435), .A4(n85436), .ZN(
        n85432) );
  OAI21_X1 U71033 ( .B1(n101155), .B2(n105823), .A(n85437), .ZN(n85436) );
  AOI22_X1 U71034 ( .A1(n85226), .A2(n110784), .B1(n85227), .B2(n110788), .ZN(
        n85437) );
  NAND2_X1 U71035 ( .A1(n85438), .A2(n85439), .ZN(n85435) );
  AOI22_X1 U71036 ( .A1(n85230), .A2(n110811), .B1(n74196), .B2(n105819), .ZN(
        n85439) );
  AOI22_X1 U71037 ( .A1(n85232), .A2(n110791), .B1(n74172), .B2(n105817), .ZN(
        n85438) );
  NAND2_X1 U71038 ( .A1(n85440), .A2(n85441), .ZN(n85434) );
  AOI22_X1 U71039 ( .A1(n105816), .A2(n110801), .B1(n74208), .B2(n105815), 
        .ZN(n85441) );
  AOI22_X1 U71040 ( .A1(n74212), .A2(n105814), .B1(n105813), .B2(n110808), 
        .ZN(n85440) );
  NAND2_X1 U71041 ( .A1(n85442), .A2(n85443), .ZN(n85433) );
  AOI22_X1 U71042 ( .A1(n105812), .A2(n110819), .B1(n85243), .B2(n110817), 
        .ZN(n85443) );
  AOI22_X1 U71043 ( .A1(n85244), .A2(n110815), .B1(n105809), .B2(n110823), 
        .ZN(n85442) );
  NOR4_X1 U71044 ( .A1(n85444), .A2(n85445), .A3(n85446), .A4(n85447), .ZN(
        n85431) );
  OAI21_X1 U71045 ( .B1(n102655), .B2(n85250), .A(n85448), .ZN(n85447) );
  AOI22_X1 U71046 ( .A1(n85252), .A2(n110837), .B1(n74267), .B2(n85253), .ZN(
        n85448) );
  NAND2_X1 U71047 ( .A1(n85449), .A2(n85450), .ZN(n85446) );
  AOI22_X1 U71048 ( .A1(n74140), .A2(n105804), .B1(n85257), .B2(n74247), .ZN(
        n85450) );
  AOI22_X1 U71049 ( .A1(n105802), .A2(n110833), .B1(n85259), .B2(n110825), 
        .ZN(n85449) );
  OAI21_X1 U71050 ( .B1(n102653), .B2(n85260), .A(n85451), .ZN(n85445) );
  AOI22_X1 U71051 ( .A1(n105799), .A2(n110753), .B1(n85263), .B2(n110799), 
        .ZN(n85451) );
  NAND2_X1 U71052 ( .A1(n85452), .A2(n85453), .ZN(n85444) );
  AOI22_X1 U71053 ( .A1(n105797), .A2(n110776), .B1(n85267), .B2(n110771), 
        .ZN(n85453) );
  AOI22_X1 U71054 ( .A1(n85268), .A2(n110769), .B1(n85269), .B2(n110762), .ZN(
        n85452) );
  NOR2_X1 U71055 ( .A1(n101056), .A2(n85270), .ZN(n85428) );
  AOI22_X1 U71056 ( .A1(n105100), .A2(n110771), .B1(n74208), .B2(n105175), 
        .ZN(n85426) );
  AOI22_X1 U71057 ( .A1(n105170), .A2(n110815), .B1(n105792), .B2(n110759), 
        .ZN(n85425) );
  AOI22_X1 U71058 ( .A1(n85272), .A2(n110829), .B1(n85273), .B2(n110841), .ZN(
        n85424) );
  NAND4_X2 U71059 ( .A1(n85454), .A2(n85455), .A3(n85456), .A4(n85457), .ZN(
        n58793) );
  NOR3_X1 U71060 ( .A1(n85458), .A2(n85459), .A3(n85460), .ZN(n85457) );
  NOR2_X1 U71061 ( .A1(n102630), .A2(n85217), .ZN(n85460) );
  AOI21_X1 U71062 ( .B1(n85461), .B2(n85462), .A(n106325), .ZN(n85459) );
  NOR4_X1 U71063 ( .A1(n85463), .A2(n85464), .A3(n85465), .A4(n85466), .ZN(
        n85462) );
  OAI21_X1 U71064 ( .B1(n100771), .B2(n105823), .A(n85467), .ZN(n85466) );
  AOI22_X1 U71065 ( .A1(n85226), .A2(n110884), .B1(n85227), .B2(n110888), .ZN(
        n85467) );
  NAND2_X1 U71066 ( .A1(n85468), .A2(n85469), .ZN(n85465) );
  AOI22_X1 U71067 ( .A1(n85230), .A2(n110911), .B1(n74336), .B2(n105819), .ZN(
        n85469) );
  AOI22_X1 U71068 ( .A1(n85232), .A2(n110891), .B1(n74312), .B2(n105817), .ZN(
        n85468) );
  NAND2_X1 U71069 ( .A1(n85470), .A2(n85471), .ZN(n85464) );
  AOI22_X1 U71070 ( .A1(n105816), .A2(n110898), .B1(n74348), .B2(n105815), 
        .ZN(n85471) );
  AOI22_X1 U71071 ( .A1(n105814), .A2(n110903), .B1(n105813), .B2(n110907), 
        .ZN(n85470) );
  NAND2_X1 U71072 ( .A1(n85472), .A2(n85473), .ZN(n85463) );
  AOI22_X1 U71073 ( .A1(n105812), .A2(n110920), .B1(n85243), .B2(n110917), 
        .ZN(n85473) );
  AOI22_X1 U71074 ( .A1(n85244), .A2(n110915), .B1(n105809), .B2(n110924), 
        .ZN(n85472) );
  NOR4_X1 U71075 ( .A1(n85474), .A2(n85475), .A3(n85476), .A4(n85477), .ZN(
        n85461) );
  OAI21_X1 U71076 ( .B1(n102639), .B2(n85250), .A(n85478), .ZN(n85477) );
  AOI22_X1 U71077 ( .A1(n85252), .A2(n110938), .B1(n74407), .B2(n105805), .ZN(
        n85478) );
  NAND2_X1 U71078 ( .A1(n85479), .A2(n85480), .ZN(n85476) );
  AOI22_X1 U71079 ( .A1(n74280), .A2(n105804), .B1(n74387), .B2(n105803), .ZN(
        n85480) );
  AOI22_X1 U71080 ( .A1(n105802), .A2(n110934), .B1(n85259), .B2(n110926), 
        .ZN(n85479) );
  OAI21_X1 U71081 ( .B1(n102637), .B2(n85260), .A(n85481), .ZN(n85475) );
  AOI22_X1 U71082 ( .A1(n105799), .A2(n110854), .B1(n85263), .B2(n110897), 
        .ZN(n85481) );
  NAND2_X1 U71083 ( .A1(n85482), .A2(n85483), .ZN(n85474) );
  AOI22_X1 U71084 ( .A1(n105797), .A2(n110877), .B1(n85267), .B2(n110872), 
        .ZN(n85483) );
  AOI22_X1 U71085 ( .A1(n85268), .A2(n110870), .B1(n85269), .B2(n110863), .ZN(
        n85482) );
  NOR2_X1 U71086 ( .A1(n101057), .A2(n85270), .ZN(n85458) );
  AOI22_X1 U71087 ( .A1(n105099), .A2(n110872), .B1(n74348), .B2(n105175), 
        .ZN(n85456) );
  AOI22_X1 U71088 ( .A1(n105171), .A2(n110915), .B1(n105792), .B2(n110860), 
        .ZN(n85455) );
  AOI22_X1 U71089 ( .A1(n85272), .A2(n110930), .B1(n85273), .B2(n110942), .ZN(
        n85454) );
  NAND4_X2 U71090 ( .A1(n85484), .A2(n85485), .A3(n85486), .A4(n85487), .ZN(
        n58792) );
  NOR3_X1 U71091 ( .A1(n85488), .A2(n85489), .A3(n85490), .ZN(n85487) );
  NOR2_X1 U71092 ( .A1(n102614), .A2(n85217), .ZN(n85490) );
  AOI21_X1 U71093 ( .B1(n85491), .B2(n85492), .A(n106325), .ZN(n85489) );
  NOR4_X1 U71094 ( .A1(n85493), .A2(n85494), .A3(n85495), .A4(n85496), .ZN(
        n85492) );
  OAI21_X1 U71095 ( .B1(n101156), .B2(n105823), .A(n85497), .ZN(n85496) );
  AOI22_X1 U71096 ( .A1(n85226), .A2(n110479), .B1(n85227), .B2(n110482), .ZN(
        n85497) );
  NAND2_X1 U71097 ( .A1(n85498), .A2(n85499), .ZN(n85495) );
  AOI22_X1 U71098 ( .A1(n85230), .A2(n110506), .B1(n73772), .B2(n105819), .ZN(
        n85499) );
  AOI22_X1 U71099 ( .A1(n85232), .A2(n110485), .B1(n73748), .B2(n105817), .ZN(
        n85498) );
  NAND2_X1 U71100 ( .A1(n85500), .A2(n85501), .ZN(n85494) );
  AOI22_X1 U71101 ( .A1(n73780), .A2(n105816), .B1(n85237), .B2(n73784), .ZN(
        n85501) );
  AOI22_X1 U71102 ( .A1(n85238), .A2(n110498), .B1(n105813), .B2(n110502), 
        .ZN(n85500) );
  NAND2_X1 U71103 ( .A1(n85502), .A2(n85503), .ZN(n85493) );
  AOI22_X1 U71104 ( .A1(n105812), .A2(n110514), .B1(n85243), .B2(n110512), 
        .ZN(n85503) );
  AOI22_X1 U71105 ( .A1(n85244), .A2(n110510), .B1(n73812), .B2(n105809), .ZN(
        n85502) );
  NOR4_X1 U71106 ( .A1(n85504), .A2(n85505), .A3(n85506), .A4(n85507), .ZN(
        n85491) );
  OAI21_X1 U71107 ( .B1(n102622), .B2(n85250), .A(n85508), .ZN(n85507) );
  AOI22_X1 U71108 ( .A1(n85252), .A2(n110531), .B1(n73843), .B2(n105805), .ZN(
        n85508) );
  NAND2_X1 U71109 ( .A1(n85509), .A2(n85510), .ZN(n85506) );
  AOI22_X1 U71110 ( .A1(n73716), .A2(n105804), .B1(n73823), .B2(n105803), .ZN(
        n85510) );
  AOI22_X1 U71111 ( .A1(n85258), .A2(n110527), .B1(n85259), .B2(n110519), .ZN(
        n85509) );
  OAI21_X1 U71112 ( .B1(n102620), .B2(n85260), .A(n85511), .ZN(n85505) );
  AOI22_X1 U71113 ( .A1(n85262), .A2(n110449), .B1(n85263), .B2(n110492), .ZN(
        n85511) );
  NAND2_X1 U71114 ( .A1(n85512), .A2(n85513), .ZN(n85504) );
  AOI22_X1 U71115 ( .A1(n73744), .A2(n105797), .B1(n85267), .B2(n110467), .ZN(
        n85513) );
  AOI22_X1 U71116 ( .A1(n85268), .A2(n110465), .B1(n85269), .B2(n110458), .ZN(
        n85512) );
  NOR2_X1 U71117 ( .A1(n101058), .A2(n85270), .ZN(n85488) );
  AOI22_X1 U71118 ( .A1(n105101), .A2(n110467), .B1(n73784), .B2(n105175), 
        .ZN(n85486) );
  AOI22_X1 U71119 ( .A1(n106745), .A2(n110510), .B1(n105792), .B2(n110455), 
        .ZN(n85485) );
  AOI22_X1 U71120 ( .A1(n85272), .A2(n110523), .B1(n85273), .B2(n110535), .ZN(
        n85484) );
  NAND4_X2 U71121 ( .A1(n85514), .A2(n85515), .A3(n85516), .A4(n85517), .ZN(
        n58791) );
  NOR3_X1 U71122 ( .A1(n85518), .A2(n85519), .A3(n85520), .ZN(n85517) );
  NOR2_X1 U71123 ( .A1(n102600), .A2(n85217), .ZN(n85520) );
  AOI21_X1 U71124 ( .B1(n85521), .B2(n85522), .A(n106325), .ZN(n85519) );
  NOR4_X1 U71125 ( .A1(n85523), .A2(n85524), .A3(n85525), .A4(n85526), .ZN(
        n85522) );
  OAI21_X1 U71126 ( .B1(n101157), .B2(n105823), .A(n85527), .ZN(n85526) );
  AOI22_X1 U71127 ( .A1(n85226), .A2(n110261), .B1(n85227), .B2(n110264), .ZN(
        n85527) );
  NAND2_X1 U71128 ( .A1(n85528), .A2(n85529), .ZN(n85525) );
  AOI22_X1 U71129 ( .A1(n85230), .A2(n110289), .B1(n73476), .B2(n105819), .ZN(
        n85529) );
  AOI22_X1 U71130 ( .A1(n85232), .A2(n110267), .B1(n73452), .B2(n105817), .ZN(
        n85528) );
  NAND2_X1 U71131 ( .A1(n85530), .A2(n85531), .ZN(n85524) );
  AOI22_X1 U71132 ( .A1(n73484), .A2(n105816), .B1(n73488), .B2(n105815), .ZN(
        n85531) );
  AOI22_X1 U71133 ( .A1(n105814), .A2(n110281), .B1(n105813), .B2(n110285), 
        .ZN(n85530) );
  NAND2_X1 U71134 ( .A1(n85532), .A2(n85533), .ZN(n85523) );
  AOI22_X1 U71135 ( .A1(n105812), .A2(n110298), .B1(n85243), .B2(n110295), 
        .ZN(n85533) );
  AOI22_X1 U71136 ( .A1(n85244), .A2(n110293), .B1(n105809), .B2(n110302), 
        .ZN(n85532) );
  NOR4_X1 U71137 ( .A1(n85534), .A2(n85535), .A3(n85536), .A4(n85537), .ZN(
        n85521) );
  OAI21_X1 U71138 ( .B1(n102608), .B2(n85250), .A(n85538), .ZN(n85537) );
  AOI22_X1 U71139 ( .A1(n85252), .A2(n110316), .B1(n73547), .B2(n105805), .ZN(
        n85538) );
  NAND2_X1 U71140 ( .A1(n85539), .A2(n85540), .ZN(n85536) );
  AOI22_X1 U71141 ( .A1(n73420), .A2(n105804), .B1(n105803), .B2(n73527), .ZN(
        n85540) );
  AOI22_X1 U71142 ( .A1(n85258), .A2(n110312), .B1(n85259), .B2(n110304), .ZN(
        n85539) );
  OAI21_X1 U71143 ( .B1(n102606), .B2(n85260), .A(n85541), .ZN(n85535) );
  AOI22_X1 U71144 ( .A1(n85262), .A2(n111020), .B1(n85263), .B2(n110275), .ZN(
        n85541) );
  NAND2_X1 U71145 ( .A1(n85542), .A2(n85543), .ZN(n85534) );
  AOI22_X1 U71146 ( .A1(n73448), .A2(n105797), .B1(n85267), .B2(n110249), .ZN(
        n85543) );
  AOI22_X1 U71147 ( .A1(n85268), .A2(n110247), .B1(n85269), .B2(n110240), .ZN(
        n85542) );
  NOR2_X1 U71148 ( .A1(n101059), .A2(n85270), .ZN(n85518) );
  AOI22_X1 U71149 ( .A1(n105100), .A2(n110249), .B1(n73488), .B2(n105175), 
        .ZN(n85516) );
  AOI22_X1 U71150 ( .A1(n105172), .A2(n110293), .B1(n105792), .B2(n110237), 
        .ZN(n85515) );
  AOI22_X1 U71151 ( .A1(n85272), .A2(n110308), .B1(n85273), .B2(n110320), .ZN(
        n85514) );
  NAND4_X2 U71152 ( .A1(n85544), .A2(n85545), .A3(n85546), .A4(n85547), .ZN(
        n58790) );
  NOR3_X1 U71153 ( .A1(n85548), .A2(n85549), .A3(n85550), .ZN(n85547) );
  NOR2_X1 U71154 ( .A1(n102585), .A2(n85217), .ZN(n85550) );
  AOI21_X1 U71155 ( .B1(n85551), .B2(n85552), .A(n106325), .ZN(n85549) );
  NOR4_X1 U71156 ( .A1(n85553), .A2(n85554), .A3(n85555), .A4(n85556), .ZN(
        n85552) );
  OAI21_X1 U71157 ( .B1(n101158), .B2(n105823), .A(n85557), .ZN(n85556) );
  AOI22_X1 U71158 ( .A1(n85226), .A2(n110578), .B1(n85227), .B2(n110582), .ZN(
        n85557) );
  NAND2_X1 U71159 ( .A1(n85558), .A2(n85559), .ZN(n85555) );
  AOI22_X1 U71160 ( .A1(n85230), .A2(n110609), .B1(n73913), .B2(n105819), .ZN(
        n85559) );
  AOI22_X1 U71161 ( .A1(n85232), .A2(n110585), .B1(n73889), .B2(n105817), .ZN(
        n85558) );
  NAND2_X1 U71162 ( .A1(n85560), .A2(n85561), .ZN(n85554) );
  AOI22_X1 U71163 ( .A1(n105816), .A2(n110595), .B1(n85237), .B2(n73925), .ZN(
        n85561) );
  AOI22_X1 U71164 ( .A1(n105814), .A2(n110601), .B1(n105813), .B2(n110605), 
        .ZN(n85560) );
  NAND2_X1 U71165 ( .A1(n85562), .A2(n85563), .ZN(n85553) );
  AOI22_X1 U71166 ( .A1(n105812), .A2(n110619), .B1(n85243), .B2(n110615), 
        .ZN(n85563) );
  AOI22_X1 U71167 ( .A1(n85244), .A2(n110613), .B1(n73953), .B2(n105809), .ZN(
        n85562) );
  NOR4_X1 U71168 ( .A1(n85564), .A2(n85565), .A3(n85566), .A4(n85567), .ZN(
        n85551) );
  OAI21_X1 U71169 ( .B1(n102593), .B2(n85250), .A(n85568), .ZN(n85567) );
  AOI22_X1 U71170 ( .A1(n85252), .A2(n110636), .B1(n73984), .B2(n105805), .ZN(
        n85568) );
  NAND2_X1 U71171 ( .A1(n85569), .A2(n85570), .ZN(n85566) );
  AOI22_X1 U71172 ( .A1(n73857), .A2(n105804), .B1(n73964), .B2(n105803), .ZN(
        n85570) );
  AOI22_X1 U71173 ( .A1(n85258), .A2(n110632), .B1(n85259), .B2(n110624), .ZN(
        n85569) );
  OAI21_X1 U71174 ( .B1(n102591), .B2(n85260), .A(n85571), .ZN(n85565) );
  AOI22_X1 U71175 ( .A1(n85262), .A2(n111018), .B1(n85263), .B2(n110593), .ZN(
        n85571) );
  NAND2_X1 U71176 ( .A1(n85572), .A2(n85573), .ZN(n85564) );
  AOI22_X1 U71177 ( .A1(n73885), .A2(n105797), .B1(n85267), .B2(n110566), .ZN(
        n85573) );
  AOI22_X1 U71178 ( .A1(n85268), .A2(n110564), .B1(n85269), .B2(n110557), .ZN(
        n85572) );
  NOR2_X1 U71179 ( .A1(n101060), .A2(n85270), .ZN(n85548) );
  AOI22_X1 U71180 ( .A1(n105101), .A2(n110566), .B1(n73925), .B2(n105175), 
        .ZN(n85546) );
  AOI22_X1 U71181 ( .A1(n105170), .A2(n110613), .B1(n105792), .B2(n110554), 
        .ZN(n85545) );
  AOI22_X1 U71182 ( .A1(n85272), .A2(n110628), .B1(n85273), .B2(n110640), .ZN(
        n85544) );
  NAND4_X2 U71183 ( .A1(n85574), .A2(n85575), .A3(n85576), .A4(n85577), .ZN(
        n58789) );
  NOR3_X1 U71184 ( .A1(n85578), .A2(n85579), .A3(n85580), .ZN(n85577) );
  NOR2_X1 U71185 ( .A1(n102570), .A2(n105824), .ZN(n85580) );
  AOI21_X1 U71186 ( .B1(n85581), .B2(n85582), .A(n106325), .ZN(n85579) );
  NOR4_X1 U71187 ( .A1(n85583), .A2(n85584), .A3(n85585), .A4(n85586), .ZN(
        n85582) );
  OAI21_X1 U71188 ( .B1(n101159), .B2(n105823), .A(n85587), .ZN(n85586) );
  AOI22_X1 U71189 ( .A1(n105822), .A2(n110369), .B1(n85227), .B2(n110373), 
        .ZN(n85587) );
  NAND2_X1 U71190 ( .A1(n85588), .A2(n85589), .ZN(n85585) );
  AOI22_X1 U71191 ( .A1(n105820), .A2(n110398), .B1(n73625), .B2(n105819), 
        .ZN(n85589) );
  AOI22_X1 U71192 ( .A1(n105818), .A2(n110376), .B1(n73601), .B2(n105817), 
        .ZN(n85588) );
  NAND2_X1 U71193 ( .A1(n85590), .A2(n85591), .ZN(n85584) );
  AOI22_X1 U71194 ( .A1(n105816), .A2(n110385), .B1(n85237), .B2(n73637), .ZN(
        n85591) );
  AOI22_X1 U71195 ( .A1(n105814), .A2(n110390), .B1(n105813), .B2(n110394), 
        .ZN(n85590) );
  NAND2_X1 U71196 ( .A1(n85592), .A2(n85593), .ZN(n85583) );
  AOI22_X1 U71197 ( .A1(n105812), .A2(n110407), .B1(n85243), .B2(n110404), 
        .ZN(n85593) );
  AOI22_X1 U71198 ( .A1(n105810), .A2(n110402), .B1(n105809), .B2(n110411), 
        .ZN(n85592) );
  NOR4_X1 U71199 ( .A1(n85594), .A2(n85595), .A3(n85596), .A4(n85597), .ZN(
        n85581) );
  OAI21_X1 U71200 ( .B1(n102578), .B2(n85250), .A(n85598), .ZN(n85597) );
  AOI22_X1 U71201 ( .A1(n105807), .A2(n110425), .B1(n73696), .B2(n105805), 
        .ZN(n85598) );
  NAND2_X1 U71202 ( .A1(n85599), .A2(n85600), .ZN(n85596) );
  AOI22_X1 U71203 ( .A1(n73569), .A2(n105804), .B1(n105803), .B2(n73676), .ZN(
        n85600) );
  AOI22_X1 U71204 ( .A1(n85258), .A2(n110421), .B1(n85259), .B2(n110413), .ZN(
        n85599) );
  OAI21_X1 U71205 ( .B1(n102576), .B2(n85260), .A(n85601), .ZN(n85595) );
  AOI22_X1 U71206 ( .A1(n85262), .A2(n111019), .B1(n85263), .B2(n110383), .ZN(
        n85601) );
  NAND2_X1 U71207 ( .A1(n85602), .A2(n85603), .ZN(n85594) );
  AOI22_X1 U71208 ( .A1(n73597), .A2(n105797), .B1(n85267), .B2(n110357), .ZN(
        n85603) );
  AOI22_X1 U71209 ( .A1(n105795), .A2(n110355), .B1(n85269), .B2(n110348), 
        .ZN(n85602) );
  NOR2_X1 U71210 ( .A1(n101061), .A2(n105793), .ZN(n85578) );
  AOI22_X1 U71211 ( .A1(n105100), .A2(n110357), .B1(n73637), .B2(n105175), 
        .ZN(n85576) );
  AOI22_X1 U71212 ( .A1(n106745), .A2(n110402), .B1(n105792), .B2(n110345), 
        .ZN(n85575) );
  AOI22_X1 U71213 ( .A1(n105791), .A2(n110417), .B1(n105790), .B2(n110429), 
        .ZN(n85574) );
  NAND4_X2 U71214 ( .A1(n85604), .A2(n85605), .A3(n85606), .A4(n85607), .ZN(
        n58788) );
  NOR3_X1 U71215 ( .A1(n85608), .A2(n85609), .A3(n85610), .ZN(n85607) );
  NOR2_X1 U71216 ( .A1(n102554), .A2(n105824), .ZN(n85610) );
  AOI21_X1 U71217 ( .B1(n85611), .B2(n85612), .A(n106325), .ZN(n85609) );
  NOR4_X1 U71218 ( .A1(n85613), .A2(n85614), .A3(n85615), .A4(n85616), .ZN(
        n85612) );
  OAI21_X1 U71219 ( .B1(n101160), .B2(n85224), .A(n85617), .ZN(n85616) );
  AOI22_X1 U71220 ( .A1(n105822), .A2(n110045), .B1(n105821), .B2(n110049), 
        .ZN(n85617) );
  NAND2_X1 U71221 ( .A1(n85618), .A2(n85619), .ZN(n85615) );
  AOI22_X1 U71222 ( .A1(n105820), .A2(n110076), .B1(n105819), .B2(n110058), 
        .ZN(n85619) );
  AOI22_X1 U71223 ( .A1(n105818), .A2(n110052), .B1(n73163), .B2(n105817), 
        .ZN(n85618) );
  NAND2_X1 U71224 ( .A1(n85620), .A2(n85621), .ZN(n85614) );
  AOI22_X1 U71225 ( .A1(n105816), .A2(n110063), .B1(n73199), .B2(n105815), 
        .ZN(n85621) );
  AOI22_X1 U71226 ( .A1(n85238), .A2(n110068), .B1(n105813), .B2(n110072), 
        .ZN(n85620) );
  NAND2_X1 U71227 ( .A1(n85622), .A2(n85623), .ZN(n85613) );
  AOI22_X1 U71228 ( .A1(n105812), .A2(n110085), .B1(n105811), .B2(n110082), 
        .ZN(n85623) );
  AOI22_X1 U71229 ( .A1(n105810), .A2(n110080), .B1(n105809), .B2(n110089), 
        .ZN(n85622) );
  NOR4_X1 U71230 ( .A1(n85624), .A2(n85625), .A3(n85626), .A4(n85627), .ZN(
        n85611) );
  OAI21_X1 U71231 ( .B1(n102562), .B2(n105808), .A(n85628), .ZN(n85627) );
  AOI22_X1 U71232 ( .A1(n105807), .A2(n110103), .B1(n73258), .B2(n105805), 
        .ZN(n85628) );
  NAND2_X1 U71233 ( .A1(n85629), .A2(n85630), .ZN(n85626) );
  AOI22_X1 U71234 ( .A1(n73131), .A2(n85256), .B1(n85257), .B2(n73238), .ZN(
        n85630) );
  AOI22_X1 U71235 ( .A1(n85258), .A2(n110099), .B1(n105801), .B2(n110091), 
        .ZN(n85629) );
  OAI21_X1 U71236 ( .B1(n102560), .B2(n105800), .A(n85631), .ZN(n85625) );
  AOI22_X1 U71237 ( .A1(n85262), .A2(n110014), .B1(n105798), .B2(n110061), 
        .ZN(n85631) );
  NAND2_X1 U71238 ( .A1(n85632), .A2(n85633), .ZN(n85624) );
  AOI22_X1 U71239 ( .A1(n105797), .A2(n73159), .B1(n105796), .B2(n110032), 
        .ZN(n85633) );
  AOI22_X1 U71240 ( .A1(n105795), .A2(n110030), .B1(n105794), .B2(n110023), 
        .ZN(n85632) );
  NOR2_X1 U71241 ( .A1(n101062), .A2(n105793), .ZN(n85608) );
  AOI22_X1 U71242 ( .A1(n105100), .A2(n110032), .B1(n73199), .B2(n105175), 
        .ZN(n85606) );
  AOI22_X1 U71243 ( .A1(n105171), .A2(n110080), .B1(n105792), .B2(n110020), 
        .ZN(n85605) );
  AOI22_X1 U71244 ( .A1(n105791), .A2(n110095), .B1(n105790), .B2(n110107), 
        .ZN(n85604) );
  NAND4_X2 U71245 ( .A1(n85634), .A2(n85635), .A3(n85636), .A4(n85637), .ZN(
        n58787) );
  NOR3_X1 U71246 ( .A1(n85638), .A2(n85639), .A3(n85640), .ZN(n85637) );
  NOR2_X1 U71247 ( .A1(n102537), .A2(n105824), .ZN(n85640) );
  AOI21_X1 U71248 ( .B1(n85641), .B2(n85642), .A(n106325), .ZN(n85639) );
  NOR4_X1 U71249 ( .A1(n85643), .A2(n85644), .A3(n85645), .A4(n85646), .ZN(
        n85642) );
  OAI21_X1 U71250 ( .B1(n101161), .B2(n105823), .A(n85647), .ZN(n85646) );
  AOI22_X1 U71251 ( .A1(n105822), .A2(n110152), .B1(n105821), .B2(n110156), 
        .ZN(n85647) );
  NAND2_X1 U71252 ( .A1(n85648), .A2(n85649), .ZN(n85645) );
  AOI22_X1 U71253 ( .A1(n105820), .A2(n110183), .B1(n105819), .B2(n110165), 
        .ZN(n85649) );
  AOI22_X1 U71254 ( .A1(n105818), .A2(n110159), .B1(n73305), .B2(n105817), 
        .ZN(n85648) );
  NAND2_X1 U71255 ( .A1(n85650), .A2(n85651), .ZN(n85644) );
  AOI22_X1 U71256 ( .A1(n105816), .A2(n110170), .B1(n105815), .B2(n73341), 
        .ZN(n85651) );
  AOI22_X1 U71257 ( .A1(n85238), .A2(n110175), .B1(n105813), .B2(n110179), 
        .ZN(n85650) );
  NAND2_X1 U71258 ( .A1(n85652), .A2(n85653), .ZN(n85643) );
  AOI22_X1 U71259 ( .A1(n105812), .A2(n110192), .B1(n105811), .B2(n110189), 
        .ZN(n85653) );
  AOI22_X1 U71260 ( .A1(n105810), .A2(n110187), .B1(n105809), .B2(n110196), 
        .ZN(n85652) );
  NOR4_X1 U71261 ( .A1(n85654), .A2(n85655), .A3(n85656), .A4(n85657), .ZN(
        n85641) );
  OAI21_X1 U71262 ( .B1(n102545), .B2(n85250), .A(n85658), .ZN(n85657) );
  AOI22_X1 U71263 ( .A1(n105807), .A2(n110210), .B1(n73400), .B2(n105805), 
        .ZN(n85658) );
  NAND2_X1 U71264 ( .A1(n85659), .A2(n85660), .ZN(n85656) );
  AOI22_X1 U71265 ( .A1(n73273), .A2(n85256), .B1(n105803), .B2(n73380), .ZN(
        n85660) );
  AOI22_X1 U71266 ( .A1(n85258), .A2(n110206), .B1(n105801), .B2(n110198), 
        .ZN(n85659) );
  OAI21_X1 U71267 ( .B1(n102543), .B2(n85260), .A(n85661), .ZN(n85655) );
  AOI22_X1 U71268 ( .A1(n85262), .A2(n111021), .B1(n105798), .B2(n110168), 
        .ZN(n85661) );
  NAND2_X1 U71269 ( .A1(n85662), .A2(n85663), .ZN(n85654) );
  AOI22_X1 U71270 ( .A1(n73301), .A2(n105797), .B1(n105796), .B2(n110139), 
        .ZN(n85663) );
  AOI22_X1 U71271 ( .A1(n105795), .A2(n110137), .B1(n105794), .B2(n110130), 
        .ZN(n85662) );
  NOR2_X1 U71272 ( .A1(n101063), .A2(n105793), .ZN(n85638) );
  AOI22_X1 U71273 ( .A1(n105099), .A2(n110139), .B1(n73341), .B2(n105175), 
        .ZN(n85636) );
  AOI22_X1 U71274 ( .A1(n105170), .A2(n110187), .B1(n105792), .B2(n110127), 
        .ZN(n85635) );
  AOI22_X1 U71275 ( .A1(n105791), .A2(n110202), .B1(n105790), .B2(n110214), 
        .ZN(n85634) );
  NAND4_X2 U71276 ( .A1(n85664), .A2(n85665), .A3(n85666), .A4(n85667), .ZN(
        n58786) );
  NOR3_X1 U71277 ( .A1(n85668), .A2(n85669), .A3(n85670), .ZN(n85667) );
  NOR2_X1 U71278 ( .A1(n102520), .A2(n105824), .ZN(n85670) );
  AOI21_X1 U71279 ( .B1(n85671), .B2(n85672), .A(n106325), .ZN(n85669) );
  NOR4_X1 U71280 ( .A1(n85673), .A2(n85674), .A3(n85675), .A4(n85676), .ZN(
        n85672) );
  OAI21_X1 U71281 ( .B1(n101162), .B2(n85224), .A(n85677), .ZN(n85676) );
  AOI22_X1 U71282 ( .A1(n105822), .A2(n109936), .B1(n105821), .B2(n109940), 
        .ZN(n85677) );
  NAND2_X1 U71283 ( .A1(n85678), .A2(n85679), .ZN(n85675) );
  AOI22_X1 U71284 ( .A1(n105820), .A2(n109968), .B1(n105819), .B2(n109949), 
        .ZN(n85679) );
  AOI22_X1 U71285 ( .A1(n105818), .A2(n109943), .B1(n73021), .B2(n105817), 
        .ZN(n85678) );
  NAND2_X1 U71286 ( .A1(n85680), .A2(n85681), .ZN(n85674) );
  AOI22_X1 U71287 ( .A1(n105816), .A2(n109954), .B1(n105815), .B2(n73057), 
        .ZN(n85681) );
  AOI22_X1 U71288 ( .A1(n85238), .A2(n109960), .B1(n105813), .B2(n109964), 
        .ZN(n85680) );
  NAND2_X1 U71289 ( .A1(n85682), .A2(n85683), .ZN(n85673) );
  AOI22_X1 U71290 ( .A1(n105812), .A2(n109977), .B1(n105811), .B2(n109974), 
        .ZN(n85683) );
  AOI22_X1 U71291 ( .A1(n105810), .A2(n109972), .B1(n105809), .B2(n109981), 
        .ZN(n85682) );
  NOR4_X1 U71292 ( .A1(n85684), .A2(n85685), .A3(n85686), .A4(n85687), .ZN(
        n85671) );
  OAI21_X1 U71293 ( .B1(n102528), .B2(n105808), .A(n85688), .ZN(n85687) );
  AOI22_X1 U71294 ( .A1(n105807), .A2(n109995), .B1(n73116), .B2(n105805), 
        .ZN(n85688) );
  NAND2_X1 U71295 ( .A1(n85689), .A2(n85690), .ZN(n85686) );
  AOI22_X1 U71296 ( .A1(n72989), .A2(n85256), .B1(n73096), .B2(n105803), .ZN(
        n85690) );
  AOI22_X1 U71297 ( .A1(n85258), .A2(n109991), .B1(n105801), .B2(n109983), 
        .ZN(n85689) );
  OAI21_X1 U71298 ( .B1(n102526), .B2(n105800), .A(n85691), .ZN(n85685) );
  AOI22_X1 U71299 ( .A1(n85262), .A2(n109905), .B1(n105798), .B2(n109952), 
        .ZN(n85691) );
  NAND2_X1 U71300 ( .A1(n85692), .A2(n85693), .ZN(n85684) );
  AOI22_X1 U71301 ( .A1(n73017), .A2(n105797), .B1(n105796), .B2(n109923), 
        .ZN(n85693) );
  AOI22_X1 U71302 ( .A1(n105795), .A2(n109921), .B1(n105794), .B2(n109914), 
        .ZN(n85692) );
  NOR2_X1 U71303 ( .A1(n102518), .A2(n105793), .ZN(n85668) );
  AOI22_X1 U71304 ( .A1(n105101), .A2(n109923), .B1(n73057), .B2(n105175), 
        .ZN(n85666) );
  AOI22_X1 U71305 ( .A1(n106745), .A2(n109972), .B1(n105792), .B2(n109911), 
        .ZN(n85665) );
  AOI22_X1 U71306 ( .A1(n105791), .A2(n109987), .B1(n105790), .B2(n109999), 
        .ZN(n85664) );
  NAND4_X2 U71307 ( .A1(n85694), .A2(n85695), .A3(n85696), .A4(n85697), .ZN(
        n58785) );
  NOR3_X1 U71308 ( .A1(n85698), .A2(n85699), .A3(n85700), .ZN(n85697) );
  NOR2_X1 U71309 ( .A1(n102500), .A2(n105824), .ZN(n85700) );
  AOI21_X1 U71310 ( .B1(n85701), .B2(n85702), .A(n106326), .ZN(n85699) );
  NOR4_X1 U71311 ( .A1(n85703), .A2(n85704), .A3(n85705), .A4(n85706), .ZN(
        n85702) );
  OAI21_X1 U71312 ( .B1(n101163), .B2(n105823), .A(n85707), .ZN(n85706) );
  AOI22_X1 U71313 ( .A1(n105822), .A2(n109819), .B1(n105821), .B2(n109823), 
        .ZN(n85707) );
  NAND2_X1 U71314 ( .A1(n85708), .A2(n85709), .ZN(n85705) );
  AOI22_X1 U71315 ( .A1(n105820), .A2(n109851), .B1(n105819), .B2(n109832), 
        .ZN(n85709) );
  AOI22_X1 U71316 ( .A1(n105818), .A2(n109826), .B1(n72871), .B2(n105817), 
        .ZN(n85708) );
  NAND2_X1 U71317 ( .A1(n85710), .A2(n85711), .ZN(n85704) );
  AOI22_X1 U71318 ( .A1(n105816), .A2(n109837), .B1(n105815), .B2(n72907), 
        .ZN(n85711) );
  AOI22_X1 U71319 ( .A1(n85238), .A2(n109843), .B1(n105813), .B2(n109847), 
        .ZN(n85710) );
  NAND2_X1 U71320 ( .A1(n85712), .A2(n85713), .ZN(n85703) );
  AOI22_X1 U71321 ( .A1(n105812), .A2(n109860), .B1(n105811), .B2(n109857), 
        .ZN(n85713) );
  AOI22_X1 U71322 ( .A1(n105810), .A2(n109855), .B1(n105809), .B2(n109864), 
        .ZN(n85712) );
  NOR4_X1 U71323 ( .A1(n85714), .A2(n85715), .A3(n85716), .A4(n85717), .ZN(
        n85701) );
  OAI21_X1 U71324 ( .B1(n102509), .B2(n85250), .A(n85718), .ZN(n85717) );
  AOI22_X1 U71325 ( .A1(n105807), .A2(n109878), .B1(n72966), .B2(n105805), 
        .ZN(n85718) );
  NAND2_X1 U71326 ( .A1(n85719), .A2(n85720), .ZN(n85716) );
  AOI22_X1 U71327 ( .A1(n72839), .A2(n105804), .B1(n72946), .B2(n105803), .ZN(
        n85720) );
  AOI22_X1 U71328 ( .A1(n105802), .A2(n109874), .B1(n105801), .B2(n109866), 
        .ZN(n85719) );
  OAI21_X1 U71329 ( .B1(n102507), .B2(n85260), .A(n85721), .ZN(n85715) );
  AOI22_X1 U71330 ( .A1(n105799), .A2(n109787), .B1(n105798), .B2(n109835), 
        .ZN(n85721) );
  NAND2_X1 U71331 ( .A1(n85722), .A2(n85723), .ZN(n85714) );
  AOI22_X1 U71332 ( .A1(n105797), .A2(n109811), .B1(n105796), .B2(n109805), 
        .ZN(n85723) );
  AOI22_X1 U71333 ( .A1(n105795), .A2(n109803), .B1(n105794), .B2(n109796), 
        .ZN(n85722) );
  NOR2_X1 U71334 ( .A1(n101064), .A2(n105793), .ZN(n85698) );
  AOI22_X1 U71335 ( .A1(n105100), .A2(n109805), .B1(n72907), .B2(n105175), 
        .ZN(n85696) );
  AOI22_X1 U71336 ( .A1(n105172), .A2(n109855), .B1(n105792), .B2(n109793), 
        .ZN(n85695) );
  AOI22_X1 U71337 ( .A1(n105791), .A2(n109870), .B1(n105790), .B2(n109882), 
        .ZN(n85694) );
  NAND4_X2 U71338 ( .A1(n85724), .A2(n85725), .A3(n85726), .A4(n85727), .ZN(
        n58784) );
  NOR3_X1 U71339 ( .A1(n85728), .A2(n85729), .A3(n85730), .ZN(n85727) );
  NOR2_X1 U71340 ( .A1(n102482), .A2(n105824), .ZN(n85730) );
  AOI21_X1 U71341 ( .B1(n85731), .B2(n85732), .A(n106325), .ZN(n85729) );
  NOR4_X1 U71342 ( .A1(n85733), .A2(n85734), .A3(n85735), .A4(n85736), .ZN(
        n85732) );
  OAI21_X1 U71343 ( .B1(n101164), .B2(n85224), .A(n85737), .ZN(n85736) );
  AOI22_X1 U71344 ( .A1(n105822), .A2(n108193), .B1(n105821), .B2(n108197), 
        .ZN(n85737) );
  NAND2_X1 U71345 ( .A1(n85738), .A2(n85739), .ZN(n85735) );
  AOI22_X1 U71346 ( .A1(n105820), .A2(n108225), .B1(n105819), .B2(n108206), 
        .ZN(n85739) );
  AOI22_X1 U71347 ( .A1(n105818), .A2(n108200), .B1(n85233), .B2(n70767), .ZN(
        n85738) );
  NAND2_X1 U71348 ( .A1(n85740), .A2(n85741), .ZN(n85734) );
  AOI22_X1 U71349 ( .A1(n105816), .A2(n108211), .B1(n105815), .B2(n70803), 
        .ZN(n85741) );
  AOI22_X1 U71350 ( .A1(n85238), .A2(n108217), .B1(n105813), .B2(n108221), 
        .ZN(n85740) );
  NAND2_X1 U71351 ( .A1(n85742), .A2(n85743), .ZN(n85733) );
  AOI22_X1 U71352 ( .A1(n105812), .A2(n108234), .B1(n105811), .B2(n108231), 
        .ZN(n85743) );
  AOI22_X1 U71353 ( .A1(n105810), .A2(n108229), .B1(n105809), .B2(n108238), 
        .ZN(n85742) );
  NOR4_X1 U71354 ( .A1(n85744), .A2(n85745), .A3(n85746), .A4(n85747), .ZN(
        n85731) );
  OAI21_X1 U71355 ( .B1(n102491), .B2(n105808), .A(n85748), .ZN(n85747) );
  AOI22_X1 U71356 ( .A1(n105807), .A2(n108252), .B1(n70862), .B2(n105806), 
        .ZN(n85748) );
  NAND2_X1 U71357 ( .A1(n85749), .A2(n85750), .ZN(n85746) );
  AOI22_X1 U71358 ( .A1(n85256), .A2(n70735), .B1(n70842), .B2(n105803), .ZN(
        n85750) );
  AOI22_X1 U71359 ( .A1(n85258), .A2(n108248), .B1(n105801), .B2(n108240), 
        .ZN(n85749) );
  OAI21_X1 U71360 ( .B1(n102489), .B2(n105800), .A(n85751), .ZN(n85745) );
  AOI22_X1 U71361 ( .A1(n85262), .A2(n108161), .B1(n105798), .B2(n108209), 
        .ZN(n85751) );
  NAND2_X1 U71362 ( .A1(n85752), .A2(n85753), .ZN(n85744) );
  AOI22_X1 U71363 ( .A1(n105797), .A2(n108185), .B1(n105796), .B2(n108179), 
        .ZN(n85753) );
  AOI22_X1 U71364 ( .A1(n105795), .A2(n108177), .B1(n105794), .B2(n108170), 
        .ZN(n85752) );
  NOR2_X1 U71365 ( .A1(n101065), .A2(n105793), .ZN(n85728) );
  AOI22_X1 U71366 ( .A1(n105099), .A2(n108179), .B1(n70803), .B2(n105174), 
        .ZN(n85726) );
  AOI22_X1 U71367 ( .A1(n105170), .A2(n108229), .B1(n105792), .B2(n108167), 
        .ZN(n85725) );
  AOI22_X1 U71368 ( .A1(n105791), .A2(n108244), .B1(n105790), .B2(n108256), 
        .ZN(n85724) );
  NAND4_X2 U71369 ( .A1(n85754), .A2(n85755), .A3(n85756), .A4(n85757), .ZN(
        n58783) );
  NOR3_X1 U71370 ( .A1(n85758), .A2(n85759), .A3(n85760), .ZN(n85757) );
  NOR2_X1 U71371 ( .A1(n102464), .A2(n105824), .ZN(n85760) );
  AOI21_X1 U71372 ( .B1(n85761), .B2(n85762), .A(n106326), .ZN(n85759) );
  NOR4_X1 U71373 ( .A1(n85763), .A2(n85764), .A3(n85765), .A4(n85766), .ZN(
        n85762) );
  OAI21_X1 U71374 ( .B1(n101165), .B2(n105823), .A(n85767), .ZN(n85766) );
  AOI22_X1 U71375 ( .A1(n105822), .A2(n108316), .B1(n105821), .B2(n108320), 
        .ZN(n85767) );
  NAND2_X1 U71376 ( .A1(n85768), .A2(n85769), .ZN(n85765) );
  AOI22_X1 U71377 ( .A1(n105820), .A2(n108348), .B1(n105819), .B2(n108329), 
        .ZN(n85769) );
  AOI22_X1 U71378 ( .A1(n105818), .A2(n108323), .B1(n105817), .B2(n70926), 
        .ZN(n85768) );
  NAND2_X1 U71379 ( .A1(n85770), .A2(n85771), .ZN(n85764) );
  AOI22_X1 U71380 ( .A1(n105816), .A2(n108334), .B1(n105815), .B2(n70962), 
        .ZN(n85771) );
  AOI22_X1 U71381 ( .A1(n85238), .A2(n108340), .B1(n105813), .B2(n108344), 
        .ZN(n85770) );
  NAND2_X1 U71382 ( .A1(n85772), .A2(n85773), .ZN(n85763) );
  AOI22_X1 U71383 ( .A1(n85242), .A2(n108357), .B1(n105811), .B2(n108354), 
        .ZN(n85773) );
  AOI22_X1 U71384 ( .A1(n105810), .A2(n108352), .B1(n105809), .B2(n108361), 
        .ZN(n85772) );
  NOR4_X1 U71385 ( .A1(n85774), .A2(n85775), .A3(n85776), .A4(n85777), .ZN(
        n85761) );
  OAI21_X1 U71386 ( .B1(n102473), .B2(n85250), .A(n85778), .ZN(n85777) );
  AOI22_X1 U71387 ( .A1(n105807), .A2(n108375), .B1(n71021), .B2(n105805), 
        .ZN(n85778) );
  NAND2_X1 U71388 ( .A1(n85779), .A2(n85780), .ZN(n85776) );
  AOI22_X1 U71389 ( .A1(n70894), .A2(n105804), .B1(n71001), .B2(n105803), .ZN(
        n85780) );
  AOI22_X1 U71390 ( .A1(n105802), .A2(n108371), .B1(n105801), .B2(n108363), 
        .ZN(n85779) );
  OAI21_X1 U71391 ( .B1(n102471), .B2(n85260), .A(n85781), .ZN(n85775) );
  AOI22_X1 U71392 ( .A1(n105799), .A2(n108284), .B1(n105798), .B2(n108332), 
        .ZN(n85781) );
  NAND2_X1 U71393 ( .A1(n85782), .A2(n85783), .ZN(n85774) );
  AOI22_X1 U71394 ( .A1(n105797), .A2(n108308), .B1(n105796), .B2(n108302), 
        .ZN(n85783) );
  AOI22_X1 U71395 ( .A1(n105795), .A2(n108300), .B1(n105794), .B2(n108293), 
        .ZN(n85782) );
  NOR2_X1 U71396 ( .A1(n102462), .A2(n105793), .ZN(n85758) );
  AOI22_X1 U71397 ( .A1(n105101), .A2(n108302), .B1(n70962), .B2(n105174), 
        .ZN(n85756) );
  AOI22_X1 U71398 ( .A1(n106745), .A2(n108352), .B1(n105792), .B2(n108290), 
        .ZN(n85755) );
  AOI22_X1 U71399 ( .A1(n105791), .A2(n108367), .B1(n105790), .B2(n108379), 
        .ZN(n85754) );
  NAND4_X2 U71400 ( .A1(n85784), .A2(n85785), .A3(n85786), .A4(n85787), .ZN(
        n58782) );
  NOR3_X1 U71401 ( .A1(n85788), .A2(n85789), .A3(n85790), .ZN(n85787) );
  NOR2_X1 U71402 ( .A1(n102444), .A2(n105824), .ZN(n85790) );
  AOI21_X1 U71403 ( .B1(n85791), .B2(n85792), .A(n106326), .ZN(n85789) );
  NOR4_X1 U71404 ( .A1(n85793), .A2(n85794), .A3(n85795), .A4(n85796), .ZN(
        n85792) );
  OAI21_X1 U71405 ( .B1(n101166), .B2(n85224), .A(n85797), .ZN(n85796) );
  AOI22_X1 U71406 ( .A1(n105822), .A2(n108427), .B1(n105821), .B2(n108431), 
        .ZN(n85797) );
  NAND2_X1 U71407 ( .A1(n85798), .A2(n85799), .ZN(n85795) );
  AOI22_X1 U71408 ( .A1(n105820), .A2(n108459), .B1(n105819), .B2(n108440), 
        .ZN(n85799) );
  AOI22_X1 U71409 ( .A1(n105818), .A2(n108434), .B1(n71071), .B2(n105817), 
        .ZN(n85798) );
  NAND2_X1 U71410 ( .A1(n85800), .A2(n85801), .ZN(n85794) );
  AOI22_X1 U71411 ( .A1(n105816), .A2(n108445), .B1(n105815), .B2(n71107), 
        .ZN(n85801) );
  AOI22_X1 U71412 ( .A1(n105814), .A2(n108451), .B1(n105813), .B2(n108455), 
        .ZN(n85800) );
  NAND2_X1 U71413 ( .A1(n85802), .A2(n85803), .ZN(n85793) );
  AOI22_X1 U71414 ( .A1(n85242), .A2(n108468), .B1(n105811), .B2(n108465), 
        .ZN(n85803) );
  AOI22_X1 U71415 ( .A1(n105810), .A2(n108463), .B1(n105809), .B2(n108472), 
        .ZN(n85802) );
  NOR4_X1 U71416 ( .A1(n85804), .A2(n85805), .A3(n85806), .A4(n85807), .ZN(
        n85791) );
  OAI21_X1 U71417 ( .B1(n102453), .B2(n105808), .A(n85808), .ZN(n85807) );
  AOI22_X1 U71418 ( .A1(n105807), .A2(n108486), .B1(n71166), .B2(n105806), 
        .ZN(n85808) );
  NAND2_X1 U71419 ( .A1(n85809), .A2(n85810), .ZN(n85806) );
  AOI22_X1 U71420 ( .A1(n71039), .A2(n105804), .B1(n71146), .B2(n105803), .ZN(
        n85810) );
  AOI22_X1 U71421 ( .A1(n85258), .A2(n108482), .B1(n105801), .B2(n108474), 
        .ZN(n85809) );
  OAI21_X1 U71422 ( .B1(n102451), .B2(n105800), .A(n85811), .ZN(n85805) );
  AOI22_X1 U71423 ( .A1(n85262), .A2(n108395), .B1(n105798), .B2(n108443), 
        .ZN(n85811) );
  NAND2_X1 U71424 ( .A1(n85812), .A2(n85813), .ZN(n85804) );
  AOI22_X1 U71425 ( .A1(n105797), .A2(n108419), .B1(n105796), .B2(n108413), 
        .ZN(n85813) );
  AOI22_X1 U71426 ( .A1(n105795), .A2(n108411), .B1(n105794), .B2(n108404), 
        .ZN(n85812) );
  NOR2_X1 U71427 ( .A1(n101066), .A2(n105793), .ZN(n85788) );
  AOI22_X1 U71428 ( .A1(n105099), .A2(n108413), .B1(n71107), .B2(n105174), 
        .ZN(n85786) );
  AOI22_X1 U71429 ( .A1(n106745), .A2(n108463), .B1(n105792), .B2(n108401), 
        .ZN(n85785) );
  AOI22_X1 U71430 ( .A1(n105791), .A2(n108478), .B1(n105790), .B2(n108490), 
        .ZN(n85784) );
  NAND4_X2 U71431 ( .A1(n85814), .A2(n85815), .A3(n85816), .A4(n85817), .ZN(
        n58781) );
  NOR3_X1 U71432 ( .A1(n85818), .A2(n85819), .A3(n85820), .ZN(n85817) );
  NOR2_X1 U71433 ( .A1(n102426), .A2(n105824), .ZN(n85820) );
  AOI21_X1 U71434 ( .B1(n85821), .B2(n85822), .A(n106326), .ZN(n85819) );
  NOR4_X1 U71435 ( .A1(n85823), .A2(n85824), .A3(n85825), .A4(n85826), .ZN(
        n85822) );
  OAI21_X1 U71436 ( .B1(n101167), .B2(n105823), .A(n85827), .ZN(n85826) );
  AOI22_X1 U71437 ( .A1(n105822), .A2(n107665), .B1(n105821), .B2(n107669), 
        .ZN(n85827) );
  NAND2_X1 U71438 ( .A1(n85828), .A2(n85829), .ZN(n85825) );
  AOI22_X1 U71439 ( .A1(n105820), .A2(n107697), .B1(n85231), .B2(n107678), 
        .ZN(n85829) );
  AOI22_X1 U71440 ( .A1(n105818), .A2(n107672), .B1(n70032), .B2(n85233), .ZN(
        n85828) );
  NAND2_X1 U71441 ( .A1(n85830), .A2(n85831), .ZN(n85824) );
  AOI22_X1 U71442 ( .A1(n105816), .A2(n107683), .B1(n70068), .B2(n105815), 
        .ZN(n85831) );
  AOI22_X1 U71443 ( .A1(n85238), .A2(n107689), .B1(n105813), .B2(n107693), 
        .ZN(n85830) );
  NAND2_X1 U71444 ( .A1(n85832), .A2(n85833), .ZN(n85823) );
  AOI22_X1 U71445 ( .A1(n85242), .A2(n107706), .B1(n105811), .B2(n107703), 
        .ZN(n85833) );
  AOI22_X1 U71446 ( .A1(n105810), .A2(n107701), .B1(n85245), .B2(n107710), 
        .ZN(n85832) );
  NOR4_X1 U71447 ( .A1(n85834), .A2(n85835), .A3(n85836), .A4(n85837), .ZN(
        n85821) );
  OAI21_X1 U71448 ( .B1(n102435), .B2(n85250), .A(n85838), .ZN(n85837) );
  AOI22_X1 U71449 ( .A1(n105807), .A2(n107723), .B1(n70127), .B2(n105805), 
        .ZN(n85838) );
  NAND2_X1 U71450 ( .A1(n85839), .A2(n85840), .ZN(n85836) );
  AOI22_X1 U71451 ( .A1(n70000), .A2(n105804), .B1(n70107), .B2(n105803), .ZN(
        n85840) );
  AOI22_X1 U71452 ( .A1(n105802), .A2(n107719), .B1(n105801), .B2(n107711), 
        .ZN(n85839) );
  OAI21_X1 U71453 ( .B1(n102433), .B2(n85260), .A(n85841), .ZN(n85835) );
  AOI22_X1 U71454 ( .A1(n105799), .A2(n107633), .B1(n105798), .B2(n107681), 
        .ZN(n85841) );
  NAND2_X1 U71455 ( .A1(n85842), .A2(n85843), .ZN(n85834) );
  AOI22_X1 U71456 ( .A1(n105797), .A2(n107657), .B1(n105796), .B2(n107651), 
        .ZN(n85843) );
  AOI22_X1 U71457 ( .A1(n105795), .A2(n107649), .B1(n105794), .B2(n107642), 
        .ZN(n85842) );
  NOR2_X1 U71458 ( .A1(n102424), .A2(n105793), .ZN(n85818) );
  AOI22_X1 U71459 ( .A1(n105100), .A2(n107651), .B1(n70068), .B2(n105174), 
        .ZN(n85816) );
  AOI22_X1 U71460 ( .A1(n105170), .A2(n107701), .B1(n105792), .B2(n107639), 
        .ZN(n85815) );
  AOI22_X1 U71461 ( .A1(n105791), .A2(n107715), .B1(n105790), .B2(n107727), 
        .ZN(n85814) );
  NAND4_X2 U71462 ( .A1(n85844), .A2(n85845), .A3(n85846), .A4(n85847), .ZN(
        n58780) );
  NOR3_X1 U71463 ( .A1(n85848), .A2(n85849), .A3(n85850), .ZN(n85847) );
  NOR2_X1 U71464 ( .A1(n102406), .A2(n105824), .ZN(n85850) );
  AOI21_X1 U71465 ( .B1(n85851), .B2(n85852), .A(n106326), .ZN(n85849) );
  NOR4_X1 U71466 ( .A1(n85853), .A2(n85854), .A3(n85855), .A4(n85856), .ZN(
        n85852) );
  OAI21_X1 U71467 ( .B1(n101168), .B2(n85224), .A(n85857), .ZN(n85856) );
  AOI22_X1 U71468 ( .A1(n105822), .A2(n109583), .B1(n105821), .B2(n109587), 
        .ZN(n85857) );
  NAND2_X1 U71469 ( .A1(n85858), .A2(n85859), .ZN(n85855) );
  AOI22_X1 U71470 ( .A1(n105820), .A2(n109612), .B1(n85231), .B2(n109596), 
        .ZN(n85859) );
  AOI22_X1 U71471 ( .A1(n105818), .A2(n109590), .B1(n72561), .B2(n105817), 
        .ZN(n85858) );
  NAND2_X1 U71472 ( .A1(n85860), .A2(n85861), .ZN(n85854) );
  AOI22_X1 U71473 ( .A1(n85236), .A2(n109601), .B1(n105815), .B2(n72597), .ZN(
        n85861) );
  AOI22_X1 U71474 ( .A1(n105814), .A2(n109606), .B1(n85239), .B2(n109609), 
        .ZN(n85860) );
  NAND2_X1 U71475 ( .A1(n85862), .A2(n85863), .ZN(n85853) );
  AOI22_X1 U71476 ( .A1(n85242), .A2(n109621), .B1(n105811), .B2(n109618), 
        .ZN(n85863) );
  AOI22_X1 U71477 ( .A1(n105810), .A2(n109616), .B1(n85245), .B2(n109625), 
        .ZN(n85862) );
  NOR4_X1 U71478 ( .A1(n85864), .A2(n85865), .A3(n85866), .A4(n85867), .ZN(
        n85851) );
  OAI21_X1 U71479 ( .B1(n102415), .B2(n105808), .A(n85868), .ZN(n85867) );
  AOI22_X1 U71480 ( .A1(n105807), .A2(n109638), .B1(n72656), .B2(n105806), 
        .ZN(n85868) );
  NAND2_X1 U71481 ( .A1(n85869), .A2(n85870), .ZN(n85866) );
  AOI22_X1 U71482 ( .A1(n72529), .A2(n105804), .B1(n72636), .B2(n105803), .ZN(
        n85870) );
  AOI22_X1 U71483 ( .A1(n85258), .A2(n109634), .B1(n105801), .B2(n109626), 
        .ZN(n85869) );
  OAI21_X1 U71484 ( .B1(n102413), .B2(n105800), .A(n85871), .ZN(n85865) );
  AOI22_X1 U71485 ( .A1(n85262), .A2(n109551), .B1(n105798), .B2(n109599), 
        .ZN(n85871) );
  NAND2_X1 U71486 ( .A1(n85872), .A2(n85873), .ZN(n85864) );
  AOI22_X1 U71487 ( .A1(n85266), .A2(n109575), .B1(n105796), .B2(n109569), 
        .ZN(n85873) );
  AOI22_X1 U71488 ( .A1(n105795), .A2(n109567), .B1(n105794), .B2(n109560), 
        .ZN(n85872) );
  NOR2_X1 U71489 ( .A1(n102404), .A2(n105793), .ZN(n85848) );
  AOI22_X1 U71490 ( .A1(n105100), .A2(n109569), .B1(n72597), .B2(n105174), 
        .ZN(n85846) );
  AOI22_X1 U71491 ( .A1(n106745), .A2(n109616), .B1(n85271), .B2(n109557), 
        .ZN(n85845) );
  AOI22_X1 U71492 ( .A1(n105791), .A2(n109630), .B1(n105790), .B2(n109642), 
        .ZN(n85844) );
  NAND4_X2 U71493 ( .A1(n85874), .A2(n85875), .A3(n85876), .A4(n85877), .ZN(
        n58779) );
  NOR3_X1 U71494 ( .A1(n85878), .A2(n85879), .A3(n85880), .ZN(n85877) );
  NOR2_X1 U71495 ( .A1(n102386), .A2(n105824), .ZN(n85880) );
  AOI21_X1 U71496 ( .B1(n85881), .B2(n85882), .A(n106326), .ZN(n85879) );
  NOR4_X1 U71497 ( .A1(n85883), .A2(n85884), .A3(n85885), .A4(n85886), .ZN(
        n85882) );
  OAI21_X1 U71498 ( .B1(n101169), .B2(n85224), .A(n85887), .ZN(n85886) );
  AOI22_X1 U71499 ( .A1(n105822), .A2(n108544), .B1(n105821), .B2(n108548), 
        .ZN(n85887) );
  NAND2_X1 U71500 ( .A1(n85888), .A2(n85889), .ZN(n85885) );
  AOI22_X1 U71501 ( .A1(n105820), .A2(n108574), .B1(n85231), .B2(n108557), 
        .ZN(n85889) );
  AOI22_X1 U71502 ( .A1(n105818), .A2(n108551), .B1(n85233), .B2(n71220), .ZN(
        n85888) );
  NAND2_X1 U71503 ( .A1(n85890), .A2(n85891), .ZN(n85884) );
  AOI22_X1 U71504 ( .A1(n85236), .A2(n108562), .B1(n105815), .B2(n71256), .ZN(
        n85891) );
  AOI22_X1 U71505 ( .A1(n85238), .A2(n108568), .B1(n85239), .B2(n108571), .ZN(
        n85890) );
  NAND2_X1 U71506 ( .A1(n85892), .A2(n85893), .ZN(n85883) );
  AOI22_X1 U71507 ( .A1(n85242), .A2(n108583), .B1(n105811), .B2(n108580), 
        .ZN(n85893) );
  AOI22_X1 U71508 ( .A1(n105810), .A2(n108578), .B1(n85245), .B2(n108587), 
        .ZN(n85892) );
  NOR4_X1 U71509 ( .A1(n85894), .A2(n85895), .A3(n85896), .A4(n85897), .ZN(
        n85881) );
  OAI21_X1 U71510 ( .B1(n102395), .B2(n105808), .A(n85898), .ZN(n85897) );
  AOI22_X1 U71511 ( .A1(n105807), .A2(n108600), .B1(n71315), .B2(n105806), 
        .ZN(n85898) );
  NAND2_X1 U71512 ( .A1(n85899), .A2(n85900), .ZN(n85896) );
  AOI22_X1 U71513 ( .A1(n71188), .A2(n105804), .B1(n71295), .B2(n105803), .ZN(
        n85900) );
  AOI22_X1 U71514 ( .A1(n85258), .A2(n108596), .B1(n105801), .B2(n108588), 
        .ZN(n85899) );
  OAI21_X1 U71515 ( .B1(n102393), .B2(n105800), .A(n85901), .ZN(n85895) );
  AOI22_X1 U71516 ( .A1(n85262), .A2(n108512), .B1(n105798), .B2(n108560), 
        .ZN(n85901) );
  NAND2_X1 U71517 ( .A1(n85902), .A2(n85903), .ZN(n85894) );
  AOI22_X1 U71518 ( .A1(n85266), .A2(n108536), .B1(n105796), .B2(n108530), 
        .ZN(n85903) );
  AOI22_X1 U71519 ( .A1(n105795), .A2(n108528), .B1(n105794), .B2(n108521), 
        .ZN(n85902) );
  NOR2_X1 U71520 ( .A1(n102384), .A2(n105793), .ZN(n85878) );
  AOI22_X1 U71521 ( .A1(n105101), .A2(n108530), .B1(n71256), .B2(n105174), 
        .ZN(n85876) );
  AOI22_X1 U71522 ( .A1(n106745), .A2(n108578), .B1(n85271), .B2(n108518), 
        .ZN(n85875) );
  AOI22_X1 U71523 ( .A1(n105791), .A2(n108592), .B1(n105790), .B2(n108604), 
        .ZN(n85874) );
  NAND4_X2 U71524 ( .A1(n85904), .A2(n85905), .A3(n85906), .A4(n85907), .ZN(
        n58778) );
  NOR3_X1 U71525 ( .A1(n85908), .A2(n85909), .A3(n85910), .ZN(n85907) );
  NOR2_X1 U71526 ( .A1(n102366), .A2(n105824), .ZN(n85910) );
  AOI21_X1 U71527 ( .B1(n85911), .B2(n85912), .A(n106326), .ZN(n85909) );
  NOR4_X1 U71528 ( .A1(n85913), .A2(n85914), .A3(n85915), .A4(n85916), .ZN(
        n85912) );
  OAI21_X1 U71529 ( .B1(n101170), .B2(n85224), .A(n85917), .ZN(n85916) );
  AOI22_X1 U71530 ( .A1(n105822), .A2(n109688), .B1(n105821), .B2(n109692), 
        .ZN(n85917) );
  NAND2_X1 U71531 ( .A1(n85918), .A2(n85919), .ZN(n85915) );
  AOI22_X1 U71532 ( .A1(n105820), .A2(n109719), .B1(n85231), .B2(n109701), 
        .ZN(n85919) );
  AOI22_X1 U71533 ( .A1(n105818), .A2(n109695), .B1(n72703), .B2(n85233), .ZN(
        n85918) );
  NAND2_X1 U71534 ( .A1(n85920), .A2(n85921), .ZN(n85914) );
  AOI22_X1 U71535 ( .A1(n85236), .A2(n109706), .B1(n72739), .B2(n105815), .ZN(
        n85921) );
  AOI22_X1 U71536 ( .A1(n105814), .A2(n109712), .B1(n85239), .B2(n109715), 
        .ZN(n85920) );
  NAND2_X1 U71537 ( .A1(n85922), .A2(n85923), .ZN(n85913) );
  AOI22_X1 U71538 ( .A1(n85242), .A2(n109728), .B1(n105811), .B2(n109725), 
        .ZN(n85923) );
  AOI22_X1 U71539 ( .A1(n105810), .A2(n109723), .B1(n85245), .B2(n109732), 
        .ZN(n85922) );
  NOR4_X1 U71540 ( .A1(n85924), .A2(n85925), .A3(n85926), .A4(n85927), .ZN(
        n85911) );
  OAI21_X1 U71541 ( .B1(n102375), .B2(n105808), .A(n85928), .ZN(n85927) );
  AOI22_X1 U71542 ( .A1(n105807), .A2(n109745), .B1(n72798), .B2(n105806), 
        .ZN(n85928) );
  NAND2_X1 U71543 ( .A1(n85929), .A2(n85930), .ZN(n85926) );
  AOI22_X1 U71544 ( .A1(n72671), .A2(n105804), .B1(n72778), .B2(n105803), .ZN(
        n85930) );
  AOI22_X1 U71545 ( .A1(n105802), .A2(n109741), .B1(n105801), .B2(n109733), 
        .ZN(n85929) );
  OAI21_X1 U71546 ( .B1(n102373), .B2(n105800), .A(n85931), .ZN(n85925) );
  AOI22_X1 U71547 ( .A1(n105799), .A2(n109656), .B1(n105798), .B2(n109704), 
        .ZN(n85931) );
  NAND2_X1 U71548 ( .A1(n85932), .A2(n85933), .ZN(n85924) );
  AOI22_X1 U71549 ( .A1(n85266), .A2(n109680), .B1(n105796), .B2(n109674), 
        .ZN(n85933) );
  AOI22_X1 U71550 ( .A1(n105795), .A2(n109672), .B1(n105794), .B2(n109665), 
        .ZN(n85932) );
  NOR2_X1 U71551 ( .A1(n101067), .A2(n105793), .ZN(n85908) );
  AOI22_X1 U71552 ( .A1(n105099), .A2(n109674), .B1(n72739), .B2(n105174), 
        .ZN(n85906) );
  AOI22_X1 U71553 ( .A1(n105170), .A2(n109723), .B1(n85271), .B2(n109662), 
        .ZN(n85905) );
  AOI22_X1 U71554 ( .A1(n105791), .A2(n109737), .B1(n105790), .B2(n109749), 
        .ZN(n85904) );
  NAND4_X2 U71555 ( .A1(n85934), .A2(n85935), .A3(n85936), .A4(n85937), .ZN(
        n58777) );
  NOR3_X1 U71556 ( .A1(n85938), .A2(n85939), .A3(n85940), .ZN(n85937) );
  NOR2_X1 U71557 ( .A1(n102348), .A2(n105824), .ZN(n85940) );
  AOI21_X1 U71558 ( .B1(n85941), .B2(n85942), .A(n106326), .ZN(n85939) );
  NOR4_X1 U71559 ( .A1(n85943), .A2(n85944), .A3(n85945), .A4(n85946), .ZN(
        n85942) );
  OAI21_X1 U71560 ( .B1(n101171), .B2(n85224), .A(n85947), .ZN(n85946) );
  AOI22_X1 U71561 ( .A1(n105822), .A2(n109472), .B1(n105821), .B2(n109476), 
        .ZN(n85947) );
  NAND2_X1 U71562 ( .A1(n85948), .A2(n85949), .ZN(n85945) );
  AOI22_X1 U71563 ( .A1(n105820), .A2(n109504), .B1(n85231), .B2(n109485), 
        .ZN(n85949) );
  AOI22_X1 U71564 ( .A1(n105818), .A2(n109479), .B1(n85233), .B2(n72413), .ZN(
        n85948) );
  NAND2_X1 U71565 ( .A1(n85950), .A2(n85951), .ZN(n85944) );
  AOI22_X1 U71566 ( .A1(n85236), .A2(n109490), .B1(n85237), .B2(n72449), .ZN(
        n85951) );
  AOI22_X1 U71567 ( .A1(n105814), .A2(n109496), .B1(n85239), .B2(n109500), 
        .ZN(n85950) );
  NAND2_X1 U71568 ( .A1(n85952), .A2(n85953), .ZN(n85943) );
  AOI22_X1 U71569 ( .A1(n85242), .A2(n109513), .B1(n105811), .B2(n109510), 
        .ZN(n85953) );
  AOI22_X1 U71570 ( .A1(n105810), .A2(n109508), .B1(n85245), .B2(n109517), 
        .ZN(n85952) );
  NOR4_X1 U71571 ( .A1(n85954), .A2(n85955), .A3(n85956), .A4(n85957), .ZN(
        n85941) );
  OAI21_X1 U71572 ( .B1(n102357), .B2(n105808), .A(n85958), .ZN(n85957) );
  AOI22_X1 U71573 ( .A1(n105807), .A2(n109530), .B1(n72508), .B2(n105806), 
        .ZN(n85958) );
  NAND2_X1 U71574 ( .A1(n85959), .A2(n85960), .ZN(n85956) );
  AOI22_X1 U71575 ( .A1(n72381), .A2(n105804), .B1(n72488), .B2(n105803), .ZN(
        n85960) );
  AOI22_X1 U71576 ( .A1(n105802), .A2(n109526), .B1(n105801), .B2(n109518), 
        .ZN(n85959) );
  OAI21_X1 U71577 ( .B1(n102355), .B2(n105800), .A(n85961), .ZN(n85955) );
  AOI22_X1 U71578 ( .A1(n105799), .A2(n109440), .B1(n105798), .B2(n109488), 
        .ZN(n85961) );
  NAND2_X1 U71579 ( .A1(n85962), .A2(n85963), .ZN(n85954) );
  AOI22_X1 U71580 ( .A1(n85266), .A2(n109464), .B1(n105796), .B2(n109458), 
        .ZN(n85963) );
  AOI22_X1 U71581 ( .A1(n105795), .A2(n109456), .B1(n105794), .B2(n109449), 
        .ZN(n85962) );
  NOR2_X1 U71582 ( .A1(n102346), .A2(n105793), .ZN(n85938) );
  AOI22_X1 U71583 ( .A1(n105099), .A2(n109458), .B1(n72449), .B2(n105174), 
        .ZN(n85936) );
  AOI22_X1 U71584 ( .A1(n105170), .A2(n109508), .B1(n85271), .B2(n109446), 
        .ZN(n85935) );
  AOI22_X1 U71585 ( .A1(n105791), .A2(n109522), .B1(n105790), .B2(n109534), 
        .ZN(n85934) );
  NAND4_X2 U71586 ( .A1(n85964), .A2(n85965), .A3(n85966), .A4(n85967), .ZN(
        n58776) );
  NOR3_X1 U71587 ( .A1(n85968), .A2(n85969), .A3(n85970), .ZN(n85967) );
  NOR2_X1 U71588 ( .A1(n102328), .A2(n105824), .ZN(n85970) );
  AOI21_X1 U71589 ( .B1(n85971), .B2(n85972), .A(n106326), .ZN(n85969) );
  NOR4_X1 U71590 ( .A1(n85973), .A2(n85974), .A3(n85975), .A4(n85976), .ZN(
        n85972) );
  OAI21_X1 U71591 ( .B1(n101172), .B2(n85224), .A(n85977), .ZN(n85976) );
  AOI22_X1 U71592 ( .A1(n105822), .A2(n109009), .B1(n105821), .B2(n109013), 
        .ZN(n85977) );
  NAND2_X1 U71593 ( .A1(n85978), .A2(n85979), .ZN(n85975) );
  AOI22_X1 U71594 ( .A1(n105820), .A2(n109041), .B1(n85231), .B2(n109022), 
        .ZN(n85979) );
  AOI22_X1 U71595 ( .A1(n105818), .A2(n109016), .B1(n85233), .B2(n71813), .ZN(
        n85978) );
  NAND2_X1 U71596 ( .A1(n85980), .A2(n85981), .ZN(n85974) );
  AOI22_X1 U71597 ( .A1(n85236), .A2(n109027), .B1(n71849), .B2(n85237), .ZN(
        n85981) );
  AOI22_X1 U71598 ( .A1(n105814), .A2(n109033), .B1(n85239), .B2(n109037), 
        .ZN(n85980) );
  NAND2_X1 U71599 ( .A1(n85982), .A2(n85983), .ZN(n85973) );
  AOI22_X1 U71600 ( .A1(n85242), .A2(n109050), .B1(n105811), .B2(n109047), 
        .ZN(n85983) );
  AOI22_X1 U71601 ( .A1(n105810), .A2(n109045), .B1(n85245), .B2(n109054), 
        .ZN(n85982) );
  NOR4_X1 U71602 ( .A1(n85984), .A2(n85985), .A3(n85986), .A4(n85987), .ZN(
        n85971) );
  OAI21_X1 U71603 ( .B1(n102337), .B2(n105808), .A(n85988), .ZN(n85987) );
  AOI22_X1 U71604 ( .A1(n105807), .A2(n109068), .B1(n71908), .B2(n105806), 
        .ZN(n85988) );
  NAND2_X1 U71605 ( .A1(n85989), .A2(n85990), .ZN(n85986) );
  AOI22_X1 U71606 ( .A1(n71781), .A2(n105804), .B1(n71888), .B2(n105803), .ZN(
        n85990) );
  AOI22_X1 U71607 ( .A1(n105802), .A2(n109064), .B1(n105801), .B2(n109056), 
        .ZN(n85989) );
  OAI21_X1 U71608 ( .B1(n102335), .B2(n105800), .A(n85991), .ZN(n85985) );
  AOI22_X1 U71609 ( .A1(n105799), .A2(n108977), .B1(n105798), .B2(n109025), 
        .ZN(n85991) );
  NAND2_X1 U71610 ( .A1(n85992), .A2(n85993), .ZN(n85984) );
  AOI22_X1 U71611 ( .A1(n85266), .A2(n109001), .B1(n105796), .B2(n108995), 
        .ZN(n85993) );
  AOI22_X1 U71612 ( .A1(n105795), .A2(n108993), .B1(n105794), .B2(n108986), 
        .ZN(n85992) );
  NOR2_X1 U71613 ( .A1(n102326), .A2(n105793), .ZN(n85968) );
  AOI22_X1 U71614 ( .A1(n105100), .A2(n108995), .B1(n71849), .B2(n105174), 
        .ZN(n85966) );
  AOI22_X1 U71615 ( .A1(n106745), .A2(n109045), .B1(n85271), .B2(n108983), 
        .ZN(n85965) );
  AOI22_X1 U71616 ( .A1(n105791), .A2(n109060), .B1(n105790), .B2(n109072), 
        .ZN(n85964) );
  NAND4_X2 U71617 ( .A1(n85994), .A2(n85995), .A3(n85996), .A4(n85997), .ZN(
        n58775) );
  NOR3_X1 U71618 ( .A1(n85998), .A2(n85999), .A3(n86000), .ZN(n85997) );
  NOR2_X1 U71619 ( .A1(n102308), .A2(n105824), .ZN(n86000) );
  AOI21_X1 U71620 ( .B1(n86001), .B2(n86002), .A(n106326), .ZN(n85999) );
  NOR4_X1 U71621 ( .A1(n86003), .A2(n86004), .A3(n86005), .A4(n86006), .ZN(
        n86002) );
  OAI21_X1 U71622 ( .B1(n101173), .B2(n85224), .A(n86007), .ZN(n86006) );
  AOI22_X1 U71623 ( .A1(n105822), .A2(n109357), .B1(n105821), .B2(n109361), 
        .ZN(n86007) );
  NAND2_X1 U71624 ( .A1(n86008), .A2(n86009), .ZN(n86005) );
  AOI22_X1 U71625 ( .A1(n105820), .A2(n109389), .B1(n85231), .B2(n109370), 
        .ZN(n86009) );
  AOI22_X1 U71626 ( .A1(n105818), .A2(n109364), .B1(n72262), .B2(n85233), .ZN(
        n86008) );
  NAND2_X1 U71627 ( .A1(n86010), .A2(n86011), .ZN(n86004) );
  AOI22_X1 U71628 ( .A1(n85236), .A2(n109375), .B1(n72298), .B2(n85237), .ZN(
        n86011) );
  AOI22_X1 U71629 ( .A1(n105814), .A2(n109381), .B1(n85239), .B2(n109385), 
        .ZN(n86010) );
  NAND2_X1 U71630 ( .A1(n86012), .A2(n86013), .ZN(n86003) );
  AOI22_X1 U71631 ( .A1(n85242), .A2(n109398), .B1(n105811), .B2(n109395), 
        .ZN(n86013) );
  AOI22_X1 U71632 ( .A1(n105810), .A2(n109393), .B1(n85245), .B2(n109402), 
        .ZN(n86012) );
  NOR4_X1 U71633 ( .A1(n86014), .A2(n86015), .A3(n86016), .A4(n86017), .ZN(
        n86001) );
  OAI21_X1 U71634 ( .B1(n102317), .B2(n105808), .A(n86018), .ZN(n86017) );
  AOI22_X1 U71635 ( .A1(n105807), .A2(n109415), .B1(n72357), .B2(n105806), 
        .ZN(n86018) );
  NAND2_X1 U71636 ( .A1(n86019), .A2(n86020), .ZN(n86016) );
  AOI22_X1 U71637 ( .A1(n72230), .A2(n105804), .B1(n72337), .B2(n105803), .ZN(
        n86020) );
  AOI22_X1 U71638 ( .A1(n105802), .A2(n109411), .B1(n105801), .B2(n109403), 
        .ZN(n86019) );
  OAI21_X1 U71639 ( .B1(n102315), .B2(n105800), .A(n86021), .ZN(n86015) );
  AOI22_X1 U71640 ( .A1(n105799), .A2(n109325), .B1(n105798), .B2(n109373), 
        .ZN(n86021) );
  NAND2_X1 U71641 ( .A1(n86022), .A2(n86023), .ZN(n86014) );
  AOI22_X1 U71642 ( .A1(n85266), .A2(n109349), .B1(n105796), .B2(n109343), 
        .ZN(n86023) );
  AOI22_X1 U71643 ( .A1(n105795), .A2(n109341), .B1(n105794), .B2(n109334), 
        .ZN(n86022) );
  NOR2_X1 U71644 ( .A1(n102306), .A2(n105793), .ZN(n85998) );
  AOI22_X1 U71645 ( .A1(n105099), .A2(n109343), .B1(n72298), .B2(n105174), 
        .ZN(n85996) );
  AOI22_X1 U71646 ( .A1(n105170), .A2(n109393), .B1(n85271), .B2(n109331), 
        .ZN(n85995) );
  AOI22_X1 U71647 ( .A1(n105791), .A2(n109407), .B1(n105790), .B2(n109419), 
        .ZN(n85994) );
  NAND4_X2 U71648 ( .A1(n86024), .A2(n86025), .A3(n86026), .A4(n86027), .ZN(
        n58774) );
  NOR3_X1 U71649 ( .A1(n86028), .A2(n86029), .A3(n86030), .ZN(n86027) );
  NOR2_X1 U71650 ( .A1(n102288), .A2(n105824), .ZN(n86030) );
  AOI21_X1 U71651 ( .B1(n86031), .B2(n86032), .A(n106326), .ZN(n86029) );
  NOR4_X1 U71652 ( .A1(n86033), .A2(n86034), .A3(n86035), .A4(n86036), .ZN(
        n86032) );
  OAI21_X1 U71653 ( .B1(n101174), .B2(n85224), .A(n86037), .ZN(n86036) );
  AOI22_X1 U71654 ( .A1(n105822), .A2(n109239), .B1(n105821), .B2(n109243), 
        .ZN(n86037) );
  NAND2_X1 U71655 ( .A1(n86038), .A2(n86039), .ZN(n86035) );
  AOI22_X1 U71656 ( .A1(n105820), .A2(n109271), .B1(n85231), .B2(n109252), 
        .ZN(n86039) );
  AOI22_X1 U71657 ( .A1(n105818), .A2(n109246), .B1(n72111), .B2(n85233), .ZN(
        n86038) );
  NAND2_X1 U71658 ( .A1(n86040), .A2(n86041), .ZN(n86034) );
  AOI22_X1 U71659 ( .A1(n85236), .A2(n109257), .B1(n72147), .B2(n85237), .ZN(
        n86041) );
  AOI22_X1 U71660 ( .A1(n105814), .A2(n109263), .B1(n85239), .B2(n109267), 
        .ZN(n86040) );
  NAND2_X1 U71661 ( .A1(n86042), .A2(n86043), .ZN(n86033) );
  AOI22_X1 U71662 ( .A1(n72171), .A2(n105812), .B1(n105811), .B2(n109277), 
        .ZN(n86043) );
  AOI22_X1 U71663 ( .A1(n105810), .A2(n109275), .B1(n85245), .B2(n109283), 
        .ZN(n86042) );
  NOR4_X1 U71664 ( .A1(n86044), .A2(n86045), .A3(n86046), .A4(n86047), .ZN(
        n86031) );
  OAI21_X1 U71665 ( .B1(n102297), .B2(n105808), .A(n86048), .ZN(n86047) );
  AOI22_X1 U71666 ( .A1(n105807), .A2(n109296), .B1(n72206), .B2(n105806), 
        .ZN(n86048) );
  NAND2_X1 U71667 ( .A1(n86049), .A2(n86050), .ZN(n86046) );
  AOI22_X1 U71668 ( .A1(n72079), .A2(n105804), .B1(n72186), .B2(n105803), .ZN(
        n86050) );
  AOI22_X1 U71669 ( .A1(n105802), .A2(n109292), .B1(n105801), .B2(n109284), 
        .ZN(n86049) );
  OAI21_X1 U71670 ( .B1(n102295), .B2(n105800), .A(n86051), .ZN(n86045) );
  AOI22_X1 U71671 ( .A1(n105799), .A2(n109207), .B1(n105798), .B2(n109255), 
        .ZN(n86051) );
  NAND2_X1 U71672 ( .A1(n86052), .A2(n86053), .ZN(n86044) );
  AOI22_X1 U71673 ( .A1(n85266), .A2(n109231), .B1(n105796), .B2(n109225), 
        .ZN(n86053) );
  AOI22_X1 U71674 ( .A1(n105795), .A2(n109223), .B1(n105794), .B2(n109216), 
        .ZN(n86052) );
  NOR2_X1 U71675 ( .A1(n102286), .A2(n105793), .ZN(n86028) );
  AOI22_X1 U71676 ( .A1(n105101), .A2(n109225), .B1(n72147), .B2(n105174), 
        .ZN(n86026) );
  AOI22_X1 U71677 ( .A1(n105171), .A2(n109275), .B1(n85271), .B2(n109213), 
        .ZN(n86025) );
  AOI22_X1 U71678 ( .A1(n105791), .A2(n109288), .B1(n105790), .B2(n109300), 
        .ZN(n86024) );
  NAND4_X2 U71679 ( .A1(n86054), .A2(n86055), .A3(n86056), .A4(n86057), .ZN(
        n58773) );
  NOR3_X1 U71680 ( .A1(n86058), .A2(n86059), .A3(n86060), .ZN(n86057) );
  NOR2_X1 U71681 ( .A1(n102269), .A2(n105824), .ZN(n86060) );
  AOI21_X1 U71682 ( .B1(n86061), .B2(n86062), .A(n106327), .ZN(n86059) );
  NOR4_X1 U71683 ( .A1(n86063), .A2(n86064), .A3(n86065), .A4(n86066), .ZN(
        n86062) );
  OAI21_X1 U71684 ( .B1(n101175), .B2(n85224), .A(n86067), .ZN(n86066) );
  AOI22_X1 U71685 ( .A1(n105822), .A2(n109131), .B1(n105821), .B2(n109135), 
        .ZN(n86067) );
  NAND2_X1 U71686 ( .A1(n86068), .A2(n86069), .ZN(n86065) );
  AOI22_X1 U71687 ( .A1(n105820), .A2(n109162), .B1(n85231), .B2(n109144), 
        .ZN(n86069) );
  AOI22_X1 U71688 ( .A1(n105818), .A2(n109138), .B1(n85233), .B2(n71967), .ZN(
        n86068) );
  NAND2_X1 U71689 ( .A1(n86070), .A2(n86071), .ZN(n86064) );
  AOI22_X1 U71690 ( .A1(n85236), .A2(n109148), .B1(n72003), .B2(n105815), .ZN(
        n86071) );
  AOI22_X1 U71691 ( .A1(n105814), .A2(n109154), .B1(n85239), .B2(n109158), 
        .ZN(n86070) );
  NAND2_X1 U71692 ( .A1(n86072), .A2(n86073), .ZN(n86063) );
  AOI22_X1 U71693 ( .A1(n85242), .A2(n109171), .B1(n105811), .B2(n109168), 
        .ZN(n86073) );
  AOI22_X1 U71694 ( .A1(n105810), .A2(n109166), .B1(n85245), .B2(n109175), 
        .ZN(n86072) );
  NOR4_X1 U71695 ( .A1(n86074), .A2(n86075), .A3(n86076), .A4(n86077), .ZN(
        n86061) );
  OAI21_X1 U71696 ( .B1(n102278), .B2(n105808), .A(n86078), .ZN(n86077) );
  AOI22_X1 U71697 ( .A1(n105807), .A2(n109188), .B1(n72062), .B2(n105806), 
        .ZN(n86078) );
  NAND2_X1 U71698 ( .A1(n86079), .A2(n86080), .ZN(n86076) );
  AOI22_X1 U71699 ( .A1(n71935), .A2(n85256), .B1(n72042), .B2(n85257), .ZN(
        n86080) );
  AOI22_X1 U71700 ( .A1(n105802), .A2(n109184), .B1(n105801), .B2(n109176), 
        .ZN(n86079) );
  OAI21_X1 U71701 ( .B1(n102276), .B2(n105800), .A(n86081), .ZN(n86075) );
  AOI22_X1 U71702 ( .A1(n105799), .A2(n109099), .B1(n105798), .B2(n109147), 
        .ZN(n86081) );
  NAND2_X1 U71703 ( .A1(n86082), .A2(n86083), .ZN(n86074) );
  AOI22_X1 U71704 ( .A1(n85266), .A2(n109123), .B1(n105796), .B2(n109117), 
        .ZN(n86083) );
  AOI22_X1 U71705 ( .A1(n105795), .A2(n109115), .B1(n105794), .B2(n109108), 
        .ZN(n86082) );
  NOR2_X1 U71706 ( .A1(n102267), .A2(n105793), .ZN(n86058) );
  AOI22_X1 U71707 ( .A1(n105101), .A2(n109117), .B1(n72003), .B2(n105174), 
        .ZN(n86056) );
  AOI22_X1 U71708 ( .A1(n106745), .A2(n109166), .B1(n85271), .B2(n109105), 
        .ZN(n86055) );
  AOI22_X1 U71709 ( .A1(n105791), .A2(n109180), .B1(n105790), .B2(n109192), 
        .ZN(n86054) );
  NAND4_X2 U71710 ( .A1(n86084), .A2(n86085), .A3(n86086), .A4(n86087), .ZN(
        n58772) );
  NOR3_X1 U71711 ( .A1(n86088), .A2(n86089), .A3(n86090), .ZN(n86087) );
  NOR2_X1 U71712 ( .A1(n102249), .A2(n105824), .ZN(n86090) );
  AOI21_X1 U71713 ( .B1(n86091), .B2(n86092), .A(n106326), .ZN(n86089) );
  NOR4_X1 U71714 ( .A1(n86093), .A2(n86094), .A3(n86095), .A4(n86096), .ZN(
        n86092) );
  OAI21_X1 U71715 ( .B1(n101176), .B2(n85224), .A(n86097), .ZN(n86096) );
  AOI22_X1 U71716 ( .A1(n105822), .A2(n108666), .B1(n105821), .B2(n108670), 
        .ZN(n86097) );
  NAND2_X1 U71717 ( .A1(n86098), .A2(n86099), .ZN(n86095) );
  AOI22_X1 U71718 ( .A1(n105820), .A2(n108698), .B1(n85231), .B2(n108679), 
        .ZN(n86099) );
  AOI22_X1 U71719 ( .A1(n105818), .A2(n108673), .B1(n85233), .B2(n71369), .ZN(
        n86098) );
  NAND2_X1 U71720 ( .A1(n86100), .A2(n86101), .ZN(n86094) );
  AOI22_X1 U71721 ( .A1(n85236), .A2(n108684), .B1(n85237), .B2(n71405), .ZN(
        n86101) );
  AOI22_X1 U71722 ( .A1(n105814), .A2(n108690), .B1(n85239), .B2(n108694), 
        .ZN(n86100) );
  NAND2_X1 U71723 ( .A1(n86102), .A2(n86103), .ZN(n86093) );
  AOI22_X1 U71724 ( .A1(n71429), .A2(n105812), .B1(n105811), .B2(n108704), 
        .ZN(n86103) );
  AOI22_X1 U71725 ( .A1(n105810), .A2(n108702), .B1(n85245), .B2(n108710), 
        .ZN(n86102) );
  NOR4_X1 U71726 ( .A1(n86104), .A2(n86105), .A3(n86106), .A4(n86107), .ZN(
        n86091) );
  OAI21_X1 U71727 ( .B1(n102258), .B2(n105808), .A(n86108), .ZN(n86107) );
  AOI22_X1 U71728 ( .A1(n105807), .A2(n108723), .B1(n71464), .B2(n105806), 
        .ZN(n86108) );
  NAND2_X1 U71729 ( .A1(n86109), .A2(n86110), .ZN(n86106) );
  AOI22_X1 U71730 ( .A1(n71337), .A2(n85256), .B1(n71444), .B2(n85257), .ZN(
        n86110) );
  AOI22_X1 U71731 ( .A1(n105802), .A2(n108719), .B1(n105801), .B2(n108711), 
        .ZN(n86109) );
  OAI21_X1 U71732 ( .B1(n102256), .B2(n105800), .A(n86111), .ZN(n86105) );
  AOI22_X1 U71733 ( .A1(n105799), .A2(n108634), .B1(n105798), .B2(n108682), 
        .ZN(n86111) );
  NAND2_X1 U71734 ( .A1(n86112), .A2(n86113), .ZN(n86104) );
  AOI22_X1 U71735 ( .A1(n85266), .A2(n108658), .B1(n105796), .B2(n108652), 
        .ZN(n86113) );
  AOI22_X1 U71736 ( .A1(n105795), .A2(n108650), .B1(n105794), .B2(n108643), 
        .ZN(n86112) );
  NOR2_X1 U71737 ( .A1(n102247), .A2(n105793), .ZN(n86088) );
  AOI22_X1 U71738 ( .A1(n105099), .A2(n108652), .B1(n71405), .B2(n105174), 
        .ZN(n86086) );
  AOI22_X1 U71739 ( .A1(n105172), .A2(n108702), .B1(n85271), .B2(n108640), 
        .ZN(n86085) );
  AOI22_X1 U71740 ( .A1(n105791), .A2(n108715), .B1(n105790), .B2(n108727), 
        .ZN(n86084) );
  NAND4_X2 U71741 ( .A1(n86114), .A2(n86115), .A3(n86116), .A4(n86117), .ZN(
        n58771) );
  NOR3_X1 U71742 ( .A1(n86118), .A2(n86119), .A3(n86120), .ZN(n86117) );
  NOR2_X1 U71743 ( .A1(n102230), .A2(n105824), .ZN(n86120) );
  AOI21_X1 U71744 ( .B1(n86121), .B2(n86122), .A(n106327), .ZN(n86119) );
  NOR4_X1 U71745 ( .A1(n86123), .A2(n86124), .A3(n86125), .A4(n86126), .ZN(
        n86122) );
  OAI21_X1 U71746 ( .B1(n101177), .B2(n85224), .A(n86127), .ZN(n86126) );
  AOI22_X1 U71747 ( .A1(n105822), .A2(n108893), .B1(n105821), .B2(n108897), 
        .ZN(n86127) );
  NAND2_X1 U71748 ( .A1(n86128), .A2(n86129), .ZN(n86125) );
  AOI22_X1 U71749 ( .A1(n105820), .A2(n108925), .B1(n85231), .B2(n108906), 
        .ZN(n86129) );
  AOI22_X1 U71750 ( .A1(n105818), .A2(n108900), .B1(n85233), .B2(n71664), .ZN(
        n86128) );
  NAND2_X1 U71751 ( .A1(n86130), .A2(n86131), .ZN(n86124) );
  AOI22_X1 U71752 ( .A1(n85236), .A2(n108911), .B1(n71700), .B2(n85237), .ZN(
        n86131) );
  AOI22_X1 U71753 ( .A1(n105814), .A2(n108917), .B1(n85239), .B2(n108921), 
        .ZN(n86130) );
  NAND2_X1 U71754 ( .A1(n86132), .A2(n86133), .ZN(n86123) );
  AOI22_X1 U71755 ( .A1(n85242), .A2(n108934), .B1(n105811), .B2(n108931), 
        .ZN(n86133) );
  AOI22_X1 U71756 ( .A1(n105810), .A2(n108929), .B1(n85245), .B2(n108938), 
        .ZN(n86132) );
  NOR4_X1 U71757 ( .A1(n86134), .A2(n86135), .A3(n86136), .A4(n86137), .ZN(
        n86121) );
  OAI21_X1 U71758 ( .B1(n102239), .B2(n105808), .A(n86138), .ZN(n86137) );
  AOI22_X1 U71759 ( .A1(n105807), .A2(n108951), .B1(n71759), .B2(n105806), 
        .ZN(n86138) );
  NAND2_X1 U71760 ( .A1(n86139), .A2(n86140), .ZN(n86136) );
  AOI22_X1 U71761 ( .A1(n85256), .A2(n71632), .B1(n71739), .B2(n85257), .ZN(
        n86140) );
  AOI22_X1 U71762 ( .A1(n105802), .A2(n108947), .B1(n105801), .B2(n108939), 
        .ZN(n86139) );
  OAI21_X1 U71763 ( .B1(n102237), .B2(n105800), .A(n86141), .ZN(n86135) );
  AOI22_X1 U71764 ( .A1(n105799), .A2(n108861), .B1(n105798), .B2(n108909), 
        .ZN(n86141) );
  NAND2_X1 U71765 ( .A1(n86142), .A2(n86143), .ZN(n86134) );
  AOI22_X1 U71766 ( .A1(n85266), .A2(n108885), .B1(n105796), .B2(n108879), 
        .ZN(n86143) );
  AOI22_X1 U71767 ( .A1(n105795), .A2(n108877), .B1(n105794), .B2(n108870), 
        .ZN(n86142) );
  NOR2_X1 U71768 ( .A1(n102228), .A2(n105793), .ZN(n86118) );
  AOI22_X1 U71769 ( .A1(n105099), .A2(n108879), .B1(n71700), .B2(n105173), 
        .ZN(n86116) );
  AOI22_X1 U71770 ( .A1(n105171), .A2(n108929), .B1(n85271), .B2(n108867), 
        .ZN(n86115) );
  AOI22_X1 U71771 ( .A1(n105791), .A2(n108943), .B1(n105790), .B2(n108955), 
        .ZN(n86114) );
  NAND4_X2 U71772 ( .A1(n86144), .A2(n86145), .A3(n86146), .A4(n86147), .ZN(
        n58770) );
  NOR3_X1 U71773 ( .A1(n86148), .A2(n86149), .A3(n86150), .ZN(n86147) );
  NOR2_X1 U71774 ( .A1(n102210), .A2(n105824), .ZN(n86150) );
  AOI21_X1 U71775 ( .B1(n86151), .B2(n86152), .A(n106327), .ZN(n86149) );
  NOR4_X1 U71776 ( .A1(n86153), .A2(n86154), .A3(n86155), .A4(n86156), .ZN(
        n86152) );
  OAI21_X1 U71777 ( .B1(n101178), .B2(n85224), .A(n86157), .ZN(n86156) );
  AOI22_X1 U71778 ( .A1(n105822), .A2(n108781), .B1(n105821), .B2(n108785), 
        .ZN(n86157) );
  NAND2_X1 U71779 ( .A1(n86158), .A2(n86159), .ZN(n86155) );
  AOI22_X1 U71780 ( .A1(n105820), .A2(n108813), .B1(n85231), .B2(n108794), 
        .ZN(n86159) );
  AOI22_X1 U71781 ( .A1(n105818), .A2(n108788), .B1(n85233), .B2(n71520), .ZN(
        n86158) );
  NAND2_X1 U71782 ( .A1(n86160), .A2(n86161), .ZN(n86154) );
  AOI22_X1 U71783 ( .A1(n85236), .A2(n108799), .B1(n85237), .B2(n71556), .ZN(
        n86161) );
  AOI22_X1 U71784 ( .A1(n105814), .A2(n108805), .B1(n85239), .B2(n108809), 
        .ZN(n86160) );
  NAND2_X1 U71785 ( .A1(n86162), .A2(n86163), .ZN(n86153) );
  AOI22_X1 U71786 ( .A1(n105812), .A2(n108822), .B1(n105811), .B2(n108819), 
        .ZN(n86163) );
  AOI22_X1 U71787 ( .A1(n105810), .A2(n108817), .B1(n85245), .B2(n108826), 
        .ZN(n86162) );
  NOR4_X1 U71788 ( .A1(n86164), .A2(n86165), .A3(n86166), .A4(n86167), .ZN(
        n86151) );
  OAI21_X1 U71789 ( .B1(n102219), .B2(n105808), .A(n86168), .ZN(n86167) );
  AOI22_X1 U71790 ( .A1(n105807), .A2(n108839), .B1(n71615), .B2(n105806), 
        .ZN(n86168) );
  NAND2_X1 U71791 ( .A1(n86169), .A2(n86170), .ZN(n86166) );
  AOI22_X1 U71792 ( .A1(n71488), .A2(n85256), .B1(n71595), .B2(n85257), .ZN(
        n86170) );
  AOI22_X1 U71793 ( .A1(n105802), .A2(n108835), .B1(n105801), .B2(n108827), 
        .ZN(n86169) );
  OAI21_X1 U71794 ( .B1(n102217), .B2(n105800), .A(n86171), .ZN(n86165) );
  AOI22_X1 U71795 ( .A1(n105799), .A2(n108749), .B1(n105798), .B2(n108797), 
        .ZN(n86171) );
  NAND2_X1 U71796 ( .A1(n86172), .A2(n86173), .ZN(n86164) );
  AOI22_X1 U71797 ( .A1(n85266), .A2(n108773), .B1(n105796), .B2(n108767), 
        .ZN(n86173) );
  AOI22_X1 U71798 ( .A1(n105795), .A2(n108765), .B1(n105794), .B2(n108758), 
        .ZN(n86172) );
  NOR2_X1 U71799 ( .A1(n102208), .A2(n105793), .ZN(n86148) );
  AOI22_X1 U71800 ( .A1(n105100), .A2(n108767), .B1(n71556), .B2(n105174), 
        .ZN(n86146) );
  AOI22_X1 U71801 ( .A1(n105170), .A2(n108817), .B1(n85271), .B2(n108755), 
        .ZN(n86145) );
  AOI22_X1 U71802 ( .A1(n105791), .A2(n108831), .B1(n105790), .B2(n108843), 
        .ZN(n86144) );
  NAND4_X2 U71803 ( .A1(n86174), .A2(n86175), .A3(n86176), .A4(n86177), .ZN(
        n58769) );
  NOR3_X1 U71804 ( .A1(n86178), .A2(n86179), .A3(n86180), .ZN(n86177) );
  NOR2_X1 U71805 ( .A1(n102190), .A2(n105824), .ZN(n86180) );
  AOI21_X1 U71806 ( .B1(n106699), .B2(n81249), .A(n106284), .ZN(n85217) );
  NOR2_X1 U71807 ( .A1(n86181), .A2(n107027), .ZN(n80260) );
  NOR2_X1 U71808 ( .A1(n107024), .A2(n80203), .ZN(n81249) );
  AOI21_X1 U71809 ( .B1(n86182), .B2(n86183), .A(n106327), .ZN(n86179) );
  NOR4_X1 U71810 ( .A1(n86184), .A2(n86185), .A3(n86186), .A4(n86187), .ZN(
        n86183) );
  OAI21_X1 U71811 ( .B1(n101179), .B2(n85224), .A(n86188), .ZN(n86187) );
  AOI22_X1 U71812 ( .A1(n105822), .A2(n107321), .B1(n105821), .B2(n107325), 
        .ZN(n86188) );
  NOR2_X1 U71813 ( .A1(n86189), .A2(n81209), .ZN(n85227) );
  NOR2_X1 U71814 ( .A1(n86190), .A2(n107024), .ZN(n85226) );
  OR2_X1 U71815 ( .A1(n86191), .A2(n107026), .ZN(n85224) );
  NAND2_X1 U71816 ( .A1(n86192), .A2(n86193), .ZN(n86186) );
  AOI22_X1 U71817 ( .A1(n105820), .A2(n107353), .B1(n105819), .B2(n107334), 
        .ZN(n86193) );
  NOR2_X1 U71818 ( .A1(n86190), .A2(n107026), .ZN(n85231) );
  NOR2_X1 U71819 ( .A1(n86194), .A2(n81209), .ZN(n85230) );
  AOI22_X1 U71820 ( .A1(n105818), .A2(n107328), .B1(n69629), .B2(n105817), 
        .ZN(n86192) );
  NOR2_X1 U71821 ( .A1(n86190), .A2(n81208), .ZN(n85233) );
  NOR2_X1 U71822 ( .A1(n86190), .A2(n81209), .ZN(n85232) );
  NAND2_X1 U71825 ( .A1(n86196), .A2(n86197), .ZN(n86185) );
  AOI22_X1 U71826 ( .A1(n105816), .A2(n107339), .B1(n69665), .B2(n105815), 
        .ZN(n86197) );
  NOR2_X1 U71827 ( .A1(n86198), .A2(n107024), .ZN(n85237) );
  NOR2_X1 U71828 ( .A1(n86194), .A2(n81208), .ZN(n85236) );
  AOI22_X1 U71829 ( .A1(n105814), .A2(n107345), .B1(n85239), .B2(n107349), 
        .ZN(n86196) );
  NOR2_X1 U71830 ( .A1(n86198), .A2(n81209), .ZN(n85239) );
  NOR2_X1 U71831 ( .A1(n86194), .A2(n107024), .ZN(n85238) );
  NAND2_X1 U71832 ( .A1(n86199), .A2(n86200), .ZN(n86184) );
  AOI22_X1 U71833 ( .A1(n69689), .A2(n105812), .B1(n105811), .B2(n107359), 
        .ZN(n86200) );
  NOR2_X1 U71834 ( .A1(n86194), .A2(n107026), .ZN(n85243) );
  NAND2_X1 U71835 ( .A1(n86201), .A2(n105055), .ZN(n86194) );
  NOR2_X1 U71836 ( .A1(n62190), .A2(n106697), .ZN(n86201) );
  NOR2_X1 U71837 ( .A1(n86202), .A2(n104582), .ZN(n85242) );
  AOI22_X1 U71838 ( .A1(n105810), .A2(n107357), .B1(n105809), .B2(n107365), 
        .ZN(n86199) );
  NOR2_X1 U71839 ( .A1(n86202), .A2(n62190), .ZN(n85245) );
  NOR2_X1 U71840 ( .A1(n86198), .A2(n107026), .ZN(n85244) );
  NOR4_X1 U71841 ( .A1(n86203), .A2(n86204), .A3(n86205), .A4(n86206), .ZN(
        n86182) );
  OAI21_X1 U71842 ( .B1(n102199), .B2(n105808), .A(n86207), .ZN(n86206) );
  AOI22_X1 U71843 ( .A1(n105807), .A2(n107189), .B1(n69426), .B2(n105806), 
        .ZN(n86207) );
  NOR4_X1 U71844 ( .A1(n106700), .A2(n104582), .A3(n81208), .A4(n86208), .ZN(
        n85253) );
  NOR2_X1 U71845 ( .A1(n106698), .A2(n107024), .ZN(n85252) );
  NAND2_X1 U71846 ( .A1(n86209), .A2(n86210), .ZN(n85250) );
  NOR2_X1 U71847 ( .A1(n106700), .A2(n81208), .ZN(n86209) );
  NAND2_X1 U71848 ( .A1(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ), 
        .A2(n81238), .ZN(n86202) );
  NAND2_X1 U71849 ( .A1(n86211), .A2(n86212), .ZN(n86205) );
  AOI22_X1 U71850 ( .A1(n69597), .A2(n105804), .B1(n69466), .B2(n105803), .ZN(
        n86212) );
  NOR2_X1 U71851 ( .A1(n106698), .A2(n81209), .ZN(n85257) );
  NOR2_X1 U71852 ( .A1(n86191), .A2(n81208), .ZN(n85256) );
  AOI22_X1 U71853 ( .A1(n105802), .A2(n107197), .B1(n105801), .B2(n107213), 
        .ZN(n86211) );
  NOR2_X1 U71854 ( .A1(n106698), .A2(n107026), .ZN(n85259) );
  NOR2_X1 U71855 ( .A1(n86208), .A2(n62190), .ZN(n86210) );
  NOR2_X1 U71856 ( .A1(n86208), .A2(n81228), .ZN(n85258) );
  NAND2_X1 U71857 ( .A1(n106279), .A2(n62190), .ZN(n81228) );
  OAI21_X1 U71858 ( .B1(n102197), .B2(n105800), .A(n86213), .ZN(n86204) );
  AOI22_X1 U71859 ( .A1(n105799), .A2(n107289), .B1(n105798), .B2(n107337), 
        .ZN(n86213) );
  NOR2_X1 U71860 ( .A1(n86198), .A2(n81208), .ZN(n85263) );
  NAND2_X1 U71861 ( .A1(n86214), .A2(n105055), .ZN(n86198) );
  NOR2_X1 U71862 ( .A1(n104582), .A2(n106697), .ZN(n86214) );
  NOR2_X1 U71863 ( .A1(n86216), .A2(n81208), .ZN(n85262) );
  OR2_X1 U71864 ( .A1(n86216), .A2(n81209), .ZN(n85260) );
  NAND2_X1 U71865 ( .A1(n86217), .A2(n86218), .ZN(n86203) );
  AOI22_X1 U71866 ( .A1(n105797), .A2(n107313), .B1(n105796), .B2(n107307), 
        .ZN(n86218) );
  NOR2_X1 U71867 ( .A1(n86216), .A2(n107026), .ZN(n85267) );
  NOR2_X1 U71868 ( .A1(n86189), .A2(n81208), .ZN(n85266) );
  NAND2_X1 U71869 ( .A1(n86219), .A2(n86220), .ZN(n81208) );
  AOI22_X1 U71870 ( .A1(n105795), .A2(n107305), .B1(n105794), .B2(n107298), 
        .ZN(n86217) );
  NOR2_X1 U71871 ( .A1(n86191), .A2(n107024), .ZN(n85269) );
  NOR2_X1 U71872 ( .A1(n86191), .A2(n106278), .ZN(n85268) );
  NAND2_X1 U71873 ( .A1(n86219), .A2(n107025), .ZN(n81209) );
  NAND2_X1 U71874 ( .A1(n86221), .A2(n105055), .ZN(n86191) );
  NOR2_X1 U71875 ( .A1(n62190), .A2(n86215), .ZN(n86221) );
  NOR2_X1 U71876 ( .A1(n102188), .A2(n105793), .ZN(n86178) );
  AOI21_X1 U71877 ( .B1(n106699), .B2(n81198), .A(n80259), .ZN(n85270) );
  NOR2_X1 U71878 ( .A1(n86181), .A2(
        \dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .ZN(n80259) );
  OR2_X1 U71879 ( .A1(n81914), .A2(n86222), .ZN(n86181) );
  NAND2_X1 U71880 ( .A1(n59514), .A2(n106753), .ZN(n81914) );
  NOR2_X1 U71881 ( .A1(n107026), .A2(n80203), .ZN(n81198) );
  NAND2_X1 U71882 ( .A1(n86223), .A2(n86215), .ZN(n86189) );
  NOR2_X1 U71883 ( .A1(n105055), .A2(n104582), .ZN(n86223) );
  AOI22_X1 U71884 ( .A1(n105101), .A2(n107307), .B1(n69665), .B2(n106746), 
        .ZN(n86176) );
  NAND2_X1 U71885 ( .A1(n86224), .A2(n106747), .ZN(n84054) );
  NOR2_X1 U71886 ( .A1(n107027), .A2(n86222), .ZN(n86224) );
  NOR4_X1 U71887 ( .A1(n59514), .A2(
        \dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .A3(n106753), .A4(
        n86222), .ZN(n81199) );
  AOI22_X1 U71888 ( .A1(n105170), .A2(n107357), .B1(n105792), .B2(n107295), 
        .ZN(n86175) );
  OAI21_X1 U71889 ( .B1(n86216), .B2(n84053), .A(n106277), .ZN(n85271) );
  NOR4_X1 U71890 ( .A1(n59514), .A2(n106753), .A3(n107027), .A4(n86222), .ZN(
        n81250) );
  NAND2_X1 U71891 ( .A1(n81211), .A2(n106328), .ZN(n84053) );
  NAND2_X1 U71892 ( .A1(n86225), .A2(n105055), .ZN(n86216) );
  NOR2_X1 U71893 ( .A1(n86215), .A2(n104582), .ZN(n86225) );
  NAND2_X1 U71894 ( .A1(n86226), .A2(n106747), .ZN(n84095) );
  NOR2_X1 U71895 ( .A1(\dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .A2(
        n86222), .ZN(n86226) );
  AOI22_X1 U71896 ( .A1(n105791), .A2(n107205), .B1(n105790), .B2(n107181), 
        .ZN(n86174) );
  OAI21_X1 U71897 ( .B1(n81252), .B2(n86208), .A(n81253), .ZN(n85273) );
  NAND2_X1 U71898 ( .A1(n81912), .A2(n106958), .ZN(n81253) );
  NAND2_X1 U71899 ( .A1(n85208), .A2(n81211), .ZN(n81252) );
  NOR2_X1 U71900 ( .A1(n107025), .A2(n86219), .ZN(n81211) );
  OAI21_X1 U71901 ( .B1(n81254), .B2(n86208), .A(n106761), .ZN(n85272) );
  OR2_X1 U71904 ( .A1(n86215), .A2(n105055), .ZN(n86208) );
  XOR2_X1 U71905 ( .A(n81238), .B(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ), 
        .Z(n86215) );
  OAI21_X1 U71906 ( .B1(n59515), .B2(
        \dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .A(n86229), .ZN(
        n81238) );
  NOR2_X1 U71907 ( .A1(n106747), .A2(n81912), .ZN(n86229) );
  NOR2_X1 U71908 ( .A1(n86228), .A2(n107027), .ZN(n81912) );
  NAND2_X1 U71909 ( .A1(n85208), .A2(n81230), .ZN(n81254) );
  NOR2_X1 U71910 ( .A1(n86220), .A2(n86219), .ZN(n81230) );
  NOR2_X1 U71912 ( .A1(n104582), .A2(n80203), .ZN(n85208) );
  OAI21_X1 U71913 ( .B1(n80203), .B2(n86230), .A(n86231), .ZN(n58746) );
  AOI21_X1 U71914 ( .B1(n106958), .B2(n106517), .A(n105206), .ZN(n86231) );
  NAND2_X1 U71915 ( .A1(n59471), .A2(n82135), .ZN(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[1] ) );
  NOR2_X1 U71916 ( .A1(n82135), .A2(n59471), .ZN(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_0/add_38_2/carry[1] ) );
  AOI21_X1 U71917 ( .B1(IR_in[16]), .B2(n111134), .A(n111135), .ZN(n82135) );
  NAND2_X1 U71918 ( .A1(n104494), .A2(n111156), .ZN(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[1] ) );
  NOR2_X1 U71919 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [0]), 
        .A2(IR_in[8]), .ZN(n82420) );
  OR2_X1 U71921 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [28]), .A2(
        \DLX_Datapath/ArithLogUnit/A_add [28]), .ZN(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_7/RCA_1/add_38_2/carry[1] ) );
  OR2_X1 U71922 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [24]), .A2(
        \DLX_Datapath/ArithLogUnit/A_add [24]), .ZN(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_6/RCA_1/add_38_2/carry[1] ) );
  OR2_X1 U71923 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [20]), .A2(
        \DLX_Datapath/ArithLogUnit/A_add [20]), .ZN(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_5/RCA_1/add_38_2/carry[1] ) );
  NOR2_X1 U71924 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [16]), .A2(
        \DLX_Datapath/ArithLogUnit/A_add [16]), .ZN(n81846) );
  OR2_X1 U71925 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [12]), .A2(
        \DLX_Datapath/ArithLogUnit/A_add [12]), .ZN(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_3/RCA_1/add_38_2/carry[1] ) );
  OR2_X1 U71926 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [8]), .A2(
        \DLX_Datapath/ArithLogUnit/A_add [8]), .ZN(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_2/RCA_1/add_38_2/carry[1] ) );
  OR2_X1 U71927 ( .A1(\DLX_Datapath/ArithLogUnit/B_add [4]), .A2(
        \DLX_Datapath/ArithLogUnit/A_add [4]), .ZN(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[1] ) );
  NAND2_X1 U71928 ( .A1(n107620), .A2(n108858), .ZN(
        \add_1_root_DLX_Datapath/ArithLogUnit/ALU_adder/P4_SumGen/CSel_i_0/RCA_1/add_38_2/carry[1] ) );
  OAI21_X1 U71929 ( .B1(n107366), .B2(n105195), .A(n86232), .ZN(DataOut[9]) );
  AOI22_X1 U71930 ( .A1(n86233), .A2(n109761), .B1(n105788), .B2(n111075), 
        .ZN(n86232) );
  OAI21_X1 U71931 ( .B1(n107368), .B2(n106934), .A(n86235), .ZN(DataOut[8]) );
  AOI22_X1 U71932 ( .A1(n105789), .A2(n109544), .B1(n105788), .B2(n111076), 
        .ZN(n86235) );
  OAI21_X1 U71933 ( .B1(n111098), .B2(n105195), .A(n86236), .ZN(DataOut[7]) );
  AOI22_X1 U71934 ( .A1(n86233), .A2(n109084), .B1(n105788), .B2(n111088), 
        .ZN(n86236) );
  OAI21_X1 U71935 ( .B1(n111099), .B2(n106934), .A(n86237), .ZN(DataOut[6]) );
  AOI22_X1 U71936 ( .A1(n105789), .A2(n109431), .B1(n105788), .B2(n111083), 
        .ZN(n86237) );
  OAI21_X1 U71937 ( .B1(n111100), .B2(n105195), .A(n86238), .ZN(DataOut[5]) );
  AOI22_X1 U71938 ( .A1(n86233), .A2(n109312), .B1(n105788), .B2(n111077), 
        .ZN(n86238) );
  OAI21_X1 U71939 ( .B1(n111101), .B2(n106934), .A(n86239), .ZN(DataOut[4]) );
  AOI22_X1 U71940 ( .A1(n105789), .A2(n109203), .B1(n105788), .B2(n111089), 
        .ZN(n86239) );
  OAI21_X1 U71941 ( .B1(n111102), .B2(n105195), .A(n86240), .ZN(DataOut[3]) );
  AOI22_X1 U71942 ( .A1(n86233), .A2(n108739), .B1(n105788), .B2(n111084), 
        .ZN(n86240) );
  OAI21_X1 U71943 ( .B1(n107370), .B2(n106934), .A(n86241), .ZN(DataOut[31])
         );
  AOI22_X1 U71944 ( .A1(n105789), .A2(n107948), .B1(n105788), .B2(n111069), 
        .ZN(n86241) );
  OAI21_X1 U71945 ( .B1(n107372), .B2(n105195), .A(n86242), .ZN(DataOut[30])
         );
  AOI22_X1 U71946 ( .A1(n105789), .A2(n108044), .B1(n105788), .B2(n111090), 
        .ZN(n86242) );
  OAI21_X1 U71947 ( .B1(n111103), .B2(n105195), .A(n86243), .ZN(DataOut[2]) );
  AOI22_X1 U71948 ( .A1(n86233), .A2(n108965), .B1(n86234), .B2(n111085), .ZN(
        n86243) );
  OAI21_X1 U71949 ( .B1(n107374), .B2(n105195), .A(n86244), .ZN(DataOut[29])
         );
  AOI22_X1 U71950 ( .A1(n105789), .A2(n107414), .B1(n86234), .B2(n111070), 
        .ZN(n86244) );
  OAI21_X1 U71951 ( .B1(n107375), .B2(n105195), .A(n86245), .ZN(DataOut[28])
         );
  AOI22_X1 U71952 ( .A1(n86233), .A2(n107853), .B1(n86234), .B2(n111091), .ZN(
        n86245) );
  OAI21_X1 U71953 ( .B1(n107377), .B2(n105195), .A(n86246), .ZN(DataOut[27])
         );
  AOI22_X1 U71954 ( .A1(n105789), .A2(n110750), .B1(n86234), .B2(n111092), 
        .ZN(n86246) );
  OAI21_X1 U71955 ( .B1(n107379), .B2(n105195), .A(n86247), .ZN(DataOut[26])
         );
  AOI22_X1 U71956 ( .A1(n86233), .A2(n108154), .B1(n86234), .B2(n111093), .ZN(
        n86247) );
  OAI21_X1 U71957 ( .B1(n107381), .B2(n105195), .A(n86248), .ZN(DataOut[25])
         );
  AOI22_X1 U71958 ( .A1(n105789), .A2(n110851), .B1(n86234), .B2(n111094), 
        .ZN(n86248) );
  OAI21_X1 U71959 ( .B1(n107383), .B2(n105195), .A(n86249), .ZN(DataOut[24])
         );
  AOI22_X1 U71960 ( .A1(n86233), .A2(n110952), .B1(n86234), .B2(n111095), .ZN(
        n86249) );
  OAI21_X1 U71961 ( .B1(n107385), .B2(n105195), .A(n86250), .ZN(DataOut[23])
         );
  AOI22_X1 U71962 ( .A1(n105789), .A2(n110546), .B1(n86234), .B2(n111071), 
        .ZN(n86250) );
  OAI21_X1 U71963 ( .B1(n107387), .B2(n105195), .A(n86251), .ZN(DataOut[22])
         );
  AOI22_X1 U71964 ( .A1(n86233), .A2(n110332), .B1(n105788), .B2(n111066), 
        .ZN(n86251) );
  OAI21_X1 U71965 ( .B1(n107389), .B2(n105195), .A(n86252), .ZN(DataOut[21])
         );
  AOI22_X1 U71966 ( .A1(n105789), .A2(n110652), .B1(n86234), .B2(n111067), 
        .ZN(n86252) );
  OAI21_X1 U71967 ( .B1(n107391), .B2(n105195), .A(n86253), .ZN(DataOut[20])
         );
  AOI22_X1 U71968 ( .A1(n86233), .A2(n110439), .B1(n105788), .B2(n111068), 
        .ZN(n86253) );
  OAI21_X1 U71969 ( .B1(n111104), .B2(n106934), .A(n86254), .ZN(DataOut[1]) );
  AOI22_X1 U71970 ( .A1(n105789), .A2(n108854), .B1(n86234), .B2(n111086), 
        .ZN(n86254) );
  OAI21_X1 U71971 ( .B1(n107393), .B2(n106934), .A(n86255), .ZN(DataOut[19])
         );
  AOI22_X1 U71972 ( .A1(n86233), .A2(n110119), .B1(n105788), .B2(n111072), 
        .ZN(n86255) );
  OAI21_X1 U71973 ( .B1(n107395), .B2(n106934), .A(n86256), .ZN(DataOut[18])
         );
  AOI22_X1 U71974 ( .A1(n105789), .A2(n110226), .B1(n86234), .B2(n111073), 
        .ZN(n86256) );
  OAI21_X1 U71975 ( .B1(n107397), .B2(n106934), .A(n86257), .ZN(DataOut[17])
         );
  AOI22_X1 U71976 ( .A1(n105789), .A2(n110010), .B1(n105788), .B2(n111078), 
        .ZN(n86257) );
  OAI21_X1 U71977 ( .B1(n107399), .B2(n106934), .A(n86258), .ZN(DataOut[16])
         );
  AOI22_X1 U71978 ( .A1(n105789), .A2(n109895), .B1(n105788), .B2(n111074), 
        .ZN(n86258) );
  OAI21_X1 U71979 ( .B1(n107401), .B2(n106934), .A(n86259), .ZN(DataOut[15])
         );
  AOI22_X1 U71980 ( .A1(n105789), .A2(n108270), .B1(n105788), .B2(n111096), 
        .ZN(n86259) );
  OAI21_X1 U71981 ( .B1(n107403), .B2(n106934), .A(n86260), .ZN(DataOut[14])
         );
  AOI22_X1 U71982 ( .A1(n105789), .A2(n108391), .B1(n105788), .B2(n111079), 
        .ZN(n86260) );
  OAI21_X1 U71983 ( .B1(n107405), .B2(n106934), .A(n86261), .ZN(DataOut[13])
         );
  AOI22_X1 U71984 ( .A1(n105789), .A2(n108500), .B1(n105788), .B2(n111080), 
        .ZN(n86261) );
  OAI21_X1 U71985 ( .B1(n107407), .B2(n106934), .A(n86262), .ZN(DataOut[12])
         );
  AOI22_X1 U71986 ( .A1(n105789), .A2(n107741), .B1(n105788), .B2(n111097), 
        .ZN(n86262) );
  OAI21_X1 U71987 ( .B1(n107409), .B2(n106934), .A(n86263), .ZN(DataOut[11])
         );
  AOI22_X1 U71988 ( .A1(n105789), .A2(n109654), .B1(n105788), .B2(n111081), 
        .ZN(n86263) );
  OAI21_X1 U71989 ( .B1(n107411), .B2(n106934), .A(n86264), .ZN(DataOut[10])
         );
  AOI22_X1 U71990 ( .A1(n105789), .A2(n109766), .B1(n105788), .B2(n111082), 
        .ZN(n86264) );
  OAI21_X1 U71991 ( .B1(n111105), .B2(n106934), .A(n86265), .ZN(DataOut[0]) );
  AOI22_X1 U71992 ( .A1(n105789), .A2(n107415), .B1(n105788), .B2(n111087), 
        .ZN(n86265) );
  NOR2_X1 U71993 ( .A1(n86234), .A2(n86266), .ZN(n86233) );
  NOR2_X1 U71994 ( .A1(n86267), .A2(n106941), .ZN(n86234) );
  OR2_X1 U71995 ( .A1(n86268), .A2(n86269), .ZN(n86267) );
  AOI22_X1 U71996 ( .A1(n86270), .A2(n86271), .B1(n107101), .B2(n83105), .ZN(
        n86268) );
  NOR4_X1 U71997 ( .A1(n86273), .A2(n86274), .A3(n86275), .A4(n86276), .ZN(
        n86271) );
  XOR2_X1 U71998 ( .A(n100422), .B(n54618), .Z(n86276) );
  XOR2_X1 U71999 ( .A(n100423), .B(n54616), .Z(n86275) );
  XOR2_X1 U72000 ( .A(n100796), .B(n54614), .Z(n86274) );
  NOR4_X1 U72001 ( .A1(n86277), .A2(n86278), .A3(n86279), .A4(n86280), .ZN(
        n86270) );
  XOR2_X1 U72002 ( .A(n86281), .B(n86282), .Z(n86280) );
  XOR2_X1 U72003 ( .A(n107102), .B(n86283), .Z(n86279) );
  XOR2_X1 U72004 ( .A(n104723), .B(n86285), .Z(n86278) );
  XOR2_X1 U72005 ( .A(n100894), .B(n64267), .Z(n86277) );
  NOR4_X1 U72006 ( .A1(n106935), .A2(n86269), .A3(n106941), .A4(n86272), .ZN(
        n86266) );
  NAND2_X1 U72007 ( .A1(n86286), .A2(n86287), .ZN(n86272) );
  NOR4_X1 U72008 ( .A1(n86288), .A2(n86289), .A3(n86290), .A4(n86291), .ZN(
        n86287) );
  XOR2_X1 U72009 ( .A(n64267), .B(n54620), .Z(n86291) );
  XOR2_X1 U72010 ( .A(n100422), .B(n100630), .Z(n86290) );
  XOR2_X1 U72011 ( .A(n100423), .B(n100631), .Z(n86289) );
  XOR2_X1 U72012 ( .A(n100632), .B(n100796), .Z(n86288) );
  NOR3_X1 U72013 ( .A1(n86292), .A2(n86293), .A3(n86294), .ZN(n86286) );
  XOR2_X1 U72014 ( .A(n104723), .B(n86295), .Z(n86294) );
  XOR2_X1 U72015 ( .A(n86281), .B(n86296), .Z(n86293) );
  XOR2_X1 U72016 ( .A(n86297), .B(n107102), .Z(n86292) );
  NOR4_X1 U72017 ( .A1(n69323), .A2(n59326), .A3(n59325), .A4(n111022), .ZN(
        n86298) );
  XOR2_X1 U72018 ( .A(n57378), .B(n59323), .Z(n86269) );
  OAI21_X1 U72019 ( .B1(n86219), .B2(n81889), .A(n86299), .ZN(
        \DLX_Datapath/RegisterFile/next_to_transfer [1]) );
  NOR2_X1 U72020 ( .A1(n111026), .A2(n111023), .ZN(n86219) );
  OAI21_X1 U72021 ( .B1(n81889), .B2(n104582), .A(n86299), .ZN(
        \DLX_Datapath/RegisterFile/next_to_transfer [0]) );
  AOI21_X1 U72026 ( .B1(n86302), .B2(n86303), .A(n86304), .ZN(n86301) );
  OAI21_X1 U72027 ( .B1(n86305), .B2(n86306), .A(n86307), .ZN(n86304) );
  OAI21_X1 U72028 ( .B1(n86308), .B2(n86309), .A(n105786), .ZN(n86307) );
  OAI21_X1 U72029 ( .B1(n107945), .B2(n86311), .A(n86312), .ZN(n86309) );
  AOI22_X1 U72030 ( .A1(n86313), .A2(n70422), .B1(n105784), .B2(n107943), .ZN(
        n86312) );
  NAND2_X1 U72031 ( .A1(n86315), .A2(n86316), .ZN(n86308) );
  AOI22_X1 U72032 ( .A1(n86317), .A2(n107941), .B1(n86318), .B2(n107946), .ZN(
        n86316) );
  AOI22_X1 U72033 ( .A1(n86319), .A2(n107944), .B1(n86320), .B2(n107942), .ZN(
        n86315) );
  NOR4_X1 U72034 ( .A1(n86321), .A2(n86322), .A3(n86323), .A4(n86324), .ZN(
        n86305) );
  NAND2_X1 U72035 ( .A1(n86325), .A2(n86326), .ZN(n86324) );
  NOR4_X1 U72036 ( .A1(n86327), .A2(n86328), .A3(n86329), .A4(n86330), .ZN(
        n86326) );
  NAND2_X1 U72037 ( .A1(n86331), .A2(n86332), .ZN(n86330) );
  AOI22_X1 U72038 ( .A1(n86333), .A2(n107922), .B1(n86334), .B2(n107923), .ZN(
        n86332) );
  AOI22_X1 U72039 ( .A1(n86335), .A2(n107931), .B1(n86336), .B2(n107929), .ZN(
        n86331) );
  NAND2_X1 U72040 ( .A1(n86337), .A2(n86338), .ZN(n86329) );
  AOI22_X1 U72041 ( .A1(n86339), .A2(n70291), .B1(n86340), .B2(n107926), .ZN(
        n86338) );
  AOI22_X1 U72042 ( .A1(n86341), .A2(n70395), .B1(n86342), .B2(n107855), .ZN(
        n86337) );
  NAND2_X1 U72043 ( .A1(n86343), .A2(n86344), .ZN(n86328) );
  AOI22_X1 U72044 ( .A1(n86345), .A2(n107859), .B1(n105770), .B2(n70295), .ZN(
        n86344) );
  AOI22_X1 U72045 ( .A1(n86347), .A2(n107927), .B1(n86348), .B2(n107924), .ZN(
        n86343) );
  NAND2_X1 U72046 ( .A1(n86349), .A2(n86350), .ZN(n86327) );
  AOI22_X1 U72047 ( .A1(n86351), .A2(n107857), .B1(n86352), .B2(n107861), .ZN(
        n86350) );
  AOI22_X1 U72048 ( .A1(n86353), .A2(n107860), .B1(n86354), .B2(n70297), .ZN(
        n86349) );
  NOR4_X1 U72049 ( .A1(n86355), .A2(n86356), .A3(n86357), .A4(n86358), .ZN(
        n86325) );
  NAND2_X1 U72050 ( .A1(n86359), .A2(n86360), .ZN(n86358) );
  AOI22_X1 U72051 ( .A1(n86361), .A2(n107932), .B1(n86362), .B2(n107935), .ZN(
        n86360) );
  AOI22_X1 U72052 ( .A1(n105761), .A2(n107936), .B1(n105760), .B2(n107938), 
        .ZN(n86359) );
  NAND2_X1 U72053 ( .A1(n86365), .A2(n86366), .ZN(n86357) );
  AOI22_X1 U72054 ( .A1(n86367), .A2(n107937), .B1(n105758), .B2(n107933), 
        .ZN(n86366) );
  AOI22_X1 U72055 ( .A1(n86369), .A2(n107939), .B1(n86370), .B2(n107934), .ZN(
        n86365) );
  NAND2_X1 U72056 ( .A1(n86371), .A2(n86372), .ZN(n86356) );
  AOI22_X1 U72057 ( .A1(n86373), .A2(n70405), .B1(n86374), .B2(n70404), .ZN(
        n86372) );
  AOI22_X1 U72058 ( .A1(n86375), .A2(n70407), .B1(n86376), .B2(n107940), .ZN(
        n86371) );
  NAND2_X1 U72059 ( .A1(n86377), .A2(n86378), .ZN(n86355) );
  AOI22_X1 U72060 ( .A1(n86379), .A2(n107925), .B1(n86380), .B2(n107930), .ZN(
        n86378) );
  AOI22_X1 U72061 ( .A1(n86381), .A2(n70402), .B1(n105748), .B2(n107928), .ZN(
        n86377) );
  NAND2_X1 U72062 ( .A1(n86383), .A2(n86384), .ZN(n86323) );
  NOR4_X1 U72063 ( .A1(n86385), .A2(n86386), .A3(n86387), .A4(n86388), .ZN(
        n86384) );
  NAND2_X1 U72064 ( .A1(n86389), .A2(n86390), .ZN(n86388) );
  AOI22_X1 U72065 ( .A1(n86391), .A2(n107869), .B1(n86392), .B2(n107871), .ZN(
        n86390) );
  AOI22_X1 U72066 ( .A1(n86393), .A2(n70320), .B1(n86394), .B2(n107870), .ZN(
        n86389) );
  NAND2_X1 U72067 ( .A1(n86395), .A2(n86396), .ZN(n86387) );
  AOI22_X1 U72068 ( .A1(n86397), .A2(n70324), .B1(n86398), .B2(n70326), .ZN(
        n86396) );
  AOI22_X1 U72069 ( .A1(n86399), .A2(n107875), .B1(n105740), .B2(n107876), 
        .ZN(n86395) );
  NAND2_X1 U72070 ( .A1(n86401), .A2(n86402), .ZN(n86386) );
  AOI22_X1 U72071 ( .A1(n105739), .A2(n107873), .B1(n86404), .B2(n70321), .ZN(
        n86402) );
  AOI22_X1 U72072 ( .A1(n86405), .A2(n107877), .B1(n105736), .B2(n107874), 
        .ZN(n86401) );
  NAND2_X1 U72073 ( .A1(n86407), .A2(n86408), .ZN(n86385) );
  AOI22_X1 U72074 ( .A1(n86409), .A2(n107881), .B1(n86410), .B2(n70331), .ZN(
        n86408) );
  AOI22_X1 U72075 ( .A1(n105733), .A2(n107880), .B1(n86412), .B2(n70329), .ZN(
        n86407) );
  NOR4_X1 U72076 ( .A1(n86413), .A2(n86414), .A3(n86415), .A4(n86416), .ZN(
        n86383) );
  NAND2_X1 U72077 ( .A1(n86417), .A2(n86418), .ZN(n86416) );
  AOI22_X1 U72078 ( .A1(n86419), .A2(n107864), .B1(n86420), .B2(n107856), .ZN(
        n86418) );
  AOI22_X1 U72079 ( .A1(n86421), .A2(n107858), .B1(n86422), .B2(n70303), .ZN(
        n86417) );
  NAND2_X1 U72080 ( .A1(n86423), .A2(n86424), .ZN(n86415) );
  AOI22_X1 U72081 ( .A1(n86425), .A2(n107863), .B1(n105726), .B2(n107866), 
        .ZN(n86424) );
  AOI22_X1 U72082 ( .A1(n105725), .A2(n107868), .B1(n105724), .B2(n107865), 
        .ZN(n86423) );
  NAND2_X1 U72083 ( .A1(n86429), .A2(n86430), .ZN(n86414) );
  AOI22_X1 U72084 ( .A1(n86431), .A2(n70312), .B1(n86432), .B2(n107862), .ZN(
        n86430) );
  AOI22_X1 U72085 ( .A1(n86433), .A2(n70304), .B1(n86434), .B2(n70308), .ZN(
        n86429) );
  NAND2_X1 U72086 ( .A1(n86435), .A2(n86436), .ZN(n86413) );
  AOI22_X1 U72087 ( .A1(n86437), .A2(n70317), .B1(n86438), .B2(n70316), .ZN(
        n86436) );
  AOI22_X1 U72088 ( .A1(n86439), .A2(n70314), .B1(n105716), .B2(n107872), .ZN(
        n86435) );
  NAND2_X1 U72089 ( .A1(n86441), .A2(n86442), .ZN(n86322) );
  NOR4_X1 U72090 ( .A1(n86443), .A2(n86444), .A3(n86445), .A4(n86446), .ZN(
        n86442) );
  NAND2_X1 U72091 ( .A1(n86447), .A2(n86448), .ZN(n86446) );
  AOI22_X1 U72092 ( .A1(n86449), .A2(n70354), .B1(n105714), .B2(n107890), .ZN(
        n86448) );
  AOI22_X1 U72093 ( .A1(n86451), .A2(n107893), .B1(n86452), .B2(n70350), .ZN(
        n86447) );
  NAND2_X1 U72094 ( .A1(n86453), .A2(n86454), .ZN(n86445) );
  AOI22_X1 U72095 ( .A1(n105711), .A2(n107897), .B1(n86456), .B2(n107896), 
        .ZN(n86454) );
  AOI22_X1 U72096 ( .A1(n105709), .A2(n107889), .B1(n105708), .B2(n107891), 
        .ZN(n86453) );
  NAND2_X1 U72097 ( .A1(n86459), .A2(n86460), .ZN(n86444) );
  AOI22_X1 U72098 ( .A1(n86461), .A2(n107898), .B1(n86462), .B2(n107895), .ZN(
        n86460) );
  AOI22_X1 U72099 ( .A1(n86463), .A2(n70358), .B1(n86464), .B2(n70360), .ZN(
        n86459) );
  NAND2_X1 U72100 ( .A1(n86465), .A2(n86466), .ZN(n86443) );
  AOI22_X1 U72101 ( .A1(n105703), .A2(n70363), .B1(n86468), .B2(n70366), .ZN(
        n86466) );
  AOI22_X1 U72102 ( .A1(n86469), .A2(n107894), .B1(n86470), .B2(n70355), .ZN(
        n86465) );
  NOR4_X1 U72103 ( .A1(n86471), .A2(n86472), .A3(n86473), .A4(n86474), .ZN(
        n86441) );
  NAND2_X1 U72104 ( .A1(n86475), .A2(n86476), .ZN(n86474) );
  AOI22_X1 U72105 ( .A1(n86477), .A2(n70330), .B1(n86478), .B2(n107884), .ZN(
        n86476) );
  AOI22_X1 U72106 ( .A1(n105697), .A2(n107879), .B1(n86480), .B2(n70334), .ZN(
        n86475) );
  NAND2_X1 U72107 ( .A1(n86481), .A2(n86482), .ZN(n86473) );
  AOI22_X1 U72108 ( .A1(n86483), .A2(n70343), .B1(n105694), .B2(n107886), .ZN(
        n86482) );
  AOI22_X1 U72109 ( .A1(n86485), .A2(n107887), .B1(n86486), .B2(n107878), .ZN(
        n86481) );
  NAND2_X1 U72110 ( .A1(n86487), .A2(n86488), .ZN(n86472) );
  AOI22_X1 U72111 ( .A1(n86489), .A2(n107885), .B1(n105690), .B2(n70342), .ZN(
        n86488) );
  AOI22_X1 U72112 ( .A1(n86491), .A2(n107883), .B1(n86492), .B2(n107888), .ZN(
        n86487) );
  NAND2_X1 U72113 ( .A1(n86493), .A2(n86494), .ZN(n86471) );
  AOI22_X1 U72114 ( .A1(n105687), .A2(n70348), .B1(n86496), .B2(n107892), .ZN(
        n86494) );
  AOI22_X1 U72115 ( .A1(n86497), .A2(n70346), .B1(n86498), .B2(n107882), .ZN(
        n86493) );
  NAND2_X1 U72116 ( .A1(n86499), .A2(n86500), .ZN(n86321) );
  NOR4_X1 U72117 ( .A1(n86501), .A2(n86502), .A3(n86503), .A4(n86504), .ZN(
        n86500) );
  NAND2_X1 U72118 ( .A1(n86505), .A2(n86506), .ZN(n86504) );
  AOI22_X1 U72119 ( .A1(n86507), .A2(n107914), .B1(n86508), .B2(n107913), .ZN(
        n86506) );
  AOI22_X1 U72120 ( .A1(n86509), .A2(n70382), .B1(n86510), .B2(n107911), .ZN(
        n86505) );
  NAND2_X1 U72121 ( .A1(n86511), .A2(n86512), .ZN(n86503) );
  AOI22_X1 U72122 ( .A1(n86513), .A2(n107909), .B1(n105678), .B2(n107912), 
        .ZN(n86512) );
  AOI22_X1 U72123 ( .A1(n86515), .A2(n70388), .B1(n105677), .B2(n107910), .ZN(
        n86511) );
  NAND2_X1 U72124 ( .A1(n86517), .A2(n86518), .ZN(n86502) );
  AOI22_X1 U72125 ( .A1(n86519), .A2(n107919), .B1(n86520), .B2(n70394), .ZN(
        n86518) );
  AOI22_X1 U72126 ( .A1(n86521), .A2(n107917), .B1(n86522), .B2(n107918), .ZN(
        n86517) );
  NAND2_X1 U72127 ( .A1(n86523), .A2(n86524), .ZN(n86501) );
  AOI22_X1 U72128 ( .A1(n86525), .A2(n70386), .B1(n86526), .B2(n107916), .ZN(
        n86524) );
  AOI22_X1 U72129 ( .A1(n86527), .A2(n107920), .B1(n86528), .B2(n107915), .ZN(
        n86523) );
  NOR4_X1 U72130 ( .A1(n86529), .A2(n86530), .A3(n86531), .A4(n86532), .ZN(
        n86499) );
  NAND2_X1 U72131 ( .A1(n86533), .A2(n86534), .ZN(n86532) );
  AOI22_X1 U72132 ( .A1(n105675), .A2(n107900), .B1(n86536), .B2(n107901), 
        .ZN(n86534) );
  AOI22_X1 U72133 ( .A1(n86537), .A2(n70367), .B1(n86538), .B2(n70365), .ZN(
        n86533) );
  NAND2_X1 U72134 ( .A1(n86539), .A2(n86540), .ZN(n86531) );
  AOI22_X1 U72135 ( .A1(n86541), .A2(n107906), .B1(n86542), .B2(n107899), .ZN(
        n86540) );
  AOI22_X1 U72136 ( .A1(n86543), .A2(n70364), .B1(n105668), .B2(n107903), .ZN(
        n86539) );
  NAND2_X1 U72137 ( .A1(n86545), .A2(n86546), .ZN(n86530) );
  AOI22_X1 U72138 ( .A1(n86547), .A2(n107902), .B1(n86548), .B2(n107907), .ZN(
        n86546) );
  AOI22_X1 U72139 ( .A1(n105665), .A2(n107908), .B1(n86550), .B2(n107905), 
        .ZN(n86545) );
  NAND2_X1 U72140 ( .A1(n86551), .A2(n86552), .ZN(n86529) );
  AOI22_X1 U72141 ( .A1(n86553), .A2(n70383), .B1(n86554), .B2(n70369), .ZN(
        n86552) );
  AOI22_X1 U72142 ( .A1(n105661), .A2(n70372), .B1(n86556), .B2(n70376), .ZN(
        n86551) );
  AOI21_X1 U72143 ( .B1(n86302), .B2(n86558), .A(n86559), .ZN(n86557) );
  OAI21_X1 U72144 ( .B1(n86560), .B2(n86306), .A(n86561), .ZN(n86559) );
  OAI21_X1 U72145 ( .B1(n86562), .B2(n86563), .A(n105786), .ZN(n86561) );
  OAI21_X1 U72146 ( .B1(n108041), .B2(n86311), .A(n86564), .ZN(n86563) );
  AOI22_X1 U72147 ( .A1(n86313), .A2(n70564), .B1(n105784), .B2(n108039), .ZN(
        n86564) );
  NAND2_X1 U72148 ( .A1(n86565), .A2(n86566), .ZN(n86562) );
  AOI22_X1 U72149 ( .A1(n86317), .A2(n108037), .B1(n86318), .B2(n108042), .ZN(
        n86566) );
  AOI22_X1 U72150 ( .A1(n86319), .A2(n108040), .B1(n86320), .B2(n108038), .ZN(
        n86565) );
  NOR4_X1 U72151 ( .A1(n86567), .A2(n86568), .A3(n86569), .A4(n86570), .ZN(
        n86560) );
  NAND2_X1 U72152 ( .A1(n86571), .A2(n86572), .ZN(n86570) );
  NOR4_X1 U72153 ( .A1(n86573), .A2(n86574), .A3(n86575), .A4(n86576), .ZN(
        n86572) );
  NAND2_X1 U72154 ( .A1(n86577), .A2(n86578), .ZN(n86576) );
  AOI22_X1 U72155 ( .A1(n86333), .A2(n108018), .B1(n86334), .B2(n108019), .ZN(
        n86578) );
  AOI22_X1 U72156 ( .A1(n86335), .A2(n108027), .B1(n86336), .B2(n108025), .ZN(
        n86577) );
  NAND2_X1 U72157 ( .A1(n86579), .A2(n86580), .ZN(n86575) );
  AOI22_X1 U72158 ( .A1(n86339), .A2(n70433), .B1(n86340), .B2(n108022), .ZN(
        n86580) );
  AOI22_X1 U72159 ( .A1(n86341), .A2(n70537), .B1(n86342), .B2(n107952), .ZN(
        n86579) );
  NAND2_X1 U72160 ( .A1(n86581), .A2(n86582), .ZN(n86574) );
  AOI22_X1 U72161 ( .A1(n86345), .A2(n107956), .B1(n105770), .B2(n70437), .ZN(
        n86582) );
  AOI22_X1 U72162 ( .A1(n86347), .A2(n108023), .B1(n86348), .B2(n108020), .ZN(
        n86581) );
  NAND2_X1 U72163 ( .A1(n86583), .A2(n86584), .ZN(n86573) );
  AOI22_X1 U72164 ( .A1(n86351), .A2(n107954), .B1(n86352), .B2(n107958), .ZN(
        n86584) );
  AOI22_X1 U72165 ( .A1(n86353), .A2(n107957), .B1(n86354), .B2(n70439), .ZN(
        n86583) );
  NOR4_X1 U72166 ( .A1(n86585), .A2(n86586), .A3(n86587), .A4(n86588), .ZN(
        n86571) );
  NAND2_X1 U72167 ( .A1(n86589), .A2(n86590), .ZN(n86588) );
  AOI22_X1 U72168 ( .A1(n86361), .A2(n108028), .B1(n86362), .B2(n108031), .ZN(
        n86590) );
  AOI22_X1 U72169 ( .A1(n105761), .A2(n108032), .B1(n105760), .B2(n108034), 
        .ZN(n86589) );
  NAND2_X1 U72170 ( .A1(n86591), .A2(n86592), .ZN(n86587) );
  AOI22_X1 U72171 ( .A1(n86367), .A2(n108033), .B1(n105758), .B2(n108029), 
        .ZN(n86592) );
  AOI22_X1 U72172 ( .A1(n86369), .A2(n108035), .B1(n86370), .B2(n108030), .ZN(
        n86591) );
  NAND2_X1 U72173 ( .A1(n86593), .A2(n86594), .ZN(n86586) );
  AOI22_X1 U72174 ( .A1(n86373), .A2(n70547), .B1(n86374), .B2(n70546), .ZN(
        n86594) );
  AOI22_X1 U72175 ( .A1(n86375), .A2(n70549), .B1(n86376), .B2(n108036), .ZN(
        n86593) );
  NAND2_X1 U72176 ( .A1(n86595), .A2(n86596), .ZN(n86585) );
  AOI22_X1 U72177 ( .A1(n86379), .A2(n108021), .B1(n86380), .B2(n108026), .ZN(
        n86596) );
  AOI22_X1 U72178 ( .A1(n86381), .A2(n70544), .B1(n105748), .B2(n108024), .ZN(
        n86595) );
  NAND2_X1 U72179 ( .A1(n86597), .A2(n86598), .ZN(n86569) );
  NOR4_X1 U72180 ( .A1(n86599), .A2(n86600), .A3(n86601), .A4(n86602), .ZN(
        n86598) );
  NAND2_X1 U72181 ( .A1(n86603), .A2(n86604), .ZN(n86602) );
  AOI22_X1 U72182 ( .A1(n86391), .A2(n107966), .B1(n86392), .B2(n107968), .ZN(
        n86604) );
  AOI22_X1 U72183 ( .A1(n86393), .A2(n70462), .B1(n86394), .B2(n107967), .ZN(
        n86603) );
  NAND2_X1 U72184 ( .A1(n86605), .A2(n86606), .ZN(n86601) );
  AOI22_X1 U72185 ( .A1(n86397), .A2(n70466), .B1(n86398), .B2(n70468), .ZN(
        n86606) );
  AOI22_X1 U72186 ( .A1(n86399), .A2(n107972), .B1(n105740), .B2(n107973), 
        .ZN(n86605) );
  NAND2_X1 U72187 ( .A1(n86607), .A2(n86608), .ZN(n86600) );
  AOI22_X1 U72188 ( .A1(n105739), .A2(n107971), .B1(n86404), .B2(n70463), .ZN(
        n86608) );
  AOI22_X1 U72189 ( .A1(n86405), .A2(n107974), .B1(n105736), .B2(n70461), .ZN(
        n86607) );
  NAND2_X1 U72190 ( .A1(n86609), .A2(n86610), .ZN(n86599) );
  AOI22_X1 U72191 ( .A1(n86409), .A2(n107976), .B1(n86410), .B2(n70473), .ZN(
        n86610) );
  AOI22_X1 U72192 ( .A1(n105733), .A2(n70474), .B1(n86412), .B2(n70471), .ZN(
        n86609) );
  NOR4_X1 U72193 ( .A1(n86611), .A2(n86612), .A3(n86613), .A4(n86614), .ZN(
        n86597) );
  NAND2_X1 U72194 ( .A1(n86615), .A2(n86616), .ZN(n86614) );
  AOI22_X1 U72195 ( .A1(n86419), .A2(n107961), .B1(n86420), .B2(n107953), .ZN(
        n86616) );
  AOI22_X1 U72196 ( .A1(n86421), .A2(n107955), .B1(n86422), .B2(n70445), .ZN(
        n86615) );
  NAND2_X1 U72197 ( .A1(n86617), .A2(n86618), .ZN(n86613) );
  AOI22_X1 U72198 ( .A1(n86425), .A2(n107960), .B1(n105726), .B2(n107963), 
        .ZN(n86618) );
  AOI22_X1 U72199 ( .A1(n105725), .A2(n107965), .B1(n105724), .B2(n107962), 
        .ZN(n86617) );
  NAND2_X1 U72200 ( .A1(n86619), .A2(n86620), .ZN(n86612) );
  AOI22_X1 U72201 ( .A1(n86431), .A2(n70454), .B1(n86432), .B2(n107959), .ZN(
        n86620) );
  AOI22_X1 U72202 ( .A1(n86433), .A2(n70446), .B1(n86434), .B2(n70450), .ZN(
        n86619) );
  NAND2_X1 U72203 ( .A1(n86621), .A2(n86622), .ZN(n86611) );
  AOI22_X1 U72204 ( .A1(n86437), .A2(n107970), .B1(n86438), .B2(n70458), .ZN(
        n86622) );
  AOI22_X1 U72205 ( .A1(n86439), .A2(n70456), .B1(n105716), .B2(n107969), .ZN(
        n86621) );
  NAND2_X1 U72206 ( .A1(n86623), .A2(n86624), .ZN(n86568) );
  NOR4_X1 U72207 ( .A1(n86625), .A2(n86626), .A3(n86627), .A4(n86628), .ZN(
        n86624) );
  NAND2_X1 U72208 ( .A1(n86629), .A2(n86630), .ZN(n86628) );
  AOI22_X1 U72209 ( .A1(n86449), .A2(n70496), .B1(n105714), .B2(n107985), .ZN(
        n86630) );
  AOI22_X1 U72210 ( .A1(n86451), .A2(n107988), .B1(n86452), .B2(n70492), .ZN(
        n86629) );
  NAND2_X1 U72211 ( .A1(n86631), .A2(n86632), .ZN(n86627) );
  AOI22_X1 U72212 ( .A1(n105711), .A2(n107991), .B1(n86456), .B2(n107990), 
        .ZN(n86632) );
  AOI22_X1 U72213 ( .A1(n105709), .A2(n107984), .B1(n105708), .B2(n107986), 
        .ZN(n86631) );
  NAND2_X1 U72214 ( .A1(n86633), .A2(n86634), .ZN(n86626) );
  AOI22_X1 U72215 ( .A1(n86461), .A2(n107992), .B1(n86462), .B2(n107989), .ZN(
        n86634) );
  AOI22_X1 U72216 ( .A1(n86463), .A2(n70500), .B1(n86464), .B2(n70502), .ZN(
        n86633) );
  NAND2_X1 U72217 ( .A1(n86635), .A2(n86636), .ZN(n86625) );
  AOI22_X1 U72218 ( .A1(n105703), .A2(n107995), .B1(n86468), .B2(n70508), .ZN(
        n86636) );
  AOI22_X1 U72219 ( .A1(n86469), .A2(n70494), .B1(n86470), .B2(n70497), .ZN(
        n86635) );
  NOR4_X1 U72220 ( .A1(n86637), .A2(n86638), .A3(n86639), .A4(n86640), .ZN(
        n86623) );
  NAND2_X1 U72221 ( .A1(n86641), .A2(n86642), .ZN(n86640) );
  AOI22_X1 U72222 ( .A1(n86477), .A2(n70472), .B1(n86478), .B2(n107979), .ZN(
        n86642) );
  AOI22_X1 U72223 ( .A1(n105697), .A2(n70470), .B1(n86480), .B2(n70476), .ZN(
        n86641) );
  NAND2_X1 U72224 ( .A1(n86643), .A2(n86644), .ZN(n86639) );
  AOI22_X1 U72225 ( .A1(n86483), .A2(n70485), .B1(n105694), .B2(n107981), .ZN(
        n86644) );
  AOI22_X1 U72226 ( .A1(n86485), .A2(n107982), .B1(n86486), .B2(n107975), .ZN(
        n86643) );
  NAND2_X1 U72227 ( .A1(n86645), .A2(n86646), .ZN(n86638) );
  AOI22_X1 U72228 ( .A1(n86489), .A2(n107980), .B1(n105690), .B2(n70484), .ZN(
        n86646) );
  AOI22_X1 U72229 ( .A1(n86491), .A2(n107978), .B1(n86492), .B2(n107983), .ZN(
        n86645) );
  NAND2_X1 U72230 ( .A1(n86647), .A2(n86648), .ZN(n86637) );
  AOI22_X1 U72231 ( .A1(n105687), .A2(n70490), .B1(n86496), .B2(n107987), .ZN(
        n86648) );
  AOI22_X1 U72232 ( .A1(n86497), .A2(n70488), .B1(n86498), .B2(n107977), .ZN(
        n86647) );
  NAND2_X1 U72233 ( .A1(n86649), .A2(n86650), .ZN(n86567) );
  NOR4_X1 U72234 ( .A1(n86651), .A2(n86652), .A3(n86653), .A4(n86654), .ZN(
        n86650) );
  NAND2_X1 U72235 ( .A1(n86655), .A2(n86656), .ZN(n86654) );
  AOI22_X1 U72236 ( .A1(n86507), .A2(n108010), .B1(n86508), .B2(n108009), .ZN(
        n86656) );
  AOI22_X1 U72237 ( .A1(n86509), .A2(n70524), .B1(n86510), .B2(n108007), .ZN(
        n86655) );
  NAND2_X1 U72238 ( .A1(n86657), .A2(n86658), .ZN(n86653) );
  AOI22_X1 U72239 ( .A1(n86513), .A2(n108005), .B1(n105678), .B2(n108008), 
        .ZN(n86658) );
  AOI22_X1 U72240 ( .A1(n86515), .A2(n70530), .B1(n105677), .B2(n108006), .ZN(
        n86657) );
  NAND2_X1 U72241 ( .A1(n86659), .A2(n86660), .ZN(n86652) );
  AOI22_X1 U72242 ( .A1(n86519), .A2(n108016), .B1(n86520), .B2(n70536), .ZN(
        n86660) );
  AOI22_X1 U72243 ( .A1(n86521), .A2(n108014), .B1(n86522), .B2(n108015), .ZN(
        n86659) );
  NAND2_X1 U72244 ( .A1(n86661), .A2(n86662), .ZN(n86651) );
  AOI22_X1 U72245 ( .A1(n86525), .A2(n108011), .B1(n86526), .B2(n108013), .ZN(
        n86662) );
  AOI22_X1 U72246 ( .A1(n86527), .A2(n70535), .B1(n86528), .B2(n108012), .ZN(
        n86661) );
  NOR4_X1 U72247 ( .A1(n86663), .A2(n86664), .A3(n86665), .A4(n86666), .ZN(
        n86649) );
  NAND2_X1 U72248 ( .A1(n86667), .A2(n86668), .ZN(n86666) );
  AOI22_X1 U72249 ( .A1(n105675), .A2(n107994), .B1(n86536), .B2(n107997), 
        .ZN(n86668) );
  AOI22_X1 U72250 ( .A1(n86537), .A2(n107996), .B1(n86538), .B2(n70507), .ZN(
        n86667) );
  NAND2_X1 U72251 ( .A1(n86669), .A2(n86670), .ZN(n86665) );
  AOI22_X1 U72252 ( .A1(n86541), .A2(n108002), .B1(n86542), .B2(n107993), .ZN(
        n86670) );
  AOI22_X1 U72253 ( .A1(n86543), .A2(n70506), .B1(n105668), .B2(n107999), .ZN(
        n86669) );
  NAND2_X1 U72254 ( .A1(n86671), .A2(n86672), .ZN(n86664) );
  AOI22_X1 U72255 ( .A1(n86547), .A2(n107998), .B1(n86548), .B2(n108003), .ZN(
        n86672) );
  AOI22_X1 U72256 ( .A1(n105665), .A2(n108004), .B1(n86550), .B2(n108001), 
        .ZN(n86671) );
  NAND2_X1 U72257 ( .A1(n86673), .A2(n86674), .ZN(n86663) );
  AOI22_X1 U72258 ( .A1(n86553), .A2(n70525), .B1(n86554), .B2(n70511), .ZN(
        n86674) );
  AOI22_X1 U72259 ( .A1(n105661), .A2(n70514), .B1(n86556), .B2(n70518), .ZN(
        n86673) );
  AOI21_X1 U72260 ( .B1(n86302), .B2(n86676), .A(n86677), .ZN(n86675) );
  OAI21_X1 U72261 ( .B1(n86678), .B2(n86306), .A(n86679), .ZN(n86677) );
  OAI21_X1 U72262 ( .B1(n86680), .B2(n86681), .A(n105786), .ZN(n86679) );
  OAI21_X1 U72263 ( .B1(n107166), .B2(n86311), .A(n86682), .ZN(n86681) );
  AOI22_X1 U72264 ( .A1(n86313), .A2(n69429), .B1(n105784), .B2(n107170), .ZN(
        n86682) );
  NAND2_X1 U72265 ( .A1(n86683), .A2(n86684), .ZN(n86680) );
  AOI22_X1 U72266 ( .A1(n86317), .A2(n107174), .B1(n86318), .B2(n106838), .ZN(
        n86684) );
  AOI22_X1 U72267 ( .A1(n86319), .A2(n107168), .B1(n86320), .B2(n107172), .ZN(
        n86683) );
  NOR4_X1 U72268 ( .A1(n86685), .A2(n86686), .A3(n86687), .A4(n86688), .ZN(
        n86678) );
  NAND2_X1 U72269 ( .A1(n86689), .A2(n86690), .ZN(n86688) );
  NOR4_X1 U72270 ( .A1(n86691), .A2(n86692), .A3(n86693), .A4(n86694), .ZN(
        n86690) );
  NAND2_X1 U72271 ( .A1(n86695), .A2(n86696), .ZN(n86694) );
  AOI22_X1 U72272 ( .A1(n86333), .A2(n107212), .B1(n86334), .B2(n107210), .ZN(
        n86696) );
  AOI22_X1 U72273 ( .A1(n86335), .A2(n107194), .B1(n86336), .B2(n107198), .ZN(
        n86695) );
  NAND2_X1 U72274 ( .A1(n86697), .A2(n86698), .ZN(n86693) );
  AOI22_X1 U72275 ( .A1(n86339), .A2(n69486), .B1(n86340), .B2(n107204), .ZN(
        n86698) );
  AOI22_X1 U72276 ( .A1(n86341), .A2(n69483), .B1(n86342), .B2(n107214), .ZN(
        n86697) );
  NAND2_X1 U72277 ( .A1(n86699), .A2(n86700), .ZN(n86692) );
  AOI22_X1 U72278 ( .A1(n86345), .A2(n107218), .B1(n105770), .B2(n69490), .ZN(
        n86700) );
  AOI22_X1 U72279 ( .A1(n86347), .A2(n107202), .B1(n86348), .B2(n107208), .ZN(
        n86699) );
  NAND2_X1 U72280 ( .A1(n86701), .A2(n86702), .ZN(n86691) );
  AOI22_X1 U72281 ( .A1(n86351), .A2(n107216), .B1(n86352), .B2(n107220), .ZN(
        n86702) );
  AOI22_X1 U72282 ( .A1(n86353), .A2(n107219), .B1(n86354), .B2(n69492), .ZN(
        n86701) );
  NOR4_X1 U72283 ( .A1(n86703), .A2(n86704), .A3(n86705), .A4(n86706), .ZN(
        n86689) );
  NAND2_X1 U72284 ( .A1(n86707), .A2(n86708), .ZN(n86706) );
  AOI22_X1 U72285 ( .A1(n86361), .A2(n107192), .B1(n86362), .B2(n107186), .ZN(
        n86708) );
  AOI22_X1 U72286 ( .A1(n105761), .A2(n107184), .B1(n105760), .B2(n107180), 
        .ZN(n86707) );
  NAND2_X1 U72287 ( .A1(n86709), .A2(n86710), .ZN(n86705) );
  AOI22_X1 U72288 ( .A1(n86367), .A2(n107182), .B1(n105758), .B2(n107190), 
        .ZN(n86710) );
  AOI22_X1 U72289 ( .A1(n86369), .A2(n107178), .B1(n86370), .B2(n107188), .ZN(
        n86709) );
  NAND2_X1 U72290 ( .A1(n86711), .A2(n86712), .ZN(n86704) );
  AOI22_X1 U72291 ( .A1(n86373), .A2(n69463), .B1(n86374), .B2(n69465), .ZN(
        n86712) );
  AOI22_X1 U72292 ( .A1(n86375), .A2(n69459), .B1(n86376), .B2(n107176), .ZN(
        n86711) );
  NAND2_X1 U72293 ( .A1(n86713), .A2(n86714), .ZN(n86703) );
  AOI22_X1 U72294 ( .A1(n86379), .A2(n107206), .B1(n86380), .B2(n107196), .ZN(
        n86714) );
  AOI22_X1 U72295 ( .A1(n86381), .A2(n69469), .B1(n105748), .B2(n107200), .ZN(
        n86713) );
  NAND2_X1 U72296 ( .A1(n86715), .A2(n86716), .ZN(n86687) );
  NOR4_X1 U72297 ( .A1(n86717), .A2(n86718), .A3(n86719), .A4(n86720), .ZN(
        n86716) );
  NAND2_X1 U72298 ( .A1(n86721), .A2(n86722), .ZN(n86720) );
  AOI22_X1 U72299 ( .A1(n86391), .A2(n107229), .B1(n86392), .B2(n107231), .ZN(
        n86722) );
  AOI22_X1 U72300 ( .A1(n86393), .A2(n69515), .B1(n86394), .B2(n107230), .ZN(
        n86721) );
  NAND2_X1 U72301 ( .A1(n86723), .A2(n86724), .ZN(n86719) );
  AOI22_X1 U72302 ( .A1(n86397), .A2(n69519), .B1(n86398), .B2(n69521), .ZN(
        n86724) );
  AOI22_X1 U72303 ( .A1(n86399), .A2(n107236), .B1(n105740), .B2(n107237), 
        .ZN(n86723) );
  NAND2_X1 U72304 ( .A1(n86725), .A2(n86726), .ZN(n86718) );
  AOI22_X1 U72305 ( .A1(n105739), .A2(n107234), .B1(n86404), .B2(n107235), 
        .ZN(n86726) );
  AOI22_X1 U72306 ( .A1(n86405), .A2(n107238), .B1(n105736), .B2(n69514), .ZN(
        n86725) );
  NAND2_X1 U72307 ( .A1(n86727), .A2(n86728), .ZN(n86717) );
  AOI22_X1 U72308 ( .A1(n86409), .A2(n107243), .B1(n86410), .B2(n69526), .ZN(
        n86728) );
  AOI22_X1 U72309 ( .A1(n105733), .A2(n107242), .B1(n86412), .B2(n69524), .ZN(
        n86727) );
  NOR4_X1 U72310 ( .A1(n86729), .A2(n86730), .A3(n86731), .A4(n86732), .ZN(
        n86715) );
  NAND2_X1 U72311 ( .A1(n86733), .A2(n86734), .ZN(n86732) );
  AOI22_X1 U72312 ( .A1(n86419), .A2(n107224), .B1(n86420), .B2(n107215), .ZN(
        n86734) );
  AOI22_X1 U72313 ( .A1(n86421), .A2(n107217), .B1(n86422), .B2(n69498), .ZN(
        n86733) );
  NAND2_X1 U72314 ( .A1(n86735), .A2(n86736), .ZN(n86731) );
  AOI22_X1 U72315 ( .A1(n86425), .A2(n107222), .B1(n105726), .B2(n107226), 
        .ZN(n86736) );
  AOI22_X1 U72316 ( .A1(n105725), .A2(n107228), .B1(n105724), .B2(n107225), 
        .ZN(n86735) );
  NAND2_X1 U72317 ( .A1(n86737), .A2(n86738), .ZN(n86730) );
  AOI22_X1 U72318 ( .A1(n86431), .A2(n69507), .B1(n86432), .B2(n107221), .ZN(
        n86738) );
  AOI22_X1 U72319 ( .A1(n86433), .A2(n107223), .B1(n86434), .B2(n69503), .ZN(
        n86737) );
  NAND2_X1 U72320 ( .A1(n86739), .A2(n86740), .ZN(n86729) );
  AOI22_X1 U72321 ( .A1(n86437), .A2(n107233), .B1(n86438), .B2(n69511), .ZN(
        n86740) );
  AOI22_X1 U72322 ( .A1(n86439), .A2(n69509), .B1(n105716), .B2(n107232), .ZN(
        n86739) );
  NAND2_X1 U72323 ( .A1(n86741), .A2(n86742), .ZN(n86686) );
  NOR4_X1 U72324 ( .A1(n86743), .A2(n86744), .A3(n86745), .A4(n86746), .ZN(
        n86742) );
  NAND2_X1 U72325 ( .A1(n86747), .A2(n86748), .ZN(n86746) );
  AOI22_X1 U72326 ( .A1(n86449), .A2(n69549), .B1(n105714), .B2(n107253), .ZN(
        n86748) );
  AOI22_X1 U72327 ( .A1(n86451), .A2(n107256), .B1(n86452), .B2(n69545), .ZN(
        n86747) );
  NAND2_X1 U72328 ( .A1(n86749), .A2(n86750), .ZN(n86745) );
  AOI22_X1 U72329 ( .A1(n105711), .A2(n107261), .B1(n86456), .B2(n107260), 
        .ZN(n86750) );
  AOI22_X1 U72330 ( .A1(n105709), .A2(n107252), .B1(n105708), .B2(n107254), 
        .ZN(n86749) );
  NAND2_X1 U72331 ( .A1(n86751), .A2(n86752), .ZN(n86744) );
  AOI22_X1 U72332 ( .A1(n86461), .A2(n107262), .B1(n86462), .B2(n107258), .ZN(
        n86752) );
  AOI22_X1 U72333 ( .A1(n86463), .A2(n69553), .B1(n86464), .B2(n69555), .ZN(
        n86751) );
  NAND2_X1 U72334 ( .A1(n86753), .A2(n86754), .ZN(n86743) );
  AOI22_X1 U72335 ( .A1(n105703), .A2(n107265), .B1(n86468), .B2(n69561), .ZN(
        n86754) );
  AOI22_X1 U72336 ( .A1(n86469), .A2(n107257), .B1(n86470), .B2(n107259), .ZN(
        n86753) );
  NOR4_X1 U72337 ( .A1(n86755), .A2(n86756), .A3(n86757), .A4(n86758), .ZN(
        n86741) );
  NAND2_X1 U72338 ( .A1(n86759), .A2(n86760), .ZN(n86758) );
  AOI22_X1 U72339 ( .A1(n86477), .A2(n107241), .B1(n86478), .B2(n107246), .ZN(
        n86760) );
  AOI22_X1 U72340 ( .A1(n105697), .A2(n107240), .B1(n86480), .B2(n69529), .ZN(
        n86759) );
  NAND2_X1 U72341 ( .A1(n86761), .A2(n86762), .ZN(n86757) );
  AOI22_X1 U72342 ( .A1(n86483), .A2(n69538), .B1(n105694), .B2(n107248), .ZN(
        n86762) );
  AOI22_X1 U72343 ( .A1(n86485), .A2(n107249), .B1(n86486), .B2(n107239), .ZN(
        n86761) );
  NAND2_X1 U72344 ( .A1(n86763), .A2(n86764), .ZN(n86756) );
  AOI22_X1 U72345 ( .A1(n86489), .A2(n107247), .B1(n105690), .B2(n107251), 
        .ZN(n86764) );
  AOI22_X1 U72346 ( .A1(n86491), .A2(n107245), .B1(n86492), .B2(n107250), .ZN(
        n86763) );
  NAND2_X1 U72347 ( .A1(n86765), .A2(n86766), .ZN(n86755) );
  AOI22_X1 U72348 ( .A1(n105687), .A2(n69543), .B1(n86496), .B2(n107255), .ZN(
        n86766) );
  AOI22_X1 U72349 ( .A1(n86497), .A2(n69541), .B1(n86498), .B2(n107244), .ZN(
        n86765) );
  NAND2_X1 U72350 ( .A1(n86767), .A2(n86768), .ZN(n86685) );
  NOR4_X1 U72351 ( .A1(n86769), .A2(n86770), .A3(n86771), .A4(n86772), .ZN(
        n86768) );
  NAND2_X1 U72352 ( .A1(n86773), .A2(n86774), .ZN(n86772) );
  AOI22_X1 U72353 ( .A1(n86507), .A2(n107281), .B1(n86508), .B2(n107280), .ZN(
        n86774) );
  AOI22_X1 U72354 ( .A1(n86509), .A2(n69577), .B1(n86510), .B2(n107278), .ZN(
        n86773) );
  NAND2_X1 U72355 ( .A1(n86775), .A2(n86776), .ZN(n86771) );
  AOI22_X1 U72356 ( .A1(n86513), .A2(n107276), .B1(n105678), .B2(n107279), 
        .ZN(n86776) );
  AOI22_X1 U72357 ( .A1(n86515), .A2(n69583), .B1(n105677), .B2(n107277), .ZN(
        n86775) );
  NAND2_X1 U72358 ( .A1(n86777), .A2(n86778), .ZN(n86770) );
  AOI22_X1 U72359 ( .A1(n86519), .A2(n107286), .B1(n86520), .B2(n69589), .ZN(
        n86778) );
  AOI22_X1 U72360 ( .A1(n86521), .A2(n107284), .B1(n86522), .B2(n107285), .ZN(
        n86777) );
  NAND2_X1 U72361 ( .A1(n86779), .A2(n86780), .ZN(n86769) );
  AOI22_X1 U72362 ( .A1(n86525), .A2(n69581), .B1(n86526), .B2(n107283), .ZN(
        n86780) );
  AOI22_X1 U72363 ( .A1(n86527), .A2(n69588), .B1(n86528), .B2(n107282), .ZN(
        n86779) );
  NOR4_X1 U72364 ( .A1(n86781), .A2(n86782), .A3(n86783), .A4(n86784), .ZN(
        n86767) );
  NAND2_X1 U72365 ( .A1(n86785), .A2(n86786), .ZN(n86784) );
  AOI22_X1 U72366 ( .A1(n105675), .A2(n107264), .B1(n86536), .B2(n107268), 
        .ZN(n86786) );
  AOI22_X1 U72367 ( .A1(n86537), .A2(n107267), .B1(n86538), .B2(n69560), .ZN(
        n86785) );
  NAND2_X1 U72368 ( .A1(n86787), .A2(n86788), .ZN(n86783) );
  AOI22_X1 U72369 ( .A1(n86541), .A2(n107273), .B1(n86542), .B2(n107263), .ZN(
        n86788) );
  AOI22_X1 U72370 ( .A1(n86543), .A2(n107266), .B1(n105668), .B2(n107270), 
        .ZN(n86787) );
  NAND2_X1 U72371 ( .A1(n86789), .A2(n86790), .ZN(n86782) );
  AOI22_X1 U72372 ( .A1(n86547), .A2(n107269), .B1(n86548), .B2(n107274), .ZN(
        n86790) );
  AOI22_X1 U72373 ( .A1(n105665), .A2(n107275), .B1(n86550), .B2(n107272), 
        .ZN(n86789) );
  NAND2_X1 U72374 ( .A1(n86791), .A2(n86792), .ZN(n86781) );
  AOI22_X1 U72375 ( .A1(n86553), .A2(n69578), .B1(n86554), .B2(n69564), .ZN(
        n86792) );
  AOI22_X1 U72376 ( .A1(n105661), .A2(n69567), .B1(n86556), .B2(n69571), .ZN(
        n86791) );
  AOI21_X1 U72377 ( .B1(n86302), .B2(n86794), .A(n86795), .ZN(n86793) );
  OAI21_X1 U72378 ( .B1(n86796), .B2(n86306), .A(n86797), .ZN(n86795) );
  OAI21_X1 U72379 ( .B1(n86798), .B2(n86799), .A(n105786), .ZN(n86797) );
  OAI21_X1 U72380 ( .B1(n107850), .B2(n86311), .A(n86800), .ZN(n86799) );
  AOI22_X1 U72381 ( .A1(n86313), .A2(n70278), .B1(n105784), .B2(n107848), .ZN(
        n86800) );
  NAND2_X1 U72382 ( .A1(n86801), .A2(n86802), .ZN(n86798) );
  AOI22_X1 U72383 ( .A1(n86317), .A2(n107846), .B1(n86318), .B2(n107851), .ZN(
        n86802) );
  AOI22_X1 U72384 ( .A1(n86319), .A2(n107849), .B1(n86320), .B2(n107847), .ZN(
        n86801) );
  NOR4_X1 U72385 ( .A1(n86803), .A2(n86804), .A3(n86805), .A4(n86806), .ZN(
        n86796) );
  NAND2_X1 U72386 ( .A1(n86807), .A2(n86808), .ZN(n86806) );
  NOR4_X1 U72387 ( .A1(n86809), .A2(n86810), .A3(n86811), .A4(n86812), .ZN(
        n86808) );
  NAND2_X1 U72388 ( .A1(n86813), .A2(n86814), .ZN(n86812) );
  AOI22_X1 U72389 ( .A1(n86333), .A2(n107826), .B1(n86334), .B2(n107827), .ZN(
        n86814) );
  AOI22_X1 U72390 ( .A1(n86335), .A2(n107836), .B1(n86336), .B2(n107834), .ZN(
        n86813) );
  NAND2_X1 U72391 ( .A1(n86815), .A2(n86816), .ZN(n86811) );
  AOI22_X1 U72392 ( .A1(n86339), .A2(n70147), .B1(n86340), .B2(n107830), .ZN(
        n86816) );
  AOI22_X1 U72393 ( .A1(n86341), .A2(n70251), .B1(n86342), .B2(n107752), .ZN(
        n86815) );
  NAND2_X1 U72394 ( .A1(n86817), .A2(n86818), .ZN(n86810) );
  AOI22_X1 U72395 ( .A1(n86345), .A2(n107756), .B1(n105770), .B2(n70151), .ZN(
        n86818) );
  AOI22_X1 U72396 ( .A1(n86347), .A2(n107831), .B1(n86348), .B2(n107828), .ZN(
        n86817) );
  NAND2_X1 U72397 ( .A1(n86819), .A2(n86820), .ZN(n86809) );
  AOI22_X1 U72398 ( .A1(n86351), .A2(n107754), .B1(n86352), .B2(n107758), .ZN(
        n86820) );
  AOI22_X1 U72399 ( .A1(n86353), .A2(n107757), .B1(n86354), .B2(n70153), .ZN(
        n86819) );
  NOR4_X1 U72400 ( .A1(n86821), .A2(n86822), .A3(n86823), .A4(n86824), .ZN(
        n86807) );
  NAND2_X1 U72401 ( .A1(n86825), .A2(n86826), .ZN(n86824) );
  AOI22_X1 U72402 ( .A1(n86361), .A2(n107837), .B1(n86362), .B2(n107840), .ZN(
        n86826) );
  AOI22_X1 U72403 ( .A1(n105761), .A2(n107841), .B1(n105760), .B2(n107843), 
        .ZN(n86825) );
  NAND2_X1 U72404 ( .A1(n86827), .A2(n86828), .ZN(n86823) );
  AOI22_X1 U72405 ( .A1(n86367), .A2(n107842), .B1(n105758), .B2(n107838), 
        .ZN(n86828) );
  AOI22_X1 U72406 ( .A1(n86369), .A2(n107844), .B1(n86370), .B2(n107839), .ZN(
        n86827) );
  NAND2_X1 U72407 ( .A1(n86829), .A2(n86830), .ZN(n86822) );
  AOI22_X1 U72408 ( .A1(n86373), .A2(n70261), .B1(n86374), .B2(n70260), .ZN(
        n86830) );
  AOI22_X1 U72409 ( .A1(n86375), .A2(n70263), .B1(n86376), .B2(n107845), .ZN(
        n86829) );
  NAND2_X1 U72410 ( .A1(n86831), .A2(n86832), .ZN(n86821) );
  AOI22_X1 U72411 ( .A1(n86379), .A2(n107829), .B1(n86380), .B2(n107835), .ZN(
        n86832) );
  AOI22_X1 U72412 ( .A1(n86381), .A2(n70258), .B1(n105748), .B2(n107833), .ZN(
        n86831) );
  NAND2_X1 U72413 ( .A1(n86833), .A2(n86834), .ZN(n86805) );
  NOR4_X1 U72414 ( .A1(n86835), .A2(n86836), .A3(n86837), .A4(n86838), .ZN(
        n86834) );
  NAND2_X1 U72415 ( .A1(n86839), .A2(n86840), .ZN(n86838) );
  AOI22_X1 U72416 ( .A1(n86391), .A2(n107767), .B1(n86392), .B2(n107769), .ZN(
        n86840) );
  AOI22_X1 U72417 ( .A1(n86393), .A2(n70176), .B1(n86394), .B2(n107768), .ZN(
        n86839) );
  NAND2_X1 U72418 ( .A1(n86841), .A2(n86842), .ZN(n86837) );
  AOI22_X1 U72419 ( .A1(n86397), .A2(n70180), .B1(n86398), .B2(n70182), .ZN(
        n86842) );
  AOI22_X1 U72420 ( .A1(n86399), .A2(n107775), .B1(n105740), .B2(n107776), 
        .ZN(n86841) );
  NAND2_X1 U72421 ( .A1(n86843), .A2(n86844), .ZN(n86836) );
  AOI22_X1 U72422 ( .A1(n105739), .A2(n107772), .B1(n86404), .B2(n107774), 
        .ZN(n86844) );
  AOI22_X1 U72423 ( .A1(n86405), .A2(n107777), .B1(n105736), .B2(n107773), 
        .ZN(n86843) );
  NAND2_X1 U72424 ( .A1(n86845), .A2(n86846), .ZN(n86835) );
  AOI22_X1 U72425 ( .A1(n86409), .A2(n107782), .B1(n86410), .B2(n70187), .ZN(
        n86846) );
  AOI22_X1 U72426 ( .A1(n105733), .A2(n107781), .B1(n86412), .B2(n70185), .ZN(
        n86845) );
  NOR4_X1 U72427 ( .A1(n86847), .A2(n86848), .A3(n86849), .A4(n86850), .ZN(
        n86833) );
  NAND2_X1 U72428 ( .A1(n86851), .A2(n86852), .ZN(n86850) );
  AOI22_X1 U72429 ( .A1(n86419), .A2(n107762), .B1(n86420), .B2(n107753), .ZN(
        n86852) );
  AOI22_X1 U72430 ( .A1(n86421), .A2(n107755), .B1(n86422), .B2(n70159), .ZN(
        n86851) );
  NAND2_X1 U72431 ( .A1(n86853), .A2(n86854), .ZN(n86849) );
  AOI22_X1 U72432 ( .A1(n86425), .A2(n107760), .B1(n105726), .B2(n107764), 
        .ZN(n86854) );
  AOI22_X1 U72433 ( .A1(n105725), .A2(n107766), .B1(n105724), .B2(n107763), 
        .ZN(n86853) );
  NAND2_X1 U72434 ( .A1(n86855), .A2(n86856), .ZN(n86848) );
  AOI22_X1 U72435 ( .A1(n86431), .A2(n70168), .B1(n86432), .B2(n107759), .ZN(
        n86856) );
  AOI22_X1 U72436 ( .A1(n86433), .A2(n107761), .B1(n86434), .B2(n107765), .ZN(
        n86855) );
  NAND2_X1 U72437 ( .A1(n86857), .A2(n86858), .ZN(n86847) );
  AOI22_X1 U72438 ( .A1(n86437), .A2(n107771), .B1(n86438), .B2(n70172), .ZN(
        n86858) );
  AOI22_X1 U72439 ( .A1(n86439), .A2(n70170), .B1(n105716), .B2(n107770), .ZN(
        n86857) );
  NAND2_X1 U72440 ( .A1(n86859), .A2(n86860), .ZN(n86804) );
  NOR4_X1 U72441 ( .A1(n86861), .A2(n86862), .A3(n86863), .A4(n86864), .ZN(
        n86860) );
  NAND2_X1 U72442 ( .A1(n86865), .A2(n86866), .ZN(n86864) );
  AOI22_X1 U72443 ( .A1(n86449), .A2(n70210), .B1(n105714), .B2(n107792), .ZN(
        n86866) );
  AOI22_X1 U72444 ( .A1(n86451), .A2(n107795), .B1(n86452), .B2(n70206), .ZN(
        n86865) );
  NAND2_X1 U72445 ( .A1(n86867), .A2(n86868), .ZN(n86863) );
  AOI22_X1 U72446 ( .A1(n105711), .A2(n107798), .B1(n86456), .B2(n107797), 
        .ZN(n86868) );
  AOI22_X1 U72447 ( .A1(n105709), .A2(n107791), .B1(n105708), .B2(n107793), 
        .ZN(n86867) );
  NAND2_X1 U72448 ( .A1(n86869), .A2(n86870), .ZN(n86862) );
  AOI22_X1 U72449 ( .A1(n86461), .A2(n107799), .B1(n86462), .B2(n70209), .ZN(
        n86870) );
  AOI22_X1 U72450 ( .A1(n86463), .A2(n70214), .B1(n86464), .B2(n70216), .ZN(
        n86869) );
  NAND2_X1 U72451 ( .A1(n86871), .A2(n86872), .ZN(n86861) );
  AOI22_X1 U72452 ( .A1(n105703), .A2(n107802), .B1(n86468), .B2(n70222), .ZN(
        n86872) );
  AOI22_X1 U72453 ( .A1(n86469), .A2(n70208), .B1(n86470), .B2(n107796), .ZN(
        n86871) );
  NOR4_X1 U72454 ( .A1(n86873), .A2(n86874), .A3(n86875), .A4(n86876), .ZN(
        n86859) );
  NAND2_X1 U72455 ( .A1(n86877), .A2(n86878), .ZN(n86876) );
  AOI22_X1 U72456 ( .A1(n86477), .A2(n107780), .B1(n86478), .B2(n107785), .ZN(
        n86878) );
  AOI22_X1 U72457 ( .A1(n105697), .A2(n107779), .B1(n86480), .B2(n70190), .ZN(
        n86877) );
  NAND2_X1 U72458 ( .A1(n86879), .A2(n86880), .ZN(n86875) );
  AOI22_X1 U72459 ( .A1(n86483), .A2(n70199), .B1(n105694), .B2(n107787), .ZN(
        n86880) );
  AOI22_X1 U72460 ( .A1(n86485), .A2(n107788), .B1(n86486), .B2(n107778), .ZN(
        n86879) );
  NAND2_X1 U72461 ( .A1(n86881), .A2(n86882), .ZN(n86874) );
  AOI22_X1 U72462 ( .A1(n86489), .A2(n107786), .B1(n105690), .B2(n107790), 
        .ZN(n86882) );
  AOI22_X1 U72463 ( .A1(n86491), .A2(n107784), .B1(n86492), .B2(n107789), .ZN(
        n86881) );
  NAND2_X1 U72464 ( .A1(n86883), .A2(n86884), .ZN(n86873) );
  AOI22_X1 U72465 ( .A1(n105687), .A2(n70204), .B1(n86496), .B2(n107794), .ZN(
        n86884) );
  AOI22_X1 U72466 ( .A1(n86497), .A2(n70202), .B1(n86498), .B2(n107783), .ZN(
        n86883) );
  NAND2_X1 U72467 ( .A1(n86885), .A2(n86886), .ZN(n86803) );
  NOR4_X1 U72468 ( .A1(n86887), .A2(n86888), .A3(n86889), .A4(n86890), .ZN(
        n86886) );
  NAND2_X1 U72469 ( .A1(n86891), .A2(n86892), .ZN(n86890) );
  AOI22_X1 U72470 ( .A1(n86507), .A2(n107819), .B1(n86508), .B2(n107818), .ZN(
        n86892) );
  AOI22_X1 U72471 ( .A1(n86509), .A2(n70238), .B1(n86510), .B2(n107816), .ZN(
        n86891) );
  NAND2_X1 U72472 ( .A1(n86893), .A2(n86894), .ZN(n86889) );
  AOI22_X1 U72473 ( .A1(n86513), .A2(n107814), .B1(n105678), .B2(n107817), 
        .ZN(n86894) );
  AOI22_X1 U72474 ( .A1(n86515), .A2(n70244), .B1(n105677), .B2(n107815), .ZN(
        n86893) );
  NAND2_X1 U72475 ( .A1(n86895), .A2(n86896), .ZN(n86888) );
  AOI22_X1 U72476 ( .A1(n86519), .A2(n107824), .B1(n86520), .B2(n70250), .ZN(
        n86896) );
  AOI22_X1 U72477 ( .A1(n86521), .A2(n107822), .B1(n86522), .B2(n107823), .ZN(
        n86895) );
  NAND2_X1 U72478 ( .A1(n86897), .A2(n86898), .ZN(n86887) );
  AOI22_X1 U72479 ( .A1(n86525), .A2(n70242), .B1(n86526), .B2(n107821), .ZN(
        n86898) );
  AOI22_X1 U72480 ( .A1(n86527), .A2(n70249), .B1(n86528), .B2(n107820), .ZN(
        n86897) );
  NOR4_X1 U72481 ( .A1(n86899), .A2(n86900), .A3(n86901), .A4(n86902), .ZN(
        n86885) );
  NAND2_X1 U72482 ( .A1(n86903), .A2(n86904), .ZN(n86902) );
  AOI22_X1 U72483 ( .A1(n105675), .A2(n107801), .B1(n86536), .B2(n107805), 
        .ZN(n86904) );
  AOI22_X1 U72484 ( .A1(n86537), .A2(n107804), .B1(n86538), .B2(n70221), .ZN(
        n86903) );
  NAND2_X1 U72485 ( .A1(n86905), .A2(n86906), .ZN(n86901) );
  AOI22_X1 U72486 ( .A1(n86541), .A2(n107810), .B1(n86542), .B2(n107800), .ZN(
        n86906) );
  AOI22_X1 U72487 ( .A1(n86543), .A2(n107803), .B1(n105668), .B2(n107807), 
        .ZN(n86905) );
  NAND2_X1 U72488 ( .A1(n86907), .A2(n86908), .ZN(n86900) );
  AOI22_X1 U72489 ( .A1(n86547), .A2(n107806), .B1(n86548), .B2(n107811), .ZN(
        n86908) );
  AOI22_X1 U72490 ( .A1(n105665), .A2(n107813), .B1(n86550), .B2(n107809), 
        .ZN(n86907) );
  NAND2_X1 U72491 ( .A1(n86909), .A2(n86910), .ZN(n86899) );
  AOI22_X1 U72492 ( .A1(n86553), .A2(n70239), .B1(n86554), .B2(n70225), .ZN(
        n86910) );
  AOI22_X1 U72493 ( .A1(n105661), .A2(n70228), .B1(n86556), .B2(n107812), .ZN(
        n86909) );
  AOI21_X1 U72494 ( .B1(n86302), .B2(n86912), .A(n86913), .ZN(n86911) );
  OAI21_X1 U72495 ( .B1(n86914), .B2(n86306), .A(n86915), .ZN(n86913) );
  OAI21_X1 U72496 ( .B1(n86916), .B2(n86917), .A(n105786), .ZN(n86915) );
  OAI21_X1 U72497 ( .B1(n110745), .B2(n86311), .A(n86918), .ZN(n86917) );
  AOI22_X1 U72498 ( .A1(n86313), .A2(n74124), .B1(n105784), .B2(n110743), .ZN(
        n86918) );
  NAND2_X1 U72499 ( .A1(n86919), .A2(n86920), .ZN(n86916) );
  AOI22_X1 U72500 ( .A1(n86317), .A2(n110741), .B1(n86318), .B2(n110746), .ZN(
        n86920) );
  AOI22_X1 U72501 ( .A1(n86319), .A2(n110744), .B1(n86320), .B2(n110742), .ZN(
        n86919) );
  NOR4_X1 U72502 ( .A1(n86921), .A2(n86922), .A3(n86923), .A4(n86924), .ZN(
        n86914) );
  NAND2_X1 U72503 ( .A1(n86925), .A2(n86926), .ZN(n86924) );
  NOR4_X1 U72504 ( .A1(n86927), .A2(n86928), .A3(n86929), .A4(n86930), .ZN(
        n86926) );
  NAND2_X1 U72505 ( .A1(n86931), .A2(n86932), .ZN(n86930) );
  AOI22_X1 U72506 ( .A1(n86333), .A2(n110722), .B1(n86334), .B2(n110723), .ZN(
        n86932) );
  AOI22_X1 U72507 ( .A1(n86335), .A2(n110731), .B1(n86336), .B2(n110729), .ZN(
        n86931) );
  NAND2_X1 U72508 ( .A1(n86933), .A2(n86934), .ZN(n86929) );
  AOI22_X1 U72509 ( .A1(n86339), .A2(n73993), .B1(n86340), .B2(n110726), .ZN(
        n86934) );
  AOI22_X1 U72510 ( .A1(n86341), .A2(n74097), .B1(n86342), .B2(n110655), .ZN(
        n86933) );
  NAND2_X1 U72511 ( .A1(n86935), .A2(n86936), .ZN(n86928) );
  AOI22_X1 U72512 ( .A1(n86345), .A2(n110659), .B1(n105770), .B2(n73997), .ZN(
        n86936) );
  AOI22_X1 U72513 ( .A1(n86347), .A2(n110727), .B1(n86348), .B2(n110724), .ZN(
        n86935) );
  NAND2_X1 U72514 ( .A1(n86937), .A2(n86938), .ZN(n86927) );
  AOI22_X1 U72515 ( .A1(n86351), .A2(n110657), .B1(n86352), .B2(n110661), .ZN(
        n86938) );
  AOI22_X1 U72516 ( .A1(n86353), .A2(n110660), .B1(n86354), .B2(n73999), .ZN(
        n86937) );
  NOR4_X1 U72517 ( .A1(n86939), .A2(n86940), .A3(n86941), .A4(n86942), .ZN(
        n86925) );
  NAND2_X1 U72518 ( .A1(n86943), .A2(n86944), .ZN(n86942) );
  AOI22_X1 U72519 ( .A1(n86361), .A2(n110732), .B1(n86362), .B2(n110735), .ZN(
        n86944) );
  AOI22_X1 U72520 ( .A1(n105761), .A2(n110736), .B1(n105760), .B2(n110738), 
        .ZN(n86943) );
  NAND2_X1 U72521 ( .A1(n86945), .A2(n86946), .ZN(n86941) );
  AOI22_X1 U72522 ( .A1(n86367), .A2(n110737), .B1(n105758), .B2(n110733), 
        .ZN(n86946) );
  AOI22_X1 U72523 ( .A1(n86369), .A2(n110739), .B1(n86370), .B2(n110734), .ZN(
        n86945) );
  NAND2_X1 U72524 ( .A1(n86947), .A2(n86948), .ZN(n86940) );
  AOI22_X1 U72525 ( .A1(n86373), .A2(n74107), .B1(n86374), .B2(n74106), .ZN(
        n86948) );
  AOI22_X1 U72526 ( .A1(n86375), .A2(n74109), .B1(n86376), .B2(n110740), .ZN(
        n86947) );
  NAND2_X1 U72527 ( .A1(n86949), .A2(n86950), .ZN(n86939) );
  AOI22_X1 U72528 ( .A1(n86379), .A2(n110725), .B1(n86380), .B2(n110730), .ZN(
        n86950) );
  AOI22_X1 U72529 ( .A1(n86381), .A2(n74104), .B1(n105748), .B2(n110728), .ZN(
        n86949) );
  NAND2_X1 U72530 ( .A1(n86951), .A2(n86952), .ZN(n86923) );
  NOR4_X1 U72531 ( .A1(n86953), .A2(n86954), .A3(n86955), .A4(n86956), .ZN(
        n86952) );
  NAND2_X1 U72532 ( .A1(n86957), .A2(n86958), .ZN(n86956) );
  AOI22_X1 U72533 ( .A1(n86391), .A2(n110670), .B1(n86392), .B2(n110672), .ZN(
        n86958) );
  AOI22_X1 U72534 ( .A1(n86393), .A2(n74022), .B1(n86394), .B2(n110671), .ZN(
        n86957) );
  NAND2_X1 U72535 ( .A1(n86959), .A2(n86960), .ZN(n86955) );
  AOI22_X1 U72536 ( .A1(n86397), .A2(n74026), .B1(n86398), .B2(n74028), .ZN(
        n86960) );
  AOI22_X1 U72537 ( .A1(n86399), .A2(n110677), .B1(n105740), .B2(n110678), 
        .ZN(n86959) );
  NAND2_X1 U72538 ( .A1(n86961), .A2(n86962), .ZN(n86954) );
  AOI22_X1 U72539 ( .A1(n105739), .A2(n110675), .B1(n86404), .B2(n110676), 
        .ZN(n86962) );
  AOI22_X1 U72540 ( .A1(n86405), .A2(n110679), .B1(n105736), .B2(n74021), .ZN(
        n86961) );
  NAND2_X1 U72541 ( .A1(n86963), .A2(n86964), .ZN(n86953) );
  AOI22_X1 U72542 ( .A1(n86409), .A2(n110683), .B1(n86410), .B2(n74033), .ZN(
        n86964) );
  AOI22_X1 U72543 ( .A1(n105733), .A2(n110682), .B1(n86412), .B2(n74031), .ZN(
        n86963) );
  NOR4_X1 U72544 ( .A1(n86965), .A2(n86966), .A3(n86967), .A4(n86968), .ZN(
        n86951) );
  NAND2_X1 U72545 ( .A1(n86969), .A2(n86970), .ZN(n86968) );
  AOI22_X1 U72546 ( .A1(n86419), .A2(n110665), .B1(n86420), .B2(n110656), .ZN(
        n86970) );
  AOI22_X1 U72547 ( .A1(n86421), .A2(n110658), .B1(n86422), .B2(n74005), .ZN(
        n86969) );
  NAND2_X1 U72548 ( .A1(n86971), .A2(n86972), .ZN(n86967) );
  AOI22_X1 U72549 ( .A1(n86425), .A2(n110663), .B1(n105726), .B2(n110667), 
        .ZN(n86972) );
  AOI22_X1 U72550 ( .A1(n105725), .A2(n110669), .B1(n105724), .B2(n110666), 
        .ZN(n86971) );
  NAND2_X1 U72551 ( .A1(n86973), .A2(n86974), .ZN(n86966) );
  AOI22_X1 U72552 ( .A1(n86431), .A2(n74014), .B1(n86432), .B2(n110662), .ZN(
        n86974) );
  AOI22_X1 U72553 ( .A1(n86433), .A2(n110664), .B1(n86434), .B2(n110668), .ZN(
        n86973) );
  NAND2_X1 U72554 ( .A1(n86975), .A2(n86976), .ZN(n86965) );
  AOI22_X1 U72555 ( .A1(n86437), .A2(n110674), .B1(n86438), .B2(n74018), .ZN(
        n86976) );
  AOI22_X1 U72556 ( .A1(n86439), .A2(n74016), .B1(n105716), .B2(n110673), .ZN(
        n86975) );
  NAND2_X1 U72557 ( .A1(n86977), .A2(n86978), .ZN(n86922) );
  NOR4_X1 U72558 ( .A1(n86979), .A2(n86980), .A3(n86981), .A4(n86982), .ZN(
        n86978) );
  NAND2_X1 U72559 ( .A1(n86983), .A2(n86984), .ZN(n86982) );
  AOI22_X1 U72560 ( .A1(n86449), .A2(n74056), .B1(n105714), .B2(n110692), .ZN(
        n86984) );
  AOI22_X1 U72561 ( .A1(n86451), .A2(n110695), .B1(n86452), .B2(n74052), .ZN(
        n86983) );
  NAND2_X1 U72562 ( .A1(n86985), .A2(n86986), .ZN(n86981) );
  AOI22_X1 U72563 ( .A1(n105711), .A2(n110698), .B1(n86456), .B2(n110697), 
        .ZN(n86986) );
  AOI22_X1 U72564 ( .A1(n105709), .A2(n110691), .B1(n105708), .B2(n110693), 
        .ZN(n86985) );
  NAND2_X1 U72565 ( .A1(n86987), .A2(n86988), .ZN(n86980) );
  AOI22_X1 U72566 ( .A1(n86461), .A2(n74061), .B1(n86462), .B2(n74055), .ZN(
        n86988) );
  AOI22_X1 U72567 ( .A1(n86463), .A2(n74060), .B1(n86464), .B2(n74062), .ZN(
        n86987) );
  NAND2_X1 U72568 ( .A1(n86989), .A2(n86990), .ZN(n86979) );
  AOI22_X1 U72569 ( .A1(n105703), .A2(n74065), .B1(n86468), .B2(n74068), .ZN(
        n86990) );
  AOI22_X1 U72570 ( .A1(n86469), .A2(n110696), .B1(n86470), .B2(n74057), .ZN(
        n86989) );
  NOR4_X1 U72571 ( .A1(n86991), .A2(n86992), .A3(n86993), .A4(n86994), .ZN(
        n86977) );
  NAND2_X1 U72572 ( .A1(n86995), .A2(n86996), .ZN(n86994) );
  AOI22_X1 U72573 ( .A1(n86477), .A2(n74032), .B1(n86478), .B2(n110686), .ZN(
        n86996) );
  AOI22_X1 U72574 ( .A1(n105697), .A2(n110681), .B1(n86480), .B2(n74036), .ZN(
        n86995) );
  NAND2_X1 U72575 ( .A1(n86997), .A2(n86998), .ZN(n86993) );
  AOI22_X1 U72576 ( .A1(n86483), .A2(n74045), .B1(n105694), .B2(n110688), .ZN(
        n86998) );
  AOI22_X1 U72577 ( .A1(n86485), .A2(n110689), .B1(n86486), .B2(n110680), .ZN(
        n86997) );
  NAND2_X1 U72578 ( .A1(n86999), .A2(n87000), .ZN(n86992) );
  AOI22_X1 U72579 ( .A1(n86489), .A2(n110687), .B1(n105690), .B2(n74044), .ZN(
        n87000) );
  AOI22_X1 U72580 ( .A1(n86491), .A2(n110685), .B1(n86492), .B2(n110690), .ZN(
        n86999) );
  NAND2_X1 U72581 ( .A1(n87001), .A2(n87002), .ZN(n86991) );
  AOI22_X1 U72582 ( .A1(n105687), .A2(n74050), .B1(n86496), .B2(n110694), .ZN(
        n87002) );
  AOI22_X1 U72583 ( .A1(n86497), .A2(n74048), .B1(n86498), .B2(n110684), .ZN(
        n87001) );
  NAND2_X1 U72584 ( .A1(n87003), .A2(n87004), .ZN(n86921) );
  NOR4_X1 U72585 ( .A1(n87005), .A2(n87006), .A3(n87007), .A4(n87008), .ZN(
        n87004) );
  NAND2_X1 U72586 ( .A1(n87009), .A2(n87010), .ZN(n87008) );
  AOI22_X1 U72587 ( .A1(n86507), .A2(n110715), .B1(n86508), .B2(n110714), .ZN(
        n87010) );
  AOI22_X1 U72588 ( .A1(n86509), .A2(n74084), .B1(n86510), .B2(n110712), .ZN(
        n87009) );
  NAND2_X1 U72589 ( .A1(n87011), .A2(n87012), .ZN(n87007) );
  AOI22_X1 U72590 ( .A1(n86513), .A2(n110710), .B1(n105678), .B2(n110713), 
        .ZN(n87012) );
  AOI22_X1 U72591 ( .A1(n86515), .A2(n74090), .B1(n105677), .B2(n110711), .ZN(
        n87011) );
  NAND2_X1 U72592 ( .A1(n87013), .A2(n87014), .ZN(n87006) );
  AOI22_X1 U72593 ( .A1(n86519), .A2(n110720), .B1(n86520), .B2(n74096), .ZN(
        n87014) );
  AOI22_X1 U72594 ( .A1(n86521), .A2(n110718), .B1(n86522), .B2(n110719), .ZN(
        n87013) );
  NAND2_X1 U72595 ( .A1(n87015), .A2(n87016), .ZN(n87005) );
  AOI22_X1 U72596 ( .A1(n86525), .A2(n74088), .B1(n86526), .B2(n110717), .ZN(
        n87016) );
  AOI22_X1 U72597 ( .A1(n86527), .A2(n74095), .B1(n86528), .B2(n110716), .ZN(
        n87015) );
  NOR4_X1 U72598 ( .A1(n87017), .A2(n87018), .A3(n87019), .A4(n87020), .ZN(
        n87003) );
  NAND2_X1 U72599 ( .A1(n87021), .A2(n87022), .ZN(n87020) );
  AOI22_X1 U72600 ( .A1(n105675), .A2(n110700), .B1(n86536), .B2(n110702), 
        .ZN(n87022) );
  AOI22_X1 U72601 ( .A1(n86537), .A2(n74069), .B1(n86538), .B2(n74067), .ZN(
        n87021) );
  NAND2_X1 U72602 ( .A1(n87023), .A2(n87024), .ZN(n87019) );
  AOI22_X1 U72603 ( .A1(n86541), .A2(n110707), .B1(n86542), .B2(n110699), .ZN(
        n87024) );
  AOI22_X1 U72604 ( .A1(n86543), .A2(n110701), .B1(n105668), .B2(n110704), 
        .ZN(n87023) );
  NAND2_X1 U72605 ( .A1(n87025), .A2(n87026), .ZN(n87018) );
  AOI22_X1 U72606 ( .A1(n86547), .A2(n110703), .B1(n86548), .B2(n74077), .ZN(
        n87026) );
  AOI22_X1 U72607 ( .A1(n105665), .A2(n110709), .B1(n86550), .B2(n110706), 
        .ZN(n87025) );
  NAND2_X1 U72608 ( .A1(n87027), .A2(n87028), .ZN(n87017) );
  AOI22_X1 U72609 ( .A1(n86553), .A2(n74085), .B1(n86554), .B2(n74071), .ZN(
        n87028) );
  AOI22_X1 U72610 ( .A1(n105661), .A2(n110705), .B1(n86556), .B2(n110708), 
        .ZN(n87027) );
  AOI21_X1 U72611 ( .B1(n86302), .B2(n87030), .A(n87031), .ZN(n87029) );
  OAI21_X1 U72612 ( .B1(n87032), .B2(n86306), .A(n87033), .ZN(n87031) );
  OAI21_X1 U72613 ( .B1(n87034), .B2(n87035), .A(n105786), .ZN(n87033) );
  OAI21_X1 U72614 ( .B1(n108150), .B2(n86311), .A(n87036), .ZN(n87035) );
  AOI22_X1 U72615 ( .A1(n86313), .A2(n70711), .B1(n105784), .B2(n108148), .ZN(
        n87036) );
  NAND2_X1 U72616 ( .A1(n87037), .A2(n87038), .ZN(n87034) );
  AOI22_X1 U72617 ( .A1(n86317), .A2(n108146), .B1(n86318), .B2(n108151), .ZN(
        n87038) );
  AOI22_X1 U72618 ( .A1(n86319), .A2(n108149), .B1(n86320), .B2(n108147), .ZN(
        n87037) );
  NOR4_X1 U72619 ( .A1(n87039), .A2(n87040), .A3(n87041), .A4(n87042), .ZN(
        n87032) );
  NAND2_X1 U72620 ( .A1(n87043), .A2(n87044), .ZN(n87042) );
  NOR4_X1 U72621 ( .A1(n87045), .A2(n87046), .A3(n87047), .A4(n87048), .ZN(
        n87044) );
  NAND2_X1 U72622 ( .A1(n87049), .A2(n87050), .ZN(n87048) );
  AOI22_X1 U72623 ( .A1(n86333), .A2(n108126), .B1(n86334), .B2(n108127), .ZN(
        n87050) );
  AOI22_X1 U72624 ( .A1(n86335), .A2(n108136), .B1(n86336), .B2(n108134), .ZN(
        n87049) );
  NAND2_X1 U72625 ( .A1(n87051), .A2(n87052), .ZN(n87047) );
  AOI22_X1 U72626 ( .A1(n86339), .A2(n70580), .B1(n86340), .B2(n108130), .ZN(
        n87052) );
  AOI22_X1 U72627 ( .A1(n86341), .A2(n70684), .B1(n86342), .B2(n108054), .ZN(
        n87051) );
  NAND2_X1 U72628 ( .A1(n87053), .A2(n87054), .ZN(n87046) );
  AOI22_X1 U72629 ( .A1(n86345), .A2(n108058), .B1(n105770), .B2(n70584), .ZN(
        n87054) );
  AOI22_X1 U72630 ( .A1(n86347), .A2(n108131), .B1(n86348), .B2(n108128), .ZN(
        n87053) );
  NAND2_X1 U72631 ( .A1(n87055), .A2(n87056), .ZN(n87045) );
  AOI22_X1 U72632 ( .A1(n86351), .A2(n108056), .B1(n86352), .B2(n108060), .ZN(
        n87056) );
  AOI22_X1 U72633 ( .A1(n86353), .A2(n108059), .B1(n86354), .B2(n70586), .ZN(
        n87055) );
  NOR4_X1 U72634 ( .A1(n87057), .A2(n87058), .A3(n87059), .A4(n87060), .ZN(
        n87043) );
  NAND2_X1 U72635 ( .A1(n87061), .A2(n87062), .ZN(n87060) );
  AOI22_X1 U72636 ( .A1(n86361), .A2(n108137), .B1(n86362), .B2(n108140), .ZN(
        n87062) );
  AOI22_X1 U72637 ( .A1(n105761), .A2(n108141), .B1(n105760), .B2(n108143), 
        .ZN(n87061) );
  NAND2_X1 U72638 ( .A1(n87063), .A2(n87064), .ZN(n87059) );
  AOI22_X1 U72639 ( .A1(n86367), .A2(n108142), .B1(n105758), .B2(n108138), 
        .ZN(n87064) );
  AOI22_X1 U72640 ( .A1(n86369), .A2(n108144), .B1(n86370), .B2(n108139), .ZN(
        n87063) );
  NAND2_X1 U72641 ( .A1(n87065), .A2(n87066), .ZN(n87058) );
  AOI22_X1 U72642 ( .A1(n86373), .A2(n70694), .B1(n86374), .B2(n70693), .ZN(
        n87066) );
  AOI22_X1 U72643 ( .A1(n86375), .A2(n70696), .B1(n86376), .B2(n108145), .ZN(
        n87065) );
  NAND2_X1 U72644 ( .A1(n87067), .A2(n87068), .ZN(n87057) );
  AOI22_X1 U72645 ( .A1(n86379), .A2(n108129), .B1(n86380), .B2(n108135), .ZN(
        n87068) );
  AOI22_X1 U72646 ( .A1(n86381), .A2(n70691), .B1(n105748), .B2(n108133), .ZN(
        n87067) );
  NAND2_X1 U72647 ( .A1(n87069), .A2(n87070), .ZN(n87041) );
  NOR4_X1 U72648 ( .A1(n87071), .A2(n87072), .A3(n87073), .A4(n87074), .ZN(
        n87070) );
  NAND2_X1 U72649 ( .A1(n87075), .A2(n87076), .ZN(n87074) );
  AOI22_X1 U72650 ( .A1(n86391), .A2(n108069), .B1(n86392), .B2(n108071), .ZN(
        n87076) );
  AOI22_X1 U72651 ( .A1(n86393), .A2(n70609), .B1(n86394), .B2(n108070), .ZN(
        n87075) );
  NAND2_X1 U72652 ( .A1(n87077), .A2(n87078), .ZN(n87073) );
  AOI22_X1 U72653 ( .A1(n86397), .A2(n70613), .B1(n86398), .B2(n70615), .ZN(
        n87078) );
  AOI22_X1 U72654 ( .A1(n86399), .A2(n108077), .B1(n105740), .B2(n108078), 
        .ZN(n87077) );
  NAND2_X1 U72655 ( .A1(n87079), .A2(n87080), .ZN(n87072) );
  AOI22_X1 U72656 ( .A1(n105739), .A2(n108074), .B1(n86404), .B2(n108076), 
        .ZN(n87080) );
  AOI22_X1 U72657 ( .A1(n86405), .A2(n108079), .B1(n105736), .B2(n108075), 
        .ZN(n87079) );
  NAND2_X1 U72658 ( .A1(n87081), .A2(n87082), .ZN(n87071) );
  AOI22_X1 U72659 ( .A1(n86409), .A2(n108083), .B1(n86410), .B2(n70620), .ZN(
        n87082) );
  AOI22_X1 U72660 ( .A1(n105733), .A2(n108082), .B1(n86412), .B2(n70618), .ZN(
        n87081) );
  NOR4_X1 U72661 ( .A1(n87083), .A2(n87084), .A3(n87085), .A4(n87086), .ZN(
        n87069) );
  NAND2_X1 U72662 ( .A1(n87087), .A2(n87088), .ZN(n87086) );
  AOI22_X1 U72663 ( .A1(n86419), .A2(n108064), .B1(n86420), .B2(n108055), .ZN(
        n87088) );
  AOI22_X1 U72664 ( .A1(n86421), .A2(n108057), .B1(n86422), .B2(n70592), .ZN(
        n87087) );
  NAND2_X1 U72665 ( .A1(n87089), .A2(n87090), .ZN(n87085) );
  AOI22_X1 U72666 ( .A1(n86425), .A2(n108062), .B1(n105726), .B2(n108066), 
        .ZN(n87090) );
  AOI22_X1 U72667 ( .A1(n105725), .A2(n108068), .B1(n105724), .B2(n108065), 
        .ZN(n87089) );
  NAND2_X1 U72668 ( .A1(n87091), .A2(n87092), .ZN(n87084) );
  AOI22_X1 U72669 ( .A1(n86431), .A2(n70601), .B1(n86432), .B2(n108061), .ZN(
        n87092) );
  AOI22_X1 U72670 ( .A1(n86433), .A2(n108063), .B1(n86434), .B2(n108067), .ZN(
        n87091) );
  NAND2_X1 U72671 ( .A1(n87093), .A2(n87094), .ZN(n87083) );
  AOI22_X1 U72672 ( .A1(n86437), .A2(n108073), .B1(n86438), .B2(n70605), .ZN(
        n87094) );
  AOI22_X1 U72673 ( .A1(n86439), .A2(n70603), .B1(n105716), .B2(n108072), .ZN(
        n87093) );
  NAND2_X1 U72674 ( .A1(n87095), .A2(n87096), .ZN(n87040) );
  NOR4_X1 U72675 ( .A1(n87097), .A2(n87098), .A3(n87099), .A4(n87100), .ZN(
        n87096) );
  NAND2_X1 U72676 ( .A1(n87101), .A2(n87102), .ZN(n87100) );
  AOI22_X1 U72677 ( .A1(n86449), .A2(n70643), .B1(n105714), .B2(n108092), .ZN(
        n87102) );
  AOI22_X1 U72678 ( .A1(n86451), .A2(n108095), .B1(n86452), .B2(n70639), .ZN(
        n87101) );
  NAND2_X1 U72679 ( .A1(n87103), .A2(n87104), .ZN(n87099) );
  AOI22_X1 U72680 ( .A1(n105711), .A2(n108100), .B1(n86456), .B2(n108099), 
        .ZN(n87104) );
  AOI22_X1 U72681 ( .A1(n105709), .A2(n108091), .B1(n86458), .B2(n108093), 
        .ZN(n87103) );
  NAND2_X1 U72682 ( .A1(n87105), .A2(n87106), .ZN(n87098) );
  AOI22_X1 U72683 ( .A1(n86461), .A2(n108101), .B1(n86462), .B2(n108097), .ZN(
        n87106) );
  AOI22_X1 U72684 ( .A1(n86463), .A2(n70647), .B1(n86464), .B2(n70649), .ZN(
        n87105) );
  NAND2_X1 U72685 ( .A1(n87107), .A2(n87108), .ZN(n87097) );
  AOI22_X1 U72686 ( .A1(n105703), .A2(n70652), .B1(n86468), .B2(n70655), .ZN(
        n87108) );
  AOI22_X1 U72687 ( .A1(n86469), .A2(n108096), .B1(n86470), .B2(n108098), .ZN(
        n87107) );
  NOR4_X1 U72688 ( .A1(n87109), .A2(n87110), .A3(n87111), .A4(n87112), .ZN(
        n87095) );
  NAND2_X1 U72689 ( .A1(n87113), .A2(n87114), .ZN(n87112) );
  AOI22_X1 U72690 ( .A1(n86477), .A2(n70619), .B1(n86478), .B2(n108086), .ZN(
        n87114) );
  AOI22_X1 U72691 ( .A1(n105697), .A2(n108081), .B1(n86480), .B2(n70623), .ZN(
        n87113) );
  NAND2_X1 U72692 ( .A1(n87115), .A2(n87116), .ZN(n87111) );
  AOI22_X1 U72693 ( .A1(n86483), .A2(n70632), .B1(n105694), .B2(n108088), .ZN(
        n87116) );
  AOI22_X1 U72694 ( .A1(n86485), .A2(n108089), .B1(n86486), .B2(n108080), .ZN(
        n87115) );
  NAND2_X1 U72695 ( .A1(n87117), .A2(n87118), .ZN(n87110) );
  AOI22_X1 U72696 ( .A1(n86489), .A2(n108087), .B1(n105690), .B2(n70631), .ZN(
        n87118) );
  AOI22_X1 U72697 ( .A1(n86491), .A2(n108085), .B1(n86492), .B2(n108090), .ZN(
        n87117) );
  NAND2_X1 U72698 ( .A1(n87119), .A2(n87120), .ZN(n87109) );
  AOI22_X1 U72699 ( .A1(n105687), .A2(n70637), .B1(n86496), .B2(n108094), .ZN(
        n87120) );
  AOI22_X1 U72700 ( .A1(n86497), .A2(n70635), .B1(n86498), .B2(n108084), .ZN(
        n87119) );
  NAND2_X1 U72701 ( .A1(n87121), .A2(n87122), .ZN(n87039) );
  NOR4_X1 U72702 ( .A1(n87123), .A2(n87124), .A3(n87125), .A4(n87126), .ZN(
        n87122) );
  NAND2_X1 U72703 ( .A1(n87127), .A2(n87128), .ZN(n87126) );
  AOI22_X1 U72704 ( .A1(n86507), .A2(n108118), .B1(n86508), .B2(n108117), .ZN(
        n87128) );
  AOI22_X1 U72705 ( .A1(n86509), .A2(n70671), .B1(n86510), .B2(n108115), .ZN(
        n87127) );
  NAND2_X1 U72706 ( .A1(n87129), .A2(n87130), .ZN(n87125) );
  AOI22_X1 U72707 ( .A1(n86513), .A2(n108113), .B1(n105678), .B2(n108116), 
        .ZN(n87130) );
  AOI22_X1 U72708 ( .A1(n86515), .A2(n70677), .B1(n105677), .B2(n108114), .ZN(
        n87129) );
  NAND2_X1 U72709 ( .A1(n87131), .A2(n87132), .ZN(n87124) );
  AOI22_X1 U72710 ( .A1(n86519), .A2(n108123), .B1(n86520), .B2(n70683), .ZN(
        n87132) );
  AOI22_X1 U72711 ( .A1(n86521), .A2(n108121), .B1(n86522), .B2(n108122), .ZN(
        n87131) );
  NAND2_X1 U72712 ( .A1(n87133), .A2(n87134), .ZN(n87123) );
  AOI22_X1 U72713 ( .A1(n86525), .A2(n70675), .B1(n86526), .B2(n108120), .ZN(
        n87134) );
  AOI22_X1 U72714 ( .A1(n86527), .A2(n108124), .B1(n86528), .B2(n108119), .ZN(
        n87133) );
  NOR4_X1 U72715 ( .A1(n87135), .A2(n87136), .A3(n87137), .A4(n87138), .ZN(
        n87121) );
  NAND2_X1 U72716 ( .A1(n87139), .A2(n87140), .ZN(n87138) );
  AOI22_X1 U72717 ( .A1(n105675), .A2(n108103), .B1(n86536), .B2(n108105), 
        .ZN(n87140) );
  AOI22_X1 U72718 ( .A1(n86537), .A2(n70656), .B1(n86538), .B2(n70654), .ZN(
        n87139) );
  NAND2_X1 U72719 ( .A1(n87141), .A2(n87142), .ZN(n87137) );
  AOI22_X1 U72720 ( .A1(n86541), .A2(n108110), .B1(n86542), .B2(n108102), .ZN(
        n87142) );
  AOI22_X1 U72721 ( .A1(n86543), .A2(n108104), .B1(n105668), .B2(n108107), 
        .ZN(n87141) );
  NAND2_X1 U72722 ( .A1(n87143), .A2(n87144), .ZN(n87136) );
  AOI22_X1 U72723 ( .A1(n86547), .A2(n108106), .B1(n86548), .B2(n70664), .ZN(
        n87144) );
  AOI22_X1 U72724 ( .A1(n105665), .A2(n108112), .B1(n86550), .B2(n108109), 
        .ZN(n87143) );
  NAND2_X1 U72725 ( .A1(n87145), .A2(n87146), .ZN(n87135) );
  AOI22_X1 U72726 ( .A1(n86553), .A2(n70672), .B1(n86554), .B2(n70658), .ZN(
        n87146) );
  AOI22_X1 U72727 ( .A1(n105661), .A2(n108108), .B1(n86556), .B2(n108111), 
        .ZN(n87145) );
  AOI21_X1 U72728 ( .B1(n86302), .B2(n87148), .A(n87149), .ZN(n87147) );
  OAI21_X1 U72729 ( .B1(n87150), .B2(n86306), .A(n87151), .ZN(n87149) );
  OAI21_X1 U72730 ( .B1(n87152), .B2(n87153), .A(n105786), .ZN(n87151) );
  OAI21_X1 U72731 ( .B1(n110848), .B2(n86311), .A(n87154), .ZN(n87153) );
  AOI22_X1 U72732 ( .A1(n86313), .A2(n74265), .B1(n105784), .B2(n110846), .ZN(
        n87154) );
  NAND2_X1 U72733 ( .A1(n87155), .A2(n87156), .ZN(n87152) );
  AOI22_X1 U72734 ( .A1(n86317), .A2(n110844), .B1(n86318), .B2(n110849), .ZN(
        n87156) );
  AOI22_X1 U72735 ( .A1(n86319), .A2(n110847), .B1(n86320), .B2(n110845), .ZN(
        n87155) );
  NOR4_X1 U72736 ( .A1(n87157), .A2(n87158), .A3(n87159), .A4(n87160), .ZN(
        n87150) );
  NAND2_X1 U72737 ( .A1(n87161), .A2(n87162), .ZN(n87160) );
  NOR4_X1 U72738 ( .A1(n87163), .A2(n87164), .A3(n87165), .A4(n87166), .ZN(
        n87162) );
  NAND2_X1 U72739 ( .A1(n87167), .A2(n87168), .ZN(n87166) );
  AOI22_X1 U72740 ( .A1(n86333), .A2(n110825), .B1(n86334), .B2(n110826), .ZN(
        n87168) );
  AOI22_X1 U72741 ( .A1(n86335), .A2(n110834), .B1(n86336), .B2(n110832), .ZN(
        n87167) );
  NAND2_X1 U72742 ( .A1(n87169), .A2(n87170), .ZN(n87165) );
  AOI22_X1 U72743 ( .A1(n86339), .A2(n74134), .B1(n86340), .B2(n110829), .ZN(
        n87170) );
  AOI22_X1 U72744 ( .A1(n86341), .A2(n74238), .B1(n86342), .B2(n110752), .ZN(
        n87169) );
  NAND2_X1 U72745 ( .A1(n87171), .A2(n87172), .ZN(n87164) );
  AOI22_X1 U72746 ( .A1(n86345), .A2(n110756), .B1(n105770), .B2(n74138), .ZN(
        n87172) );
  AOI22_X1 U72747 ( .A1(n86347), .A2(n110830), .B1(n86348), .B2(n110827), .ZN(
        n87171) );
  NAND2_X1 U72748 ( .A1(n87173), .A2(n87174), .ZN(n87163) );
  AOI22_X1 U72749 ( .A1(n86351), .A2(n110754), .B1(n86352), .B2(n110758), .ZN(
        n87174) );
  AOI22_X1 U72750 ( .A1(n86353), .A2(n110757), .B1(n86354), .B2(n74140), .ZN(
        n87173) );
  NOR4_X1 U72751 ( .A1(n87175), .A2(n87176), .A3(n87177), .A4(n87178), .ZN(
        n87161) );
  NAND2_X1 U72752 ( .A1(n87179), .A2(n87180), .ZN(n87178) );
  AOI22_X1 U72753 ( .A1(n86361), .A2(n110835), .B1(n86362), .B2(n110838), .ZN(
        n87180) );
  AOI22_X1 U72754 ( .A1(n105761), .A2(n110839), .B1(n105760), .B2(n110841), 
        .ZN(n87179) );
  NAND2_X1 U72755 ( .A1(n87181), .A2(n87182), .ZN(n87177) );
  AOI22_X1 U72756 ( .A1(n86367), .A2(n110840), .B1(n105758), .B2(n110836), 
        .ZN(n87182) );
  AOI22_X1 U72757 ( .A1(n86369), .A2(n110842), .B1(n86370), .B2(n110837), .ZN(
        n87181) );
  NAND2_X1 U72758 ( .A1(n87183), .A2(n87184), .ZN(n87176) );
  AOI22_X1 U72759 ( .A1(n86373), .A2(n74248), .B1(n86374), .B2(n74247), .ZN(
        n87184) );
  AOI22_X1 U72760 ( .A1(n86375), .A2(n74250), .B1(n86376), .B2(n110843), .ZN(
        n87183) );
  NAND2_X1 U72761 ( .A1(n87185), .A2(n87186), .ZN(n87175) );
  AOI22_X1 U72762 ( .A1(n86379), .A2(n110828), .B1(n86380), .B2(n110833), .ZN(
        n87186) );
  AOI22_X1 U72763 ( .A1(n86381), .A2(n74245), .B1(n105748), .B2(n110831), .ZN(
        n87185) );
  NAND2_X1 U72764 ( .A1(n87187), .A2(n87188), .ZN(n87159) );
  NOR4_X1 U72765 ( .A1(n87189), .A2(n87190), .A3(n87191), .A4(n87192), .ZN(
        n87188) );
  NAND2_X1 U72766 ( .A1(n87193), .A2(n87194), .ZN(n87192) );
  AOI22_X1 U72767 ( .A1(n86391), .A2(n110767), .B1(n86392), .B2(n110769), .ZN(
        n87194) );
  AOI22_X1 U72768 ( .A1(n86393), .A2(n74163), .B1(n86394), .B2(n110768), .ZN(
        n87193) );
  NAND2_X1 U72769 ( .A1(n87195), .A2(n87196), .ZN(n87191) );
  AOI22_X1 U72770 ( .A1(n86397), .A2(n74167), .B1(n86398), .B2(n74169), .ZN(
        n87196) );
  AOI22_X1 U72771 ( .A1(n86399), .A2(n110774), .B1(n105740), .B2(n110775), 
        .ZN(n87195) );
  NAND2_X1 U72772 ( .A1(n87197), .A2(n87198), .ZN(n87190) );
  AOI22_X1 U72773 ( .A1(n105739), .A2(n110772), .B1(n86404), .B2(n110773), 
        .ZN(n87198) );
  AOI22_X1 U72774 ( .A1(n86405), .A2(n110776), .B1(n105736), .B2(n74162), .ZN(
        n87197) );
  NAND2_X1 U72775 ( .A1(n87199), .A2(n87200), .ZN(n87189) );
  AOI22_X1 U72776 ( .A1(n86409), .A2(n110781), .B1(n86410), .B2(n74174), .ZN(
        n87200) );
  AOI22_X1 U72777 ( .A1(n105733), .A2(n110780), .B1(n86412), .B2(n74172), .ZN(
        n87199) );
  NOR4_X1 U72778 ( .A1(n87201), .A2(n87202), .A3(n87203), .A4(n87204), .ZN(
        n87187) );
  NAND2_X1 U72779 ( .A1(n87205), .A2(n87206), .ZN(n87204) );
  AOI22_X1 U72780 ( .A1(n86419), .A2(n110762), .B1(n86420), .B2(n110753), .ZN(
        n87206) );
  AOI22_X1 U72781 ( .A1(n86421), .A2(n110755), .B1(n86422), .B2(n74146), .ZN(
        n87205) );
  NAND2_X1 U72782 ( .A1(n87207), .A2(n87208), .ZN(n87203) );
  AOI22_X1 U72783 ( .A1(n86425), .A2(n110760), .B1(n105726), .B2(n110764), 
        .ZN(n87208) );
  AOI22_X1 U72784 ( .A1(n105725), .A2(n110766), .B1(n105724), .B2(n110763), 
        .ZN(n87207) );
  NAND2_X1 U72785 ( .A1(n87209), .A2(n87210), .ZN(n87202) );
  AOI22_X1 U72786 ( .A1(n86431), .A2(n74155), .B1(n86432), .B2(n110759), .ZN(
        n87210) );
  AOI22_X1 U72787 ( .A1(n86433), .A2(n110761), .B1(n86434), .B2(n110765), .ZN(
        n87209) );
  NAND2_X1 U72788 ( .A1(n87211), .A2(n87212), .ZN(n87201) );
  AOI22_X1 U72789 ( .A1(n86437), .A2(n110771), .B1(n86438), .B2(n74159), .ZN(
        n87212) );
  AOI22_X1 U72790 ( .A1(n86439), .A2(n74157), .B1(n105716), .B2(n110770), .ZN(
        n87211) );
  NAND2_X1 U72791 ( .A1(n87213), .A2(n87214), .ZN(n87158) );
  NOR4_X1 U72792 ( .A1(n87215), .A2(n87216), .A3(n87217), .A4(n87218), .ZN(
        n87214) );
  NAND2_X1 U72793 ( .A1(n87219), .A2(n87220), .ZN(n87218) );
  AOI22_X1 U72794 ( .A1(n86449), .A2(n74197), .B1(n105714), .B2(n110791), .ZN(
        n87220) );
  AOI22_X1 U72795 ( .A1(n86451), .A2(n110795), .B1(n86452), .B2(n110794), .ZN(
        n87219) );
  NAND2_X1 U72796 ( .A1(n87221), .A2(n87222), .ZN(n87217) );
  AOI22_X1 U72797 ( .A1(n105711), .A2(n110799), .B1(n86456), .B2(n110798), 
        .ZN(n87222) );
  AOI22_X1 U72798 ( .A1(n105709), .A2(n110790), .B1(n86458), .B2(n110792), 
        .ZN(n87221) );
  NAND2_X1 U72799 ( .A1(n87223), .A2(n87224), .ZN(n87216) );
  AOI22_X1 U72800 ( .A1(n86461), .A2(n110800), .B1(n86462), .B2(n74196), .ZN(
        n87224) );
  AOI22_X1 U72801 ( .A1(n86463), .A2(n74201), .B1(n86464), .B2(n74203), .ZN(
        n87223) );
  NAND2_X1 U72802 ( .A1(n87225), .A2(n87226), .ZN(n87215) );
  AOI22_X1 U72803 ( .A1(n105703), .A2(n74206), .B1(n86468), .B2(n74209), .ZN(
        n87226) );
  AOI22_X1 U72804 ( .A1(n86469), .A2(n110796), .B1(n86470), .B2(n110797), .ZN(
        n87225) );
  NOR4_X1 U72805 ( .A1(n87227), .A2(n87228), .A3(n87229), .A4(n87230), .ZN(
        n87213) );
  NAND2_X1 U72806 ( .A1(n87231), .A2(n87232), .ZN(n87230) );
  AOI22_X1 U72807 ( .A1(n86477), .A2(n110779), .B1(n86478), .B2(n110784), .ZN(
        n87232) );
  AOI22_X1 U72808 ( .A1(n105697), .A2(n110778), .B1(n86480), .B2(n74177), .ZN(
        n87231) );
  NAND2_X1 U72809 ( .A1(n87233), .A2(n87234), .ZN(n87229) );
  AOI22_X1 U72810 ( .A1(n86483), .A2(n74186), .B1(n105694), .B2(n110786), .ZN(
        n87234) );
  AOI22_X1 U72811 ( .A1(n86485), .A2(n110787), .B1(n86486), .B2(n110777), .ZN(
        n87233) );
  NAND2_X1 U72812 ( .A1(n87235), .A2(n87236), .ZN(n87228) );
  AOI22_X1 U72813 ( .A1(n86489), .A2(n110785), .B1(n105690), .B2(n110789), 
        .ZN(n87236) );
  AOI22_X1 U72814 ( .A1(n86491), .A2(n110783), .B1(n86492), .B2(n110788), .ZN(
        n87235) );
  NAND2_X1 U72815 ( .A1(n87237), .A2(n87238), .ZN(n87227) );
  AOI22_X1 U72816 ( .A1(n105687), .A2(n74191), .B1(n86496), .B2(n110793), .ZN(
        n87238) );
  AOI22_X1 U72817 ( .A1(n86497), .A2(n74189), .B1(n86498), .B2(n110782), .ZN(
        n87237) );
  NAND2_X1 U72818 ( .A1(n87239), .A2(n87240), .ZN(n87157) );
  NOR4_X1 U72819 ( .A1(n87241), .A2(n87242), .A3(n87243), .A4(n87244), .ZN(
        n87240) );
  NAND2_X1 U72820 ( .A1(n87245), .A2(n87246), .ZN(n87244) );
  AOI22_X1 U72821 ( .A1(n86507), .A2(n110817), .B1(n86508), .B2(n110816), .ZN(
        n87246) );
  AOI22_X1 U72822 ( .A1(n86509), .A2(n74225), .B1(n86510), .B2(n110814), .ZN(
        n87245) );
  NAND2_X1 U72823 ( .A1(n87247), .A2(n87248), .ZN(n87243) );
  AOI22_X1 U72824 ( .A1(n86513), .A2(n110812), .B1(n105678), .B2(n110815), 
        .ZN(n87248) );
  AOI22_X1 U72825 ( .A1(n86515), .A2(n74231), .B1(n105677), .B2(n110813), .ZN(
        n87247) );
  NAND2_X1 U72826 ( .A1(n87249), .A2(n87250), .ZN(n87242) );
  AOI22_X1 U72827 ( .A1(n86519), .A2(n110822), .B1(n86520), .B2(n74237), .ZN(
        n87250) );
  AOI22_X1 U72828 ( .A1(n86521), .A2(n110820), .B1(n86522), .B2(n110821), .ZN(
        n87249) );
  NAND2_X1 U72829 ( .A1(n87251), .A2(n87252), .ZN(n87241) );
  AOI22_X1 U72830 ( .A1(n86525), .A2(n74229), .B1(n86526), .B2(n110819), .ZN(
        n87252) );
  AOI22_X1 U72831 ( .A1(n86527), .A2(n110823), .B1(n86528), .B2(n110818), .ZN(
        n87251) );
  NOR4_X1 U72832 ( .A1(n87253), .A2(n87254), .A3(n87255), .A4(n87256), .ZN(
        n87239) );
  NAND2_X1 U72833 ( .A1(n87257), .A2(n87258), .ZN(n87256) );
  AOI22_X1 U72834 ( .A1(n105675), .A2(n110802), .B1(n86536), .B2(n110804), 
        .ZN(n87258) );
  AOI22_X1 U72835 ( .A1(n86537), .A2(n74210), .B1(n86538), .B2(n74208), .ZN(
        n87257) );
  NAND2_X1 U72836 ( .A1(n87259), .A2(n87260), .ZN(n87255) );
  AOI22_X1 U72837 ( .A1(n86541), .A2(n110809), .B1(n86542), .B2(n110801), .ZN(
        n87260) );
  AOI22_X1 U72838 ( .A1(n86543), .A2(n110803), .B1(n105668), .B2(n110806), 
        .ZN(n87259) );
  NAND2_X1 U72839 ( .A1(n87261), .A2(n87262), .ZN(n87254) );
  AOI22_X1 U72840 ( .A1(n86547), .A2(n110805), .B1(n86548), .B2(n74218), .ZN(
        n87262) );
  AOI22_X1 U72841 ( .A1(n105665), .A2(n110811), .B1(n86550), .B2(n110808), 
        .ZN(n87261) );
  NAND2_X1 U72842 ( .A1(n87263), .A2(n87264), .ZN(n87253) );
  AOI22_X1 U72843 ( .A1(n86553), .A2(n74226), .B1(n86554), .B2(n74212), .ZN(
        n87264) );
  AOI22_X1 U72844 ( .A1(n105661), .A2(n110807), .B1(n86556), .B2(n110810), 
        .ZN(n87263) );
  AOI21_X1 U72845 ( .B1(n86302), .B2(n87266), .A(n87267), .ZN(n87265) );
  OAI21_X1 U72846 ( .B1(n87268), .B2(n86306), .A(n87269), .ZN(n87267) );
  OAI21_X1 U72847 ( .B1(n87270), .B2(n87271), .A(n105786), .ZN(n87269) );
  OAI21_X1 U72848 ( .B1(n110949), .B2(n86311), .A(n87272), .ZN(n87271) );
  AOI22_X1 U72849 ( .A1(n86313), .A2(n74405), .B1(n105784), .B2(n110947), .ZN(
        n87272) );
  NAND2_X1 U72850 ( .A1(n87273), .A2(n87274), .ZN(n87270) );
  AOI22_X1 U72851 ( .A1(n86317), .A2(n110945), .B1(n86318), .B2(n110950), .ZN(
        n87274) );
  AOI22_X1 U72852 ( .A1(n86319), .A2(n110948), .B1(n86320), .B2(n110946), .ZN(
        n87273) );
  NOR4_X1 U72853 ( .A1(n87275), .A2(n87276), .A3(n87277), .A4(n87278), .ZN(
        n87268) );
  NAND2_X1 U72854 ( .A1(n87279), .A2(n87280), .ZN(n87278) );
  NOR4_X1 U72855 ( .A1(n87281), .A2(n87282), .A3(n87283), .A4(n87284), .ZN(
        n87280) );
  NAND2_X1 U72856 ( .A1(n87285), .A2(n87286), .ZN(n87284) );
  AOI22_X1 U72857 ( .A1(n86333), .A2(n110926), .B1(n86334), .B2(n110927), .ZN(
        n87286) );
  AOI22_X1 U72858 ( .A1(n86335), .A2(n110935), .B1(n86336), .B2(n110933), .ZN(
        n87285) );
  NAND2_X1 U72859 ( .A1(n87287), .A2(n87288), .ZN(n87283) );
  AOI22_X1 U72860 ( .A1(n86339), .A2(n74274), .B1(n86340), .B2(n110930), .ZN(
        n87288) );
  AOI22_X1 U72861 ( .A1(n86341), .A2(n74378), .B1(n86342), .B2(n110853), .ZN(
        n87287) );
  NAND2_X1 U72862 ( .A1(n87289), .A2(n87290), .ZN(n87282) );
  AOI22_X1 U72863 ( .A1(n86345), .A2(n110857), .B1(n105770), .B2(n74278), .ZN(
        n87290) );
  AOI22_X1 U72864 ( .A1(n86347), .A2(n110931), .B1(n86348), .B2(n110928), .ZN(
        n87289) );
  NAND2_X1 U72865 ( .A1(n87291), .A2(n87292), .ZN(n87281) );
  AOI22_X1 U72866 ( .A1(n86351), .A2(n110855), .B1(n86352), .B2(n110859), .ZN(
        n87292) );
  AOI22_X1 U72867 ( .A1(n86353), .A2(n110858), .B1(n86354), .B2(n74280), .ZN(
        n87291) );
  NOR4_X1 U72868 ( .A1(n87293), .A2(n87294), .A3(n87295), .A4(n87296), .ZN(
        n87279) );
  NAND2_X1 U72869 ( .A1(n87297), .A2(n87298), .ZN(n87296) );
  AOI22_X1 U72870 ( .A1(n86361), .A2(n110936), .B1(n86362), .B2(n110939), .ZN(
        n87298) );
  AOI22_X1 U72871 ( .A1(n105761), .A2(n110940), .B1(n105760), .B2(n110942), 
        .ZN(n87297) );
  NAND2_X1 U72872 ( .A1(n87299), .A2(n87300), .ZN(n87295) );
  AOI22_X1 U72873 ( .A1(n86367), .A2(n110941), .B1(n105758), .B2(n110937), 
        .ZN(n87300) );
  AOI22_X1 U72874 ( .A1(n86369), .A2(n110943), .B1(n86370), .B2(n110938), .ZN(
        n87299) );
  NAND2_X1 U72875 ( .A1(n87301), .A2(n87302), .ZN(n87294) );
  AOI22_X1 U72876 ( .A1(n86373), .A2(n74388), .B1(n86374), .B2(n74387), .ZN(
        n87302) );
  AOI22_X1 U72877 ( .A1(n86375), .A2(n74390), .B1(n86376), .B2(n110944), .ZN(
        n87301) );
  NAND2_X1 U72878 ( .A1(n87303), .A2(n87304), .ZN(n87293) );
  AOI22_X1 U72879 ( .A1(n86379), .A2(n110929), .B1(n86380), .B2(n110934), .ZN(
        n87304) );
  AOI22_X1 U72880 ( .A1(n86381), .A2(n74385), .B1(n105748), .B2(n110932), .ZN(
        n87303) );
  NAND2_X1 U72881 ( .A1(n87305), .A2(n87306), .ZN(n87277) );
  NOR4_X1 U72882 ( .A1(n87307), .A2(n87308), .A3(n87309), .A4(n87310), .ZN(
        n87306) );
  NAND2_X1 U72883 ( .A1(n87311), .A2(n87312), .ZN(n87310) );
  AOI22_X1 U72884 ( .A1(n86391), .A2(n110868), .B1(n86392), .B2(n110870), .ZN(
        n87312) );
  AOI22_X1 U72885 ( .A1(n86393), .A2(n74303), .B1(n86394), .B2(n110869), .ZN(
        n87311) );
  NAND2_X1 U72886 ( .A1(n87313), .A2(n87314), .ZN(n87309) );
  AOI22_X1 U72887 ( .A1(n86397), .A2(n74307), .B1(n86398), .B2(n74309), .ZN(
        n87314) );
  AOI22_X1 U72888 ( .A1(n86399), .A2(n110875), .B1(n105740), .B2(n110876), 
        .ZN(n87313) );
  NAND2_X1 U72889 ( .A1(n87315), .A2(n87316), .ZN(n87308) );
  AOI22_X1 U72890 ( .A1(n105739), .A2(n110873), .B1(n86404), .B2(n110874), 
        .ZN(n87316) );
  AOI22_X1 U72891 ( .A1(n86405), .A2(n110877), .B1(n105736), .B2(n74302), .ZN(
        n87315) );
  NAND2_X1 U72892 ( .A1(n87317), .A2(n87318), .ZN(n87307) );
  AOI22_X1 U72893 ( .A1(n86409), .A2(n110882), .B1(n86410), .B2(n74314), .ZN(
        n87318) );
  AOI22_X1 U72894 ( .A1(n105733), .A2(n110881), .B1(n86412), .B2(n74312), .ZN(
        n87317) );
  NOR4_X1 U72895 ( .A1(n87319), .A2(n87320), .A3(n87321), .A4(n87322), .ZN(
        n87305) );
  NAND2_X1 U72896 ( .A1(n87323), .A2(n87324), .ZN(n87322) );
  AOI22_X1 U72897 ( .A1(n86419), .A2(n110863), .B1(n86420), .B2(n110854), .ZN(
        n87324) );
  AOI22_X1 U72898 ( .A1(n86421), .A2(n110856), .B1(n86422), .B2(n74286), .ZN(
        n87323) );
  NAND2_X1 U72899 ( .A1(n87325), .A2(n87326), .ZN(n87321) );
  AOI22_X1 U72900 ( .A1(n86425), .A2(n110861), .B1(n105726), .B2(n110865), 
        .ZN(n87326) );
  AOI22_X1 U72901 ( .A1(n105725), .A2(n110867), .B1(n105724), .B2(n110864), 
        .ZN(n87325) );
  NAND2_X1 U72902 ( .A1(n87327), .A2(n87328), .ZN(n87320) );
  AOI22_X1 U72903 ( .A1(n86431), .A2(n74295), .B1(n86432), .B2(n110860), .ZN(
        n87328) );
  AOI22_X1 U72904 ( .A1(n86433), .A2(n110862), .B1(n86434), .B2(n110866), .ZN(
        n87327) );
  NAND2_X1 U72905 ( .A1(n87329), .A2(n87330), .ZN(n87319) );
  AOI22_X1 U72906 ( .A1(n86437), .A2(n110872), .B1(n86438), .B2(n74299), .ZN(
        n87330) );
  AOI22_X1 U72907 ( .A1(n86439), .A2(n74297), .B1(n105716), .B2(n110871), .ZN(
        n87329) );
  NAND2_X1 U72908 ( .A1(n87331), .A2(n87332), .ZN(n87276) );
  NOR4_X1 U72909 ( .A1(n87333), .A2(n87334), .A3(n87335), .A4(n87336), .ZN(
        n87332) );
  NAND2_X1 U72910 ( .A1(n87337), .A2(n87338), .ZN(n87336) );
  AOI22_X1 U72911 ( .A1(n86449), .A2(n74337), .B1(n105714), .B2(n110891), .ZN(
        n87338) );
  AOI22_X1 U72912 ( .A1(n86451), .A2(n110894), .B1(n86452), .B2(n110893), .ZN(
        n87337) );
  NAND2_X1 U72913 ( .A1(n87339), .A2(n87340), .ZN(n87335) );
  AOI22_X1 U72914 ( .A1(n105711), .A2(n110897), .B1(n86456), .B2(n110896), 
        .ZN(n87340) );
  AOI22_X1 U72915 ( .A1(n105709), .A2(n110890), .B1(n86458), .B2(n111016), 
        .ZN(n87339) );
  NAND2_X1 U72916 ( .A1(n87341), .A2(n87342), .ZN(n87334) );
  AOI22_X1 U72917 ( .A1(n86461), .A2(n74342), .B1(n86462), .B2(n74336), .ZN(
        n87342) );
  AOI22_X1 U72918 ( .A1(n86463), .A2(n74341), .B1(n86464), .B2(n74343), .ZN(
        n87341) );
  NAND2_X1 U72919 ( .A1(n87343), .A2(n87344), .ZN(n87333) );
  AOI22_X1 U72920 ( .A1(n105703), .A2(n111037), .B1(n86468), .B2(n74349), .ZN(
        n87344) );
  AOI22_X1 U72921 ( .A1(n86469), .A2(n110895), .B1(n86470), .B2(n74338), .ZN(
        n87343) );
  NOR4_X1 U72922 ( .A1(n87345), .A2(n87346), .A3(n87347), .A4(n87348), .ZN(
        n87331) );
  NAND2_X1 U72923 ( .A1(n87349), .A2(n87350), .ZN(n87348) );
  AOI22_X1 U72924 ( .A1(n86477), .A2(n110880), .B1(n86478), .B2(n110884), .ZN(
        n87350) );
  AOI22_X1 U72925 ( .A1(n105697), .A2(n110879), .B1(n86480), .B2(n74317), .ZN(
        n87349) );
  NAND2_X1 U72926 ( .A1(n87351), .A2(n87352), .ZN(n87347) );
  AOI22_X1 U72927 ( .A1(n86483), .A2(n74326), .B1(n105694), .B2(n110886), .ZN(
        n87352) );
  AOI22_X1 U72928 ( .A1(n86485), .A2(n110887), .B1(n86486), .B2(n110878), .ZN(
        n87351) );
  NAND2_X1 U72929 ( .A1(n87353), .A2(n87354), .ZN(n87346) );
  AOI22_X1 U72930 ( .A1(n86489), .A2(n110885), .B1(n105690), .B2(n110889), 
        .ZN(n87354) );
  AOI22_X1 U72931 ( .A1(n86491), .A2(n74319), .B1(n86492), .B2(n110888), .ZN(
        n87353) );
  NAND2_X1 U72932 ( .A1(n87355), .A2(n87356), .ZN(n87345) );
  AOI22_X1 U72933 ( .A1(n105687), .A2(n74331), .B1(n86496), .B2(n110892), .ZN(
        n87356) );
  AOI22_X1 U72934 ( .A1(n86497), .A2(n74329), .B1(n86498), .B2(n110883), .ZN(
        n87355) );
  NAND2_X1 U72935 ( .A1(n87357), .A2(n87358), .ZN(n87275) );
  NOR4_X1 U72936 ( .A1(n87359), .A2(n87360), .A3(n87361), .A4(n87362), .ZN(
        n87358) );
  NAND2_X1 U72937 ( .A1(n87363), .A2(n87364), .ZN(n87362) );
  AOI22_X1 U72938 ( .A1(n86507), .A2(n110917), .B1(n86508), .B2(n110916), .ZN(
        n87364) );
  AOI22_X1 U72939 ( .A1(n86509), .A2(n74365), .B1(n86510), .B2(n110914), .ZN(
        n87363) );
  NAND2_X1 U72940 ( .A1(n87365), .A2(n87366), .ZN(n87361) );
  AOI22_X1 U72941 ( .A1(n86513), .A2(n110912), .B1(n105678), .B2(n110915), 
        .ZN(n87366) );
  AOI22_X1 U72942 ( .A1(n86515), .A2(n74371), .B1(n105677), .B2(n110913), .ZN(
        n87365) );
  NAND2_X1 U72943 ( .A1(n87367), .A2(n87368), .ZN(n87360) );
  AOI22_X1 U72944 ( .A1(n86519), .A2(n110923), .B1(n86520), .B2(n74377), .ZN(
        n87368) );
  AOI22_X1 U72945 ( .A1(n86521), .A2(n110921), .B1(n86522), .B2(n110922), .ZN(
        n87367) );
  NAND2_X1 U72946 ( .A1(n87369), .A2(n87370), .ZN(n87359) );
  AOI22_X1 U72947 ( .A1(n86525), .A2(n110918), .B1(n86526), .B2(n110920), .ZN(
        n87370) );
  AOI22_X1 U72948 ( .A1(n86527), .A2(n110924), .B1(n86528), .B2(n110919), .ZN(
        n87369) );
  NOR4_X1 U72949 ( .A1(n87371), .A2(n87372), .A3(n87373), .A4(n87374), .ZN(
        n87357) );
  NAND2_X1 U72950 ( .A1(n87375), .A2(n87376), .ZN(n87374) );
  AOI22_X1 U72951 ( .A1(n105675), .A2(n110899), .B1(n86536), .B2(n110902), 
        .ZN(n87376) );
  AOI22_X1 U72952 ( .A1(n86537), .A2(n110901), .B1(n86538), .B2(n74348), .ZN(
        n87375) );
  NAND2_X1 U72953 ( .A1(n87377), .A2(n87378), .ZN(n87373) );
  AOI22_X1 U72954 ( .A1(n86541), .A2(n110908), .B1(n86542), .B2(n110898), .ZN(
        n87378) );
  AOI22_X1 U72955 ( .A1(n86543), .A2(n110900), .B1(n105668), .B2(n110905), 
        .ZN(n87377) );
  NAND2_X1 U72956 ( .A1(n87379), .A2(n87380), .ZN(n87372) );
  AOI22_X1 U72957 ( .A1(n86547), .A2(n110904), .B1(n86548), .B2(n110909), .ZN(
        n87380) );
  AOI22_X1 U72958 ( .A1(n105665), .A2(n110911), .B1(n86550), .B2(n110907), 
        .ZN(n87379) );
  NAND2_X1 U72959 ( .A1(n87381), .A2(n87382), .ZN(n87371) );
  AOI22_X1 U72960 ( .A1(n86553), .A2(n74366), .B1(n86554), .B2(n110903), .ZN(
        n87382) );
  AOI22_X1 U72961 ( .A1(n105661), .A2(n110906), .B1(n86556), .B2(n110910), 
        .ZN(n87381) );
  AOI21_X1 U72962 ( .B1(n86302), .B2(n87384), .A(n87385), .ZN(n87383) );
  OAI21_X1 U72963 ( .B1(n87386), .B2(n86306), .A(n87387), .ZN(n87385) );
  OAI21_X1 U72964 ( .B1(n87388), .B2(n87389), .A(n105786), .ZN(n87387) );
  OAI21_X1 U72965 ( .B1(n110542), .B2(n86311), .A(n87390), .ZN(n87389) );
  AOI22_X1 U72966 ( .A1(n86313), .A2(n73841), .B1(n105784), .B2(n110540), .ZN(
        n87390) );
  NAND2_X1 U72967 ( .A1(n87391), .A2(n87392), .ZN(n87388) );
  AOI22_X1 U72968 ( .A1(n86317), .A2(n110538), .B1(n86318), .B2(n110543), .ZN(
        n87392) );
  AOI22_X1 U72969 ( .A1(n86319), .A2(n110541), .B1(n86320), .B2(n110539), .ZN(
        n87391) );
  NOR4_X1 U72970 ( .A1(n87393), .A2(n87394), .A3(n87395), .A4(n87396), .ZN(
        n87386) );
  NAND2_X1 U72971 ( .A1(n87397), .A2(n87398), .ZN(n87396) );
  NOR4_X1 U72972 ( .A1(n87399), .A2(n87400), .A3(n87401), .A4(n87402), .ZN(
        n87398) );
  NAND2_X1 U72973 ( .A1(n87403), .A2(n87404), .ZN(n87402) );
  AOI22_X1 U72974 ( .A1(n86333), .A2(n110519), .B1(n86334), .B2(n110520), .ZN(
        n87404) );
  AOI22_X1 U72975 ( .A1(n86335), .A2(n110528), .B1(n86336), .B2(n110526), .ZN(
        n87403) );
  NAND2_X1 U72976 ( .A1(n87405), .A2(n87406), .ZN(n87401) );
  AOI22_X1 U72977 ( .A1(n86339), .A2(n73710), .B1(n86340), .B2(n110523), .ZN(
        n87406) );
  AOI22_X1 U72978 ( .A1(n86341), .A2(n73814), .B1(n86342), .B2(n110448), .ZN(
        n87405) );
  NAND2_X1 U72979 ( .A1(n87407), .A2(n87408), .ZN(n87400) );
  AOI22_X1 U72980 ( .A1(n86345), .A2(n110452), .B1(n86346), .B2(n73714), .ZN(
        n87408) );
  AOI22_X1 U72981 ( .A1(n86347), .A2(n110524), .B1(n86348), .B2(n110521), .ZN(
        n87407) );
  NAND2_X1 U72982 ( .A1(n87409), .A2(n87410), .ZN(n87399) );
  AOI22_X1 U72983 ( .A1(n86351), .A2(n110450), .B1(n86352), .B2(n110454), .ZN(
        n87410) );
  AOI22_X1 U72984 ( .A1(n86353), .A2(n110453), .B1(n86354), .B2(n73716), .ZN(
        n87409) );
  NOR4_X1 U72985 ( .A1(n87411), .A2(n87412), .A3(n87413), .A4(n87414), .ZN(
        n87397) );
  NAND2_X1 U72986 ( .A1(n87415), .A2(n87416), .ZN(n87414) );
  AOI22_X1 U72987 ( .A1(n86361), .A2(n110529), .B1(n86362), .B2(n110532), .ZN(
        n87416) );
  AOI22_X1 U72988 ( .A1(n86363), .A2(n110533), .B1(n105760), .B2(n110535), 
        .ZN(n87415) );
  NAND2_X1 U72989 ( .A1(n87417), .A2(n87418), .ZN(n87413) );
  AOI22_X1 U72990 ( .A1(n86367), .A2(n110534), .B1(n86368), .B2(n110530), .ZN(
        n87418) );
  AOI22_X1 U72991 ( .A1(n86369), .A2(n110536), .B1(n86370), .B2(n110531), .ZN(
        n87417) );
  NAND2_X1 U72992 ( .A1(n87419), .A2(n87420), .ZN(n87412) );
  AOI22_X1 U72993 ( .A1(n86373), .A2(n73824), .B1(n86374), .B2(n73823), .ZN(
        n87420) );
  AOI22_X1 U72994 ( .A1(n86375), .A2(n73826), .B1(n86376), .B2(n110537), .ZN(
        n87419) );
  NAND2_X1 U72995 ( .A1(n87421), .A2(n87422), .ZN(n87411) );
  AOI22_X1 U72996 ( .A1(n86379), .A2(n110522), .B1(n86380), .B2(n110527), .ZN(
        n87422) );
  AOI22_X1 U72997 ( .A1(n86381), .A2(n73821), .B1(n105748), .B2(n110525), .ZN(
        n87421) );
  NAND2_X1 U72998 ( .A1(n87423), .A2(n87424), .ZN(n87395) );
  NOR4_X1 U72999 ( .A1(n87425), .A2(n87426), .A3(n87427), .A4(n87428), .ZN(
        n87424) );
  NAND2_X1 U73000 ( .A1(n87429), .A2(n87430), .ZN(n87428) );
  AOI22_X1 U73001 ( .A1(n86391), .A2(n110463), .B1(n86392), .B2(n110465), .ZN(
        n87430) );
  AOI22_X1 U73002 ( .A1(n86393), .A2(n73739), .B1(n86394), .B2(n110464), .ZN(
        n87429) );
  NAND2_X1 U73003 ( .A1(n87431), .A2(n87432), .ZN(n87427) );
  AOI22_X1 U73004 ( .A1(n86397), .A2(n73743), .B1(n86398), .B2(n73745), .ZN(
        n87432) );
  AOI22_X1 U73005 ( .A1(n86399), .A2(n110470), .B1(n86400), .B2(n110471), .ZN(
        n87431) );
  NAND2_X1 U73006 ( .A1(n87433), .A2(n87434), .ZN(n87426) );
  AOI22_X1 U73007 ( .A1(n86403), .A2(n110468), .B1(n86404), .B2(n110469), .ZN(
        n87434) );
  AOI22_X1 U73008 ( .A1(n86405), .A2(n73744), .B1(n105736), .B2(n73738), .ZN(
        n87433) );
  NAND2_X1 U73009 ( .A1(n87435), .A2(n87436), .ZN(n87425) );
  AOI22_X1 U73010 ( .A1(n86409), .A2(n110476), .B1(n86410), .B2(n73750), .ZN(
        n87436) );
  AOI22_X1 U73011 ( .A1(n86411), .A2(n110475), .B1(n86412), .B2(n73748), .ZN(
        n87435) );
  NOR4_X1 U73012 ( .A1(n87437), .A2(n87438), .A3(n87439), .A4(n87440), .ZN(
        n87423) );
  NAND2_X1 U73013 ( .A1(n87441), .A2(n87442), .ZN(n87440) );
  AOI22_X1 U73014 ( .A1(n86419), .A2(n110458), .B1(n86420), .B2(n110449), .ZN(
        n87442) );
  AOI22_X1 U73015 ( .A1(n86421), .A2(n110451), .B1(n86422), .B2(n73722), .ZN(
        n87441) );
  NAND2_X1 U73016 ( .A1(n87443), .A2(n87444), .ZN(n87439) );
  AOI22_X1 U73017 ( .A1(n86425), .A2(n110456), .B1(n86426), .B2(n110460), .ZN(
        n87444) );
  AOI22_X1 U73018 ( .A1(n105725), .A2(n110462), .B1(n86428), .B2(n110459), 
        .ZN(n87443) );
  NAND2_X1 U73019 ( .A1(n87445), .A2(n87446), .ZN(n87438) );
  AOI22_X1 U73020 ( .A1(n86431), .A2(n73731), .B1(n86432), .B2(n110455), .ZN(
        n87446) );
  AOI22_X1 U73021 ( .A1(n86433), .A2(n110457), .B1(n86434), .B2(n110461), .ZN(
        n87445) );
  NAND2_X1 U73022 ( .A1(n87447), .A2(n87448), .ZN(n87437) );
  AOI22_X1 U73023 ( .A1(n86437), .A2(n110467), .B1(n86438), .B2(n73735), .ZN(
        n87448) );
  AOI22_X1 U73024 ( .A1(n86439), .A2(n73733), .B1(n105716), .B2(n110466), .ZN(
        n87447) );
  NAND2_X1 U73025 ( .A1(n87449), .A2(n87450), .ZN(n87394) );
  NOR4_X1 U73026 ( .A1(n87451), .A2(n87452), .A3(n87453), .A4(n87454), .ZN(
        n87450) );
  NAND2_X1 U73027 ( .A1(n87455), .A2(n87456), .ZN(n87454) );
  AOI22_X1 U73028 ( .A1(n86449), .A2(n73773), .B1(n86450), .B2(n110485), .ZN(
        n87456) );
  AOI22_X1 U73029 ( .A1(n86451), .A2(n110488), .B1(n86452), .B2(n110487), .ZN(
        n87455) );
  NAND2_X1 U73030 ( .A1(n87457), .A2(n87458), .ZN(n87453) );
  AOI22_X1 U73031 ( .A1(n105711), .A2(n110492), .B1(n86456), .B2(n110491), 
        .ZN(n87458) );
  AOI22_X1 U73032 ( .A1(n105709), .A2(n110484), .B1(n105708), .B2(n111017), 
        .ZN(n87457) );
  NAND2_X1 U73033 ( .A1(n87459), .A2(n87460), .ZN(n87452) );
  AOI22_X1 U73034 ( .A1(n86461), .A2(n110493), .B1(n86462), .B2(n73772), .ZN(
        n87460) );
  AOI22_X1 U73035 ( .A1(n86463), .A2(n73777), .B1(n86464), .B2(n73779), .ZN(
        n87459) );
  NAND2_X1 U73036 ( .A1(n87461), .A2(n87462), .ZN(n87451) );
  AOI22_X1 U73037 ( .A1(n86467), .A2(n111036), .B1(n86468), .B2(n73785), .ZN(
        n87462) );
  AOI22_X1 U73038 ( .A1(n86469), .A2(n110489), .B1(n86470), .B2(n110490), .ZN(
        n87461) );
  NOR4_X1 U73039 ( .A1(n87463), .A2(n87464), .A3(n87465), .A4(n87466), .ZN(
        n87449) );
  NAND2_X1 U73040 ( .A1(n87467), .A2(n87468), .ZN(n87466) );
  AOI22_X1 U73041 ( .A1(n86477), .A2(n110474), .B1(n86478), .B2(n110479), .ZN(
        n87468) );
  AOI22_X1 U73042 ( .A1(n105697), .A2(n110473), .B1(n86480), .B2(n73753), .ZN(
        n87467) );
  NAND2_X1 U73043 ( .A1(n87469), .A2(n87470), .ZN(n87465) );
  AOI22_X1 U73044 ( .A1(n86483), .A2(n73762), .B1(n105694), .B2(n110480), .ZN(
        n87470) );
  AOI22_X1 U73045 ( .A1(n86485), .A2(n110481), .B1(n86486), .B2(n110472), .ZN(
        n87469) );
  NAND2_X1 U73046 ( .A1(n87471), .A2(n87472), .ZN(n87464) );
  AOI22_X1 U73047 ( .A1(n86489), .A2(n73757), .B1(n86490), .B2(n110483), .ZN(
        n87472) );
  AOI22_X1 U73048 ( .A1(n86491), .A2(n110478), .B1(n86492), .B2(n110482), .ZN(
        n87471) );
  NAND2_X1 U73049 ( .A1(n87473), .A2(n87474), .ZN(n87463) );
  AOI22_X1 U73050 ( .A1(n105687), .A2(n73767), .B1(n86496), .B2(n110486), .ZN(
        n87474) );
  AOI22_X1 U73051 ( .A1(n86497), .A2(n73765), .B1(n86498), .B2(n110477), .ZN(
        n87473) );
  NAND2_X1 U73052 ( .A1(n87475), .A2(n87476), .ZN(n87393) );
  NOR4_X1 U73053 ( .A1(n87477), .A2(n87478), .A3(n87479), .A4(n87480), .ZN(
        n87476) );
  NAND2_X1 U73054 ( .A1(n87481), .A2(n87482), .ZN(n87480) );
  AOI22_X1 U73055 ( .A1(n86507), .A2(n110512), .B1(n86508), .B2(n110511), .ZN(
        n87482) );
  AOI22_X1 U73056 ( .A1(n86509), .A2(n73801), .B1(n86510), .B2(n110509), .ZN(
        n87481) );
  NAND2_X1 U73057 ( .A1(n87483), .A2(n87484), .ZN(n87479) );
  AOI22_X1 U73058 ( .A1(n86513), .A2(n110507), .B1(n105678), .B2(n110510), 
        .ZN(n87484) );
  AOI22_X1 U73059 ( .A1(n86515), .A2(n73807), .B1(n86516), .B2(n110508), .ZN(
        n87483) );
  NAND2_X1 U73060 ( .A1(n87485), .A2(n87486), .ZN(n87478) );
  AOI22_X1 U73061 ( .A1(n86519), .A2(n110517), .B1(n86520), .B2(n73813), .ZN(
        n87486) );
  AOI22_X1 U73062 ( .A1(n86521), .A2(n110515), .B1(n86522), .B2(n110516), .ZN(
        n87485) );
  NAND2_X1 U73063 ( .A1(n87487), .A2(n87488), .ZN(n87477) );
  AOI22_X1 U73064 ( .A1(n86525), .A2(n73805), .B1(n86526), .B2(n110514), .ZN(
        n87488) );
  AOI22_X1 U73065 ( .A1(n86527), .A2(n73812), .B1(n86528), .B2(n110513), .ZN(
        n87487) );
  NOR4_X1 U73066 ( .A1(n87489), .A2(n87490), .A3(n87491), .A4(n87492), .ZN(
        n87475) );
  NAND2_X1 U73067 ( .A1(n87493), .A2(n87494), .ZN(n87492) );
  AOI22_X1 U73068 ( .A1(n105675), .A2(n110494), .B1(n86536), .B2(n110497), 
        .ZN(n87494) );
  AOI22_X1 U73069 ( .A1(n86537), .A2(n110496), .B1(n86538), .B2(n73784), .ZN(
        n87493) );
  NAND2_X1 U73070 ( .A1(n87495), .A2(n87496), .ZN(n87491) );
  AOI22_X1 U73071 ( .A1(n86541), .A2(n110503), .B1(n86542), .B2(n73780), .ZN(
        n87496) );
  AOI22_X1 U73072 ( .A1(n86543), .A2(n110495), .B1(n105668), .B2(n110500), 
        .ZN(n87495) );
  NAND2_X1 U73073 ( .A1(n87497), .A2(n87498), .ZN(n87490) );
  AOI22_X1 U73074 ( .A1(n86547), .A2(n110499), .B1(n86548), .B2(n110504), .ZN(
        n87498) );
  AOI22_X1 U73075 ( .A1(n86549), .A2(n110506), .B1(n86550), .B2(n110502), .ZN(
        n87497) );
  NAND2_X1 U73076 ( .A1(n87499), .A2(n87500), .ZN(n87489) );
  AOI22_X1 U73077 ( .A1(n86553), .A2(n73802), .B1(n86554), .B2(n110498), .ZN(
        n87500) );
  AOI22_X1 U73078 ( .A1(n105661), .A2(n110501), .B1(n105660), .B2(n110505), 
        .ZN(n87499) );
  AOI21_X1 U73079 ( .B1(n86302), .B2(n87502), .A(n87503), .ZN(n87501) );
  OAI21_X1 U73080 ( .B1(n87504), .B2(n86306), .A(n87505), .ZN(n87503) );
  OAI21_X1 U73081 ( .B1(n87506), .B2(n87507), .A(n86310), .ZN(n87505) );
  OAI21_X1 U73082 ( .B1(n110327), .B2(n86311), .A(n87508), .ZN(n87507) );
  AOI22_X1 U73083 ( .A1(n86313), .A2(n73545), .B1(n105784), .B2(n110325), .ZN(
        n87508) );
  NAND2_X1 U73084 ( .A1(n87509), .A2(n87510), .ZN(n87506) );
  AOI22_X1 U73085 ( .A1(n86317), .A2(n110323), .B1(n86318), .B2(n110328), .ZN(
        n87510) );
  AOI22_X1 U73086 ( .A1(n86319), .A2(n110326), .B1(n86320), .B2(n110324), .ZN(
        n87509) );
  NOR4_X1 U73087 ( .A1(n87511), .A2(n87512), .A3(n87513), .A4(n87514), .ZN(
        n87504) );
  NAND2_X1 U73088 ( .A1(n87515), .A2(n87516), .ZN(n87514) );
  NOR4_X1 U73089 ( .A1(n87517), .A2(n87518), .A3(n87519), .A4(n87520), .ZN(
        n87516) );
  NAND2_X1 U73090 ( .A1(n87521), .A2(n87522), .ZN(n87520) );
  AOI22_X1 U73091 ( .A1(n86333), .A2(n110304), .B1(n86334), .B2(n110305), .ZN(
        n87522) );
  AOI22_X1 U73092 ( .A1(n86335), .A2(n110313), .B1(n86336), .B2(n110311), .ZN(
        n87521) );
  NAND2_X1 U73093 ( .A1(n87523), .A2(n87524), .ZN(n87519) );
  AOI22_X1 U73094 ( .A1(n86339), .A2(n73414), .B1(n86340), .B2(n110308), .ZN(
        n87524) );
  AOI22_X1 U73095 ( .A1(n86341), .A2(n73518), .B1(n86342), .B2(n110231), .ZN(
        n87523) );
  NAND2_X1 U73096 ( .A1(n87525), .A2(n87526), .ZN(n87518) );
  AOI22_X1 U73097 ( .A1(n86345), .A2(n110234), .B1(n86346), .B2(n73418), .ZN(
        n87526) );
  AOI22_X1 U73098 ( .A1(n86347), .A2(n110309), .B1(n86348), .B2(n110306), .ZN(
        n87525) );
  NAND2_X1 U73099 ( .A1(n87527), .A2(n87528), .ZN(n87517) );
  AOI22_X1 U73100 ( .A1(n86351), .A2(n110232), .B1(n86352), .B2(n110236), .ZN(
        n87528) );
  AOI22_X1 U73101 ( .A1(n86353), .A2(n110235), .B1(n86354), .B2(n73420), .ZN(
        n87527) );
  NOR4_X1 U73102 ( .A1(n87529), .A2(n87530), .A3(n87531), .A4(n87532), .ZN(
        n87515) );
  NAND2_X1 U73103 ( .A1(n87533), .A2(n87534), .ZN(n87532) );
  AOI22_X1 U73104 ( .A1(n86361), .A2(n110314), .B1(n86362), .B2(n110317), .ZN(
        n87534) );
  AOI22_X1 U73105 ( .A1(n86363), .A2(n110318), .B1(n105760), .B2(n110320), 
        .ZN(n87533) );
  NAND2_X1 U73106 ( .A1(n87535), .A2(n87536), .ZN(n87531) );
  AOI22_X1 U73107 ( .A1(n86367), .A2(n110319), .B1(n86368), .B2(n110315), .ZN(
        n87536) );
  AOI22_X1 U73108 ( .A1(n86369), .A2(n110321), .B1(n86370), .B2(n110316), .ZN(
        n87535) );
  NAND2_X1 U73109 ( .A1(n87537), .A2(n87538), .ZN(n87530) );
  AOI22_X1 U73110 ( .A1(n86373), .A2(n73528), .B1(n86374), .B2(n73527), .ZN(
        n87538) );
  AOI22_X1 U73111 ( .A1(n86375), .A2(n73530), .B1(n86376), .B2(n110322), .ZN(
        n87537) );
  NAND2_X1 U73112 ( .A1(n87539), .A2(n87540), .ZN(n87529) );
  AOI22_X1 U73113 ( .A1(n86379), .A2(n110307), .B1(n86380), .B2(n110312), .ZN(
        n87540) );
  AOI22_X1 U73114 ( .A1(n86381), .A2(n73525), .B1(n105748), .B2(n110310), .ZN(
        n87539) );
  NAND2_X1 U73115 ( .A1(n87541), .A2(n87542), .ZN(n87513) );
  NOR4_X1 U73116 ( .A1(n87543), .A2(n87544), .A3(n87545), .A4(n87546), .ZN(
        n87542) );
  NAND2_X1 U73117 ( .A1(n87547), .A2(n87548), .ZN(n87546) );
  AOI22_X1 U73118 ( .A1(n86391), .A2(n110245), .B1(n86392), .B2(n110247), .ZN(
        n87548) );
  AOI22_X1 U73119 ( .A1(n86393), .A2(n73443), .B1(n86394), .B2(n110246), .ZN(
        n87547) );
  NAND2_X1 U73120 ( .A1(n87549), .A2(n87550), .ZN(n87545) );
  AOI22_X1 U73121 ( .A1(n86397), .A2(n73447), .B1(n86398), .B2(n73449), .ZN(
        n87550) );
  AOI22_X1 U73122 ( .A1(n86399), .A2(n110252), .B1(n86400), .B2(n110253), .ZN(
        n87549) );
  NAND2_X1 U73123 ( .A1(n87551), .A2(n87552), .ZN(n87544) );
  AOI22_X1 U73124 ( .A1(n86403), .A2(n110250), .B1(n86404), .B2(n110251), .ZN(
        n87552) );
  AOI22_X1 U73125 ( .A1(n86405), .A2(n73448), .B1(n105736), .B2(n73442), .ZN(
        n87551) );
  NAND2_X1 U73126 ( .A1(n87553), .A2(n87554), .ZN(n87543) );
  AOI22_X1 U73127 ( .A1(n86409), .A2(n110258), .B1(n86410), .B2(n73454), .ZN(
        n87554) );
  AOI22_X1 U73128 ( .A1(n86411), .A2(n110257), .B1(n86412), .B2(n73452), .ZN(
        n87553) );
  NOR4_X1 U73129 ( .A1(n87555), .A2(n87556), .A3(n87557), .A4(n87558), .ZN(
        n87541) );
  NAND2_X1 U73130 ( .A1(n87559), .A2(n87560), .ZN(n87558) );
  AOI22_X1 U73131 ( .A1(n86419), .A2(n110240), .B1(n86420), .B2(n111020), .ZN(
        n87560) );
  AOI22_X1 U73132 ( .A1(n86421), .A2(n110233), .B1(n86422), .B2(n73426), .ZN(
        n87559) );
  NAND2_X1 U73133 ( .A1(n87561), .A2(n87562), .ZN(n87557) );
  AOI22_X1 U73134 ( .A1(n86425), .A2(n110238), .B1(n86426), .B2(n110242), .ZN(
        n87562) );
  AOI22_X1 U73135 ( .A1(n105725), .A2(n110244), .B1(n86428), .B2(n110241), 
        .ZN(n87561) );
  NAND2_X1 U73136 ( .A1(n87563), .A2(n87564), .ZN(n87556) );
  AOI22_X1 U73137 ( .A1(n86431), .A2(n73435), .B1(n86432), .B2(n110237), .ZN(
        n87564) );
  AOI22_X1 U73138 ( .A1(n86433), .A2(n110239), .B1(n86434), .B2(n110243), .ZN(
        n87563) );
  NAND2_X1 U73139 ( .A1(n87565), .A2(n87566), .ZN(n87555) );
  AOI22_X1 U73140 ( .A1(n86437), .A2(n110249), .B1(n86438), .B2(n73439), .ZN(
        n87566) );
  AOI22_X1 U73141 ( .A1(n86439), .A2(n73437), .B1(n105716), .B2(n110248), .ZN(
        n87565) );
  NAND2_X1 U73142 ( .A1(n87567), .A2(n87568), .ZN(n87512) );
  NOR4_X1 U73143 ( .A1(n87569), .A2(n87570), .A3(n87571), .A4(n87572), .ZN(
        n87568) );
  NAND2_X1 U73144 ( .A1(n87573), .A2(n87574), .ZN(n87572) );
  AOI22_X1 U73145 ( .A1(n86449), .A2(n73477), .B1(n86450), .B2(n110267), .ZN(
        n87574) );
  AOI22_X1 U73146 ( .A1(n86451), .A2(n110271), .B1(n86452), .B2(n110270), .ZN(
        n87573) );
  NAND2_X1 U73147 ( .A1(n87575), .A2(n87576), .ZN(n87571) );
  AOI22_X1 U73148 ( .A1(n105711), .A2(n110275), .B1(n86456), .B2(n110274), 
        .ZN(n87576) );
  AOI22_X1 U73149 ( .A1(n105709), .A2(n110266), .B1(n86458), .B2(n110268), 
        .ZN(n87575) );
  NAND2_X1 U73150 ( .A1(n87577), .A2(n87578), .ZN(n87570) );
  AOI22_X1 U73151 ( .A1(n86461), .A2(n110276), .B1(n86462), .B2(n73476), .ZN(
        n87578) );
  AOI22_X1 U73152 ( .A1(n86463), .A2(n73481), .B1(n86464), .B2(n73483), .ZN(
        n87577) );
  NAND2_X1 U73153 ( .A1(n87579), .A2(n87580), .ZN(n87569) );
  AOI22_X1 U73154 ( .A1(n86467), .A2(n110278), .B1(n86468), .B2(n73489), .ZN(
        n87580) );
  AOI22_X1 U73155 ( .A1(n86469), .A2(n110272), .B1(n86470), .B2(n110273), .ZN(
        n87579) );
  NOR4_X1 U73156 ( .A1(n87581), .A2(n87582), .A3(n87583), .A4(n87584), .ZN(
        n87567) );
  NAND2_X1 U73157 ( .A1(n87585), .A2(n87586), .ZN(n87584) );
  AOI22_X1 U73158 ( .A1(n86477), .A2(n110256), .B1(n86478), .B2(n110261), .ZN(
        n87586) );
  AOI22_X1 U73159 ( .A1(n105697), .A2(n110255), .B1(n86480), .B2(n73457), .ZN(
        n87585) );
  NAND2_X1 U73160 ( .A1(n87587), .A2(n87588), .ZN(n87583) );
  AOI22_X1 U73161 ( .A1(n86483), .A2(n73466), .B1(n105694), .B2(n110262), .ZN(
        n87588) );
  AOI22_X1 U73162 ( .A1(n86485), .A2(n110263), .B1(n86486), .B2(n110254), .ZN(
        n87587) );
  NAND2_X1 U73163 ( .A1(n87589), .A2(n87590), .ZN(n87582) );
  AOI22_X1 U73164 ( .A1(n86489), .A2(n73461), .B1(n86490), .B2(n110265), .ZN(
        n87590) );
  AOI22_X1 U73165 ( .A1(n86491), .A2(n110260), .B1(n86492), .B2(n110264), .ZN(
        n87589) );
  NAND2_X1 U73166 ( .A1(n87591), .A2(n87592), .ZN(n87581) );
  AOI22_X1 U73167 ( .A1(n105687), .A2(n73471), .B1(n86496), .B2(n110269), .ZN(
        n87592) );
  AOI22_X1 U73168 ( .A1(n86497), .A2(n73469), .B1(n86498), .B2(n110259), .ZN(
        n87591) );
  NAND2_X1 U73169 ( .A1(n87593), .A2(n87594), .ZN(n87511) );
  NOR4_X1 U73170 ( .A1(n87595), .A2(n87596), .A3(n87597), .A4(n87598), .ZN(
        n87594) );
  NAND2_X1 U73171 ( .A1(n87599), .A2(n87600), .ZN(n87598) );
  AOI22_X1 U73172 ( .A1(n86507), .A2(n110295), .B1(n86508), .B2(n110294), .ZN(
        n87600) );
  AOI22_X1 U73173 ( .A1(n86509), .A2(n73505), .B1(n86510), .B2(n110292), .ZN(
        n87599) );
  NAND2_X1 U73174 ( .A1(n87601), .A2(n87602), .ZN(n87597) );
  AOI22_X1 U73175 ( .A1(n86513), .A2(n110290), .B1(n105678), .B2(n110293), 
        .ZN(n87602) );
  AOI22_X1 U73176 ( .A1(n86515), .A2(n73511), .B1(n86516), .B2(n110291), .ZN(
        n87601) );
  NAND2_X1 U73177 ( .A1(n87603), .A2(n87604), .ZN(n87596) );
  AOI22_X1 U73178 ( .A1(n86519), .A2(n110301), .B1(n86520), .B2(n73517), .ZN(
        n87604) );
  AOI22_X1 U73179 ( .A1(n86521), .A2(n110299), .B1(n86522), .B2(n110300), .ZN(
        n87603) );
  NAND2_X1 U73180 ( .A1(n87605), .A2(n87606), .ZN(n87595) );
  AOI22_X1 U73181 ( .A1(n86525), .A2(n110296), .B1(n86526), .B2(n110298), .ZN(
        n87606) );
  AOI22_X1 U73182 ( .A1(n86527), .A2(n110302), .B1(n86528), .B2(n110297), .ZN(
        n87605) );
  NOR4_X1 U73183 ( .A1(n87607), .A2(n87608), .A3(n87609), .A4(n87610), .ZN(
        n87593) );
  NAND2_X1 U73184 ( .A1(n87611), .A2(n87612), .ZN(n87610) );
  AOI22_X1 U73185 ( .A1(n105675), .A2(n110277), .B1(n86536), .B2(n110280), 
        .ZN(n87612) );
  AOI22_X1 U73186 ( .A1(n86537), .A2(n111039), .B1(n86538), .B2(n73488), .ZN(
        n87611) );
  NAND2_X1 U73187 ( .A1(n87613), .A2(n87614), .ZN(n87609) );
  AOI22_X1 U73188 ( .A1(n86541), .A2(n110286), .B1(n86542), .B2(n73484), .ZN(
        n87614) );
  AOI22_X1 U73189 ( .A1(n86543), .A2(n110279), .B1(n105668), .B2(n110283), 
        .ZN(n87613) );
  NAND2_X1 U73190 ( .A1(n87615), .A2(n87616), .ZN(n87608) );
  AOI22_X1 U73191 ( .A1(n86547), .A2(n110282), .B1(n86548), .B2(n110287), .ZN(
        n87616) );
  AOI22_X1 U73192 ( .A1(n86549), .A2(n110289), .B1(n105664), .B2(n110285), 
        .ZN(n87615) );
  NAND2_X1 U73193 ( .A1(n87617), .A2(n87618), .ZN(n87607) );
  AOI22_X1 U73194 ( .A1(n86553), .A2(n73506), .B1(n86554), .B2(n110281), .ZN(
        n87618) );
  AOI22_X1 U73195 ( .A1(n105661), .A2(n110284), .B1(n105660), .B2(n110288), 
        .ZN(n87617) );
  AOI21_X1 U73196 ( .B1(n86302), .B2(n87620), .A(n87621), .ZN(n87619) );
  OAI21_X1 U73197 ( .B1(n87622), .B2(n86306), .A(n87623), .ZN(n87621) );
  OAI21_X1 U73198 ( .B1(n87624), .B2(n87625), .A(n86310), .ZN(n87623) );
  OAI21_X1 U73199 ( .B1(n110647), .B2(n86311), .A(n87626), .ZN(n87625) );
  AOI22_X1 U73200 ( .A1(n86313), .A2(n73982), .B1(n105784), .B2(n110645), .ZN(
        n87626) );
  NAND2_X1 U73201 ( .A1(n87627), .A2(n87628), .ZN(n87624) );
  AOI22_X1 U73202 ( .A1(n86317), .A2(n110643), .B1(n86318), .B2(n110648), .ZN(
        n87628) );
  AOI22_X1 U73203 ( .A1(n86319), .A2(n110646), .B1(n86320), .B2(n110644), .ZN(
        n87627) );
  NOR4_X1 U73204 ( .A1(n87629), .A2(n87630), .A3(n87631), .A4(n87632), .ZN(
        n87622) );
  NAND2_X1 U73205 ( .A1(n87633), .A2(n87634), .ZN(n87632) );
  NOR4_X1 U73206 ( .A1(n87635), .A2(n87636), .A3(n87637), .A4(n87638), .ZN(
        n87634) );
  NAND2_X1 U73207 ( .A1(n87639), .A2(n87640), .ZN(n87638) );
  AOI22_X1 U73208 ( .A1(n86333), .A2(n110624), .B1(n86334), .B2(n110625), .ZN(
        n87640) );
  AOI22_X1 U73209 ( .A1(n86335), .A2(n110633), .B1(n86336), .B2(n110631), .ZN(
        n87639) );
  NAND2_X1 U73210 ( .A1(n87641), .A2(n87642), .ZN(n87637) );
  AOI22_X1 U73211 ( .A1(n86339), .A2(n73851), .B1(n86340), .B2(n110628), .ZN(
        n87642) );
  AOI22_X1 U73212 ( .A1(n86341), .A2(n73955), .B1(n86342), .B2(n110548), .ZN(
        n87641) );
  NAND2_X1 U73213 ( .A1(n87643), .A2(n87644), .ZN(n87636) );
  AOI22_X1 U73214 ( .A1(n86345), .A2(n110551), .B1(n86346), .B2(n73855), .ZN(
        n87644) );
  AOI22_X1 U73215 ( .A1(n86347), .A2(n110629), .B1(n86348), .B2(n110626), .ZN(
        n87643) );
  NAND2_X1 U73216 ( .A1(n87645), .A2(n87646), .ZN(n87635) );
  AOI22_X1 U73217 ( .A1(n86351), .A2(n110549), .B1(n86352), .B2(n110553), .ZN(
        n87646) );
  AOI22_X1 U73218 ( .A1(n86353), .A2(n110552), .B1(n86354), .B2(n73857), .ZN(
        n87645) );
  NOR4_X1 U73219 ( .A1(n87647), .A2(n87648), .A3(n87649), .A4(n87650), .ZN(
        n87633) );
  NAND2_X1 U73220 ( .A1(n87651), .A2(n87652), .ZN(n87650) );
  AOI22_X1 U73221 ( .A1(n86361), .A2(n110634), .B1(n86362), .B2(n110637), .ZN(
        n87652) );
  AOI22_X1 U73222 ( .A1(n86363), .A2(n110638), .B1(n105760), .B2(n110640), 
        .ZN(n87651) );
  NAND2_X1 U73223 ( .A1(n87653), .A2(n87654), .ZN(n87649) );
  AOI22_X1 U73224 ( .A1(n86367), .A2(n110639), .B1(n86368), .B2(n110635), .ZN(
        n87654) );
  AOI22_X1 U73225 ( .A1(n86369), .A2(n110641), .B1(n86370), .B2(n110636), .ZN(
        n87653) );
  NAND2_X1 U73226 ( .A1(n87655), .A2(n87656), .ZN(n87648) );
  AOI22_X1 U73227 ( .A1(n86373), .A2(n73965), .B1(n86374), .B2(n73964), .ZN(
        n87656) );
  AOI22_X1 U73228 ( .A1(n86375), .A2(n73967), .B1(n86376), .B2(n110642), .ZN(
        n87655) );
  NAND2_X1 U73229 ( .A1(n87657), .A2(n87658), .ZN(n87647) );
  AOI22_X1 U73230 ( .A1(n86379), .A2(n110627), .B1(n86380), .B2(n110632), .ZN(
        n87658) );
  AOI22_X1 U73231 ( .A1(n86381), .A2(n73962), .B1(n105748), .B2(n110630), .ZN(
        n87657) );
  NAND2_X1 U73232 ( .A1(n87659), .A2(n87660), .ZN(n87631) );
  NOR4_X1 U73233 ( .A1(n87661), .A2(n87662), .A3(n87663), .A4(n87664), .ZN(
        n87660) );
  NAND2_X1 U73234 ( .A1(n87665), .A2(n87666), .ZN(n87664) );
  AOI22_X1 U73235 ( .A1(n86391), .A2(n110562), .B1(n86392), .B2(n110564), .ZN(
        n87666) );
  AOI22_X1 U73236 ( .A1(n86393), .A2(n73880), .B1(n86394), .B2(n110563), .ZN(
        n87665) );
  NAND2_X1 U73237 ( .A1(n87667), .A2(n87668), .ZN(n87663) );
  AOI22_X1 U73238 ( .A1(n86397), .A2(n73884), .B1(n86398), .B2(n73886), .ZN(
        n87668) );
  AOI22_X1 U73239 ( .A1(n86399), .A2(n110569), .B1(n86400), .B2(n110570), .ZN(
        n87667) );
  NAND2_X1 U73240 ( .A1(n87669), .A2(n87670), .ZN(n87662) );
  AOI22_X1 U73241 ( .A1(n86403), .A2(n110567), .B1(n86404), .B2(n110568), .ZN(
        n87670) );
  AOI22_X1 U73242 ( .A1(n86405), .A2(n73885), .B1(n105736), .B2(n73879), .ZN(
        n87669) );
  NAND2_X1 U73243 ( .A1(n87671), .A2(n87672), .ZN(n87661) );
  AOI22_X1 U73244 ( .A1(n86409), .A2(n110575), .B1(n86410), .B2(n73891), .ZN(
        n87672) );
  AOI22_X1 U73245 ( .A1(n86411), .A2(n110574), .B1(n86412), .B2(n73889), .ZN(
        n87671) );
  NOR4_X1 U73246 ( .A1(n87673), .A2(n87674), .A3(n87675), .A4(n87676), .ZN(
        n87659) );
  NAND2_X1 U73247 ( .A1(n87677), .A2(n87678), .ZN(n87676) );
  AOI22_X1 U73248 ( .A1(n86419), .A2(n110557), .B1(n86420), .B2(n111018), .ZN(
        n87678) );
  AOI22_X1 U73249 ( .A1(n86421), .A2(n110550), .B1(n86422), .B2(n73863), .ZN(
        n87677) );
  NAND2_X1 U73250 ( .A1(n87679), .A2(n87680), .ZN(n87675) );
  AOI22_X1 U73251 ( .A1(n86425), .A2(n110555), .B1(n86426), .B2(n110559), .ZN(
        n87680) );
  AOI22_X1 U73252 ( .A1(n105725), .A2(n110561), .B1(n86428), .B2(n110558), 
        .ZN(n87679) );
  NAND2_X1 U73253 ( .A1(n87681), .A2(n87682), .ZN(n87674) );
  AOI22_X1 U73254 ( .A1(n86431), .A2(n73872), .B1(n86432), .B2(n110554), .ZN(
        n87682) );
  AOI22_X1 U73255 ( .A1(n86433), .A2(n110556), .B1(n86434), .B2(n110560), .ZN(
        n87681) );
  NAND2_X1 U73256 ( .A1(n87683), .A2(n87684), .ZN(n87673) );
  AOI22_X1 U73257 ( .A1(n86437), .A2(n110566), .B1(n86438), .B2(n73876), .ZN(
        n87684) );
  AOI22_X1 U73258 ( .A1(n86439), .A2(n73874), .B1(n105716), .B2(n110565), .ZN(
        n87683) );
  NAND2_X1 U73259 ( .A1(n87685), .A2(n87686), .ZN(n87630) );
  NOR4_X1 U73260 ( .A1(n87687), .A2(n87688), .A3(n87689), .A4(n87690), .ZN(
        n87686) );
  NAND2_X1 U73261 ( .A1(n87691), .A2(n87692), .ZN(n87690) );
  AOI22_X1 U73262 ( .A1(n86449), .A2(n73914), .B1(n86450), .B2(n110585), .ZN(
        n87692) );
  AOI22_X1 U73263 ( .A1(n86451), .A2(n110589), .B1(n86452), .B2(n110588), .ZN(
        n87691) );
  NAND2_X1 U73264 ( .A1(n87693), .A2(n87694), .ZN(n87689) );
  AOI22_X1 U73265 ( .A1(n105711), .A2(n110593), .B1(n86456), .B2(n110592), 
        .ZN(n87694) );
  AOI22_X1 U73266 ( .A1(n105709), .A2(n110584), .B1(n105708), .B2(n110586), 
        .ZN(n87693) );
  NAND2_X1 U73267 ( .A1(n87695), .A2(n87696), .ZN(n87688) );
  AOI22_X1 U73268 ( .A1(n86461), .A2(n110594), .B1(n86462), .B2(n73913), .ZN(
        n87696) );
  AOI22_X1 U73269 ( .A1(n86463), .A2(n73918), .B1(n86464), .B2(n73920), .ZN(
        n87695) );
  NAND2_X1 U73270 ( .A1(n87697), .A2(n87698), .ZN(n87687) );
  AOI22_X1 U73271 ( .A1(n86467), .A2(n110597), .B1(n86468), .B2(n73926), .ZN(
        n87698) );
  AOI22_X1 U73272 ( .A1(n86469), .A2(n110590), .B1(n86470), .B2(n110591), .ZN(
        n87697) );
  NOR4_X1 U73273 ( .A1(n87699), .A2(n87700), .A3(n87701), .A4(n87702), .ZN(
        n87685) );
  NAND2_X1 U73274 ( .A1(n87703), .A2(n87704), .ZN(n87702) );
  AOI22_X1 U73275 ( .A1(n86477), .A2(n110573), .B1(n86478), .B2(n110578), .ZN(
        n87704) );
  AOI22_X1 U73276 ( .A1(n105697), .A2(n110572), .B1(n86480), .B2(n73894), .ZN(
        n87703) );
  NAND2_X1 U73277 ( .A1(n87705), .A2(n87706), .ZN(n87701) );
  AOI22_X1 U73278 ( .A1(n86483), .A2(n73903), .B1(n105694), .B2(n110580), .ZN(
        n87706) );
  AOI22_X1 U73279 ( .A1(n86485), .A2(n110581), .B1(n86486), .B2(n110571), .ZN(
        n87705) );
  NAND2_X1 U73280 ( .A1(n87707), .A2(n87708), .ZN(n87700) );
  AOI22_X1 U73281 ( .A1(n86489), .A2(n110579), .B1(n86490), .B2(n110583), .ZN(
        n87708) );
  AOI22_X1 U73282 ( .A1(n86491), .A2(n110577), .B1(n86492), .B2(n110582), .ZN(
        n87707) );
  NAND2_X1 U73283 ( .A1(n87709), .A2(n87710), .ZN(n87699) );
  AOI22_X1 U73284 ( .A1(n105687), .A2(n73908), .B1(n86496), .B2(n110587), .ZN(
        n87710) );
  AOI22_X1 U73285 ( .A1(n86497), .A2(n73906), .B1(n86498), .B2(n110576), .ZN(
        n87709) );
  NAND2_X1 U73286 ( .A1(n87711), .A2(n87712), .ZN(n87629) );
  NOR4_X1 U73287 ( .A1(n87713), .A2(n87714), .A3(n87715), .A4(n87716), .ZN(
        n87712) );
  NAND2_X1 U73288 ( .A1(n87717), .A2(n87718), .ZN(n87716) );
  AOI22_X1 U73289 ( .A1(n86507), .A2(n110615), .B1(n86508), .B2(n110614), .ZN(
        n87718) );
  AOI22_X1 U73290 ( .A1(n86509), .A2(n73942), .B1(n86510), .B2(n110612), .ZN(
        n87717) );
  NAND2_X1 U73291 ( .A1(n87719), .A2(n87720), .ZN(n87715) );
  AOI22_X1 U73292 ( .A1(n86513), .A2(n110610), .B1(n105678), .B2(n110613), 
        .ZN(n87720) );
  AOI22_X1 U73293 ( .A1(n86515), .A2(n110618), .B1(n86516), .B2(n110611), .ZN(
        n87719) );
  NAND2_X1 U73294 ( .A1(n87721), .A2(n87722), .ZN(n87714) );
  AOI22_X1 U73295 ( .A1(n86519), .A2(n110622), .B1(n86520), .B2(n73954), .ZN(
        n87722) );
  AOI22_X1 U73296 ( .A1(n86521), .A2(n110620), .B1(n86522), .B2(n110621), .ZN(
        n87721) );
  NAND2_X1 U73297 ( .A1(n87723), .A2(n87724), .ZN(n87713) );
  AOI22_X1 U73298 ( .A1(n86525), .A2(n110616), .B1(n86526), .B2(n110619), .ZN(
        n87724) );
  AOI22_X1 U73299 ( .A1(n86527), .A2(n73953), .B1(n86528), .B2(n110617), .ZN(
        n87723) );
  NOR4_X1 U73300 ( .A1(n87725), .A2(n87726), .A3(n87727), .A4(n87728), .ZN(
        n87711) );
  NAND2_X1 U73301 ( .A1(n87729), .A2(n87730), .ZN(n87728) );
  AOI22_X1 U73302 ( .A1(n105675), .A2(n110596), .B1(n86536), .B2(n110600), 
        .ZN(n87730) );
  AOI22_X1 U73303 ( .A1(n86537), .A2(n110599), .B1(n86538), .B2(n73925), .ZN(
        n87729) );
  NAND2_X1 U73304 ( .A1(n87731), .A2(n87732), .ZN(n87727) );
  AOI22_X1 U73305 ( .A1(n86541), .A2(n110606), .B1(n86542), .B2(n110595), .ZN(
        n87732) );
  AOI22_X1 U73306 ( .A1(n86543), .A2(n110598), .B1(n105668), .B2(n110603), 
        .ZN(n87731) );
  NAND2_X1 U73307 ( .A1(n87733), .A2(n87734), .ZN(n87726) );
  AOI22_X1 U73308 ( .A1(n86547), .A2(n110602), .B1(n86548), .B2(n110607), .ZN(
        n87734) );
  AOI22_X1 U73309 ( .A1(n86549), .A2(n110609), .B1(n105664), .B2(n110605), 
        .ZN(n87733) );
  NAND2_X1 U73310 ( .A1(n87735), .A2(n87736), .ZN(n87725) );
  AOI22_X1 U73311 ( .A1(n86553), .A2(n73943), .B1(n86554), .B2(n110601), .ZN(
        n87736) );
  AOI22_X1 U73312 ( .A1(n105661), .A2(n110604), .B1(n105660), .B2(n110608), 
        .ZN(n87735) );
  AOI21_X1 U73313 ( .B1(n86302), .B2(n87738), .A(n87739), .ZN(n87737) );
  OAI21_X1 U73314 ( .B1(n87740), .B2(n105787), .A(n87741), .ZN(n87739) );
  OAI21_X1 U73315 ( .B1(n87742), .B2(n87743), .A(n86310), .ZN(n87741) );
  OAI21_X1 U73316 ( .B1(n110436), .B2(n86311), .A(n87744), .ZN(n87743) );
  AOI22_X1 U73317 ( .A1(n86313), .A2(n73694), .B1(n105784), .B2(n110434), .ZN(
        n87744) );
  NAND2_X1 U73318 ( .A1(n87745), .A2(n87746), .ZN(n87742) );
  AOI22_X1 U73319 ( .A1(n105783), .A2(n110432), .B1(n86318), .B2(n110437), 
        .ZN(n87746) );
  AOI22_X1 U73320 ( .A1(n105781), .A2(n110435), .B1(n86320), .B2(n110433), 
        .ZN(n87745) );
  NOR4_X1 U73321 ( .A1(n87747), .A2(n87748), .A3(n87749), .A4(n87750), .ZN(
        n87740) );
  NAND2_X1 U73322 ( .A1(n87751), .A2(n87752), .ZN(n87750) );
  NOR4_X1 U73323 ( .A1(n87753), .A2(n87754), .A3(n87755), .A4(n87756), .ZN(
        n87752) );
  NAND2_X1 U73324 ( .A1(n87757), .A2(n87758), .ZN(n87756) );
  AOI22_X1 U73325 ( .A1(n105779), .A2(n110413), .B1(n86334), .B2(n110414), 
        .ZN(n87758) );
  AOI22_X1 U73326 ( .A1(n105777), .A2(n110422), .B1(n86336), .B2(n110420), 
        .ZN(n87757) );
  NAND2_X1 U73327 ( .A1(n87759), .A2(n87760), .ZN(n87755) );
  AOI22_X1 U73328 ( .A1(n105775), .A2(n73563), .B1(n86340), .B2(n110417), .ZN(
        n87760) );
  AOI22_X1 U73329 ( .A1(n105773), .A2(n73667), .B1(n86342), .B2(n110339), .ZN(
        n87759) );
  NAND2_X1 U73330 ( .A1(n87761), .A2(n87762), .ZN(n87754) );
  AOI22_X1 U73331 ( .A1(n105771), .A2(n110342), .B1(n86346), .B2(n73567), .ZN(
        n87762) );
  AOI22_X1 U73332 ( .A1(n105769), .A2(n110418), .B1(n86348), .B2(n110415), 
        .ZN(n87761) );
  NAND2_X1 U73333 ( .A1(n87763), .A2(n87764), .ZN(n87753) );
  AOI22_X1 U73334 ( .A1(n105767), .A2(n110340), .B1(n86352), .B2(n110344), 
        .ZN(n87764) );
  AOI22_X1 U73335 ( .A1(n105765), .A2(n110343), .B1(n86354), .B2(n73569), .ZN(
        n87763) );
  NOR4_X1 U73336 ( .A1(n87765), .A2(n87766), .A3(n87767), .A4(n87768), .ZN(
        n87751) );
  NAND2_X1 U73337 ( .A1(n87769), .A2(n87770), .ZN(n87768) );
  AOI22_X1 U73338 ( .A1(n105763), .A2(n110423), .B1(n86362), .B2(n110426), 
        .ZN(n87770) );
  AOI22_X1 U73339 ( .A1(n86363), .A2(n110427), .B1(n105760), .B2(n110429), 
        .ZN(n87769) );
  NAND2_X1 U73340 ( .A1(n87771), .A2(n87772), .ZN(n87767) );
  AOI22_X1 U73341 ( .A1(n105759), .A2(n110428), .B1(n86368), .B2(n110424), 
        .ZN(n87772) );
  AOI22_X1 U73342 ( .A1(n105757), .A2(n110430), .B1(n86370), .B2(n110425), 
        .ZN(n87771) );
  NAND2_X1 U73343 ( .A1(n87773), .A2(n87774), .ZN(n87766) );
  AOI22_X1 U73344 ( .A1(n105755), .A2(n73677), .B1(n86374), .B2(n73676), .ZN(
        n87774) );
  AOI22_X1 U73345 ( .A1(n105753), .A2(n73679), .B1(n86376), .B2(n110431), .ZN(
        n87773) );
  NAND2_X1 U73346 ( .A1(n87775), .A2(n87776), .ZN(n87765) );
  AOI22_X1 U73347 ( .A1(n105751), .A2(n110416), .B1(n86380), .B2(n110421), 
        .ZN(n87776) );
  AOI22_X1 U73348 ( .A1(n105749), .A2(n73674), .B1(n105748), .B2(n110419), 
        .ZN(n87775) );
  NAND2_X1 U73349 ( .A1(n87777), .A2(n87778), .ZN(n87749) );
  NOR4_X1 U73350 ( .A1(n87779), .A2(n87780), .A3(n87781), .A4(n87782), .ZN(
        n87778) );
  NAND2_X1 U73351 ( .A1(n87783), .A2(n87784), .ZN(n87782) );
  AOI22_X1 U73352 ( .A1(n105747), .A2(n110353), .B1(n86392), .B2(n110355), 
        .ZN(n87784) );
  AOI22_X1 U73353 ( .A1(n105745), .A2(n73592), .B1(n86394), .B2(n110354), .ZN(
        n87783) );
  NAND2_X1 U73354 ( .A1(n87785), .A2(n87786), .ZN(n87781) );
  AOI22_X1 U73355 ( .A1(n105743), .A2(n73596), .B1(n86398), .B2(n73598), .ZN(
        n87786) );
  AOI22_X1 U73356 ( .A1(n105741), .A2(n110360), .B1(n86400), .B2(n110361), 
        .ZN(n87785) );
  NAND2_X1 U73357 ( .A1(n87787), .A2(n87788), .ZN(n87780) );
  AOI22_X1 U73358 ( .A1(n86403), .A2(n110358), .B1(n86404), .B2(n110359), .ZN(
        n87788) );
  AOI22_X1 U73359 ( .A1(n105737), .A2(n73597), .B1(n105736), .B2(n73591), .ZN(
        n87787) );
  NAND2_X1 U73360 ( .A1(n87789), .A2(n87790), .ZN(n87779) );
  AOI22_X1 U73361 ( .A1(n105735), .A2(n110366), .B1(n86410), .B2(n73603), .ZN(
        n87790) );
  AOI22_X1 U73362 ( .A1(n86411), .A2(n110365), .B1(n86412), .B2(n73601), .ZN(
        n87789) );
  NOR4_X1 U73363 ( .A1(n87791), .A2(n87792), .A3(n87793), .A4(n87794), .ZN(
        n87777) );
  NAND2_X1 U73364 ( .A1(n87795), .A2(n87796), .ZN(n87794) );
  AOI22_X1 U73365 ( .A1(n105731), .A2(n110348), .B1(n86420), .B2(n111019), 
        .ZN(n87796) );
  AOI22_X1 U73366 ( .A1(n105729), .A2(n110341), .B1(n86422), .B2(n73575), .ZN(
        n87795) );
  NAND2_X1 U73367 ( .A1(n87797), .A2(n87798), .ZN(n87793) );
  AOI22_X1 U73368 ( .A1(n105727), .A2(n110346), .B1(n86426), .B2(n110350), 
        .ZN(n87798) );
  AOI22_X1 U73369 ( .A1(n105725), .A2(n110352), .B1(n86428), .B2(n110349), 
        .ZN(n87797) );
  NAND2_X1 U73370 ( .A1(n87799), .A2(n87800), .ZN(n87792) );
  AOI22_X1 U73371 ( .A1(n105723), .A2(n73584), .B1(n86432), .B2(n110345), .ZN(
        n87800) );
  AOI22_X1 U73372 ( .A1(n105721), .A2(n110347), .B1(n86434), .B2(n110351), 
        .ZN(n87799) );
  NAND2_X1 U73373 ( .A1(n87801), .A2(n87802), .ZN(n87791) );
  AOI22_X1 U73374 ( .A1(n105719), .A2(n110357), .B1(n86438), .B2(n73588), .ZN(
        n87802) );
  AOI22_X1 U73375 ( .A1(n105717), .A2(n73586), .B1(n105716), .B2(n110356), 
        .ZN(n87801) );
  NAND2_X1 U73376 ( .A1(n87803), .A2(n87804), .ZN(n87748) );
  NOR4_X1 U73377 ( .A1(n87805), .A2(n87806), .A3(n87807), .A4(n87808), .ZN(
        n87804) );
  NAND2_X1 U73378 ( .A1(n87809), .A2(n87810), .ZN(n87808) );
  AOI22_X1 U73379 ( .A1(n105715), .A2(n73626), .B1(n86450), .B2(n110376), .ZN(
        n87810) );
  AOI22_X1 U73380 ( .A1(n105713), .A2(n110380), .B1(n86452), .B2(n110379), 
        .ZN(n87809) );
  NAND2_X1 U73381 ( .A1(n87811), .A2(n87812), .ZN(n87807) );
  AOI22_X1 U73382 ( .A1(n105711), .A2(n110383), .B1(n86456), .B2(n110382), 
        .ZN(n87812) );
  AOI22_X1 U73383 ( .A1(n105709), .A2(n110375), .B1(n86458), .B2(n110377), 
        .ZN(n87811) );
  NAND2_X1 U73384 ( .A1(n87813), .A2(n87814), .ZN(n87806) );
  AOI22_X1 U73385 ( .A1(n105707), .A2(n110384), .B1(n86462), .B2(n73625), .ZN(
        n87814) );
  AOI22_X1 U73386 ( .A1(n105705), .A2(n73630), .B1(n86464), .B2(n73632), .ZN(
        n87813) );
  NAND2_X1 U73387 ( .A1(n87815), .A2(n87816), .ZN(n87805) );
  AOI22_X1 U73388 ( .A1(n86467), .A2(n110387), .B1(n86468), .B2(n73638), .ZN(
        n87816) );
  AOI22_X1 U73389 ( .A1(n105701), .A2(n110381), .B1(n86470), .B2(n73627), .ZN(
        n87815) );
  NOR4_X1 U73390 ( .A1(n87817), .A2(n87818), .A3(n87819), .A4(n87820), .ZN(
        n87803) );
  NAND2_X1 U73391 ( .A1(n87821), .A2(n87822), .ZN(n87820) );
  AOI22_X1 U73392 ( .A1(n105699), .A2(n110364), .B1(n86478), .B2(n110369), 
        .ZN(n87822) );
  AOI22_X1 U73393 ( .A1(n105697), .A2(n110363), .B1(n86480), .B2(n73606), .ZN(
        n87821) );
  NAND2_X1 U73394 ( .A1(n87823), .A2(n87824), .ZN(n87819) );
  AOI22_X1 U73395 ( .A1(n105695), .A2(n73615), .B1(n105694), .B2(n110371), 
        .ZN(n87824) );
  AOI22_X1 U73396 ( .A1(n105693), .A2(n110372), .B1(n86486), .B2(n110362), 
        .ZN(n87823) );
  NAND2_X1 U73397 ( .A1(n87825), .A2(n87826), .ZN(n87818) );
  AOI22_X1 U73398 ( .A1(n105691), .A2(n110370), .B1(n86490), .B2(n110374), 
        .ZN(n87826) );
  AOI22_X1 U73399 ( .A1(n105689), .A2(n110368), .B1(n86492), .B2(n110373), 
        .ZN(n87825) );
  NAND2_X1 U73400 ( .A1(n87827), .A2(n87828), .ZN(n87817) );
  AOI22_X1 U73401 ( .A1(n105687), .A2(n73620), .B1(n86496), .B2(n110378), .ZN(
        n87828) );
  AOI22_X1 U73402 ( .A1(n105685), .A2(n73618), .B1(n86498), .B2(n110367), .ZN(
        n87827) );
  NAND2_X1 U73403 ( .A1(n87829), .A2(n87830), .ZN(n87747) );
  NOR4_X1 U73404 ( .A1(n87831), .A2(n87832), .A3(n87833), .A4(n87834), .ZN(
        n87830) );
  NAND2_X1 U73405 ( .A1(n87835), .A2(n87836), .ZN(n87834) );
  AOI22_X1 U73406 ( .A1(n105683), .A2(n110404), .B1(n86508), .B2(n110403), 
        .ZN(n87836) );
  AOI22_X1 U73407 ( .A1(n105681), .A2(n73654), .B1(n86510), .B2(n110401), .ZN(
        n87835) );
  NAND2_X1 U73408 ( .A1(n87837), .A2(n87838), .ZN(n87833) );
  AOI22_X1 U73409 ( .A1(n105679), .A2(n110399), .B1(n105678), .B2(n110402), 
        .ZN(n87838) );
  AOI22_X1 U73410 ( .A1(n86515), .A2(n73660), .B1(n86516), .B2(n110400), .ZN(
        n87837) );
  NAND2_X1 U73411 ( .A1(n87839), .A2(n87840), .ZN(n87832) );
  AOI22_X1 U73412 ( .A1(n86519), .A2(n110410), .B1(n86520), .B2(n73666), .ZN(
        n87840) );
  AOI22_X1 U73413 ( .A1(n86521), .A2(n110408), .B1(n86522), .B2(n110409), .ZN(
        n87839) );
  NAND2_X1 U73414 ( .A1(n87841), .A2(n87842), .ZN(n87831) );
  AOI22_X1 U73415 ( .A1(n105676), .A2(n110405), .B1(n86526), .B2(n110407), 
        .ZN(n87842) );
  AOI22_X1 U73416 ( .A1(n86527), .A2(n110411), .B1(n86528), .B2(n110406), .ZN(
        n87841) );
  NOR4_X1 U73417 ( .A1(n87843), .A2(n87844), .A3(n87845), .A4(n87846), .ZN(
        n87829) );
  NAND2_X1 U73418 ( .A1(n87847), .A2(n87848), .ZN(n87846) );
  AOI22_X1 U73419 ( .A1(n105675), .A2(n110386), .B1(n86536), .B2(n110389), 
        .ZN(n87848) );
  AOI22_X1 U73420 ( .A1(n105673), .A2(n111038), .B1(n86538), .B2(n73637), .ZN(
        n87847) );
  NAND2_X1 U73421 ( .A1(n87849), .A2(n87850), .ZN(n87845) );
  AOI22_X1 U73422 ( .A1(n105671), .A2(n110395), .B1(n86542), .B2(n110385), 
        .ZN(n87850) );
  AOI22_X1 U73423 ( .A1(n105669), .A2(n110388), .B1(n105668), .B2(n110392), 
        .ZN(n87849) );
  NAND2_X1 U73424 ( .A1(n87851), .A2(n87852), .ZN(n87844) );
  AOI22_X1 U73425 ( .A1(n105667), .A2(n110391), .B1(n86548), .B2(n110396), 
        .ZN(n87852) );
  AOI22_X1 U73426 ( .A1(n86549), .A2(n110398), .B1(n105664), .B2(n110394), 
        .ZN(n87851) );
  NAND2_X1 U73427 ( .A1(n87853), .A2(n87854), .ZN(n87843) );
  AOI22_X1 U73428 ( .A1(n105663), .A2(n73655), .B1(n86554), .B2(n110390), .ZN(
        n87854) );
  AOI22_X1 U73429 ( .A1(n105661), .A2(n110393), .B1(n105660), .B2(n110397), 
        .ZN(n87853) );
  AOI21_X1 U73430 ( .B1(n86302), .B2(n87856), .A(n87857), .ZN(n87855) );
  OAI21_X1 U73431 ( .B1(n87858), .B2(n105787), .A(n87859), .ZN(n87857) );
  OAI21_X1 U73432 ( .B1(n87860), .B2(n87861), .A(n105786), .ZN(n87859) );
  OAI21_X1 U73433 ( .B1(n110114), .B2(n105785), .A(n87862), .ZN(n87861) );
  AOI22_X1 U73434 ( .A1(n86313), .A2(n73256), .B1(n105784), .B2(n110112), .ZN(
        n87862) );
  NAND2_X1 U73435 ( .A1(n87863), .A2(n87864), .ZN(n87860) );
  AOI22_X1 U73436 ( .A1(n105783), .A2(n110110), .B1(n105782), .B2(n110115), 
        .ZN(n87864) );
  AOI22_X1 U73437 ( .A1(n105781), .A2(n110113), .B1(n105780), .B2(n110111), 
        .ZN(n87863) );
  NOR4_X1 U73438 ( .A1(n87865), .A2(n87866), .A3(n87867), .A4(n87868), .ZN(
        n87858) );
  NAND2_X1 U73439 ( .A1(n87869), .A2(n87870), .ZN(n87868) );
  NOR4_X1 U73440 ( .A1(n87871), .A2(n87872), .A3(n87873), .A4(n87874), .ZN(
        n87870) );
  NAND2_X1 U73441 ( .A1(n87875), .A2(n87876), .ZN(n87874) );
  AOI22_X1 U73442 ( .A1(n105779), .A2(n110091), .B1(n105778), .B2(n110092), 
        .ZN(n87876) );
  AOI22_X1 U73443 ( .A1(n105777), .A2(n110100), .B1(n105776), .B2(n110098), 
        .ZN(n87875) );
  NAND2_X1 U73444 ( .A1(n87877), .A2(n87878), .ZN(n87873) );
  AOI22_X1 U73445 ( .A1(n105775), .A2(n73125), .B1(n105774), .B2(n110095), 
        .ZN(n87878) );
  AOI22_X1 U73446 ( .A1(n105773), .A2(n73229), .B1(n105772), .B2(n110013), 
        .ZN(n87877) );
  NAND2_X1 U73447 ( .A1(n87879), .A2(n87880), .ZN(n87872) );
  AOI22_X1 U73448 ( .A1(n105771), .A2(n110017), .B1(n86346), .B2(n73129), .ZN(
        n87880) );
  AOI22_X1 U73449 ( .A1(n105769), .A2(n110096), .B1(n105768), .B2(n110093), 
        .ZN(n87879) );
  NAND2_X1 U73450 ( .A1(n87881), .A2(n87882), .ZN(n87871) );
  AOI22_X1 U73451 ( .A1(n105767), .A2(n110015), .B1(n105766), .B2(n110019), 
        .ZN(n87882) );
  AOI22_X1 U73452 ( .A1(n105765), .A2(n110018), .B1(n105764), .B2(n73131), 
        .ZN(n87881) );
  NOR4_X1 U73453 ( .A1(n87883), .A2(n87884), .A3(n87885), .A4(n87886), .ZN(
        n87869) );
  NAND2_X1 U73454 ( .A1(n87887), .A2(n87888), .ZN(n87886) );
  AOI22_X1 U73455 ( .A1(n105763), .A2(n110101), .B1(n105762), .B2(n110104), 
        .ZN(n87888) );
  AOI22_X1 U73456 ( .A1(n86363), .A2(n110105), .B1(n105760), .B2(n110107), 
        .ZN(n87887) );
  NAND2_X1 U73457 ( .A1(n87889), .A2(n87890), .ZN(n87885) );
  AOI22_X1 U73458 ( .A1(n105759), .A2(n110106), .B1(n86368), .B2(n110102), 
        .ZN(n87890) );
  AOI22_X1 U73459 ( .A1(n105757), .A2(n110108), .B1(n105756), .B2(n110103), 
        .ZN(n87889) );
  NAND2_X1 U73460 ( .A1(n87891), .A2(n87892), .ZN(n87884) );
  AOI22_X1 U73461 ( .A1(n105755), .A2(n73239), .B1(n105754), .B2(n73238), .ZN(
        n87892) );
  AOI22_X1 U73462 ( .A1(n105753), .A2(n73241), .B1(n105752), .B2(n110109), 
        .ZN(n87891) );
  NAND2_X1 U73463 ( .A1(n87893), .A2(n87894), .ZN(n87883) );
  AOI22_X1 U73464 ( .A1(n105751), .A2(n110094), .B1(n105750), .B2(n110099), 
        .ZN(n87894) );
  AOI22_X1 U73465 ( .A1(n105749), .A2(n73236), .B1(n105748), .B2(n110097), 
        .ZN(n87893) );
  NAND2_X1 U73466 ( .A1(n87895), .A2(n87896), .ZN(n87867) );
  NOR4_X1 U73467 ( .A1(n87897), .A2(n87898), .A3(n87899), .A4(n87900), .ZN(
        n87896) );
  NAND2_X1 U73468 ( .A1(n87901), .A2(n87902), .ZN(n87900) );
  AOI22_X1 U73469 ( .A1(n105747), .A2(n110028), .B1(n105746), .B2(n110030), 
        .ZN(n87902) );
  AOI22_X1 U73470 ( .A1(n105745), .A2(n73154), .B1(n105744), .B2(n110029), 
        .ZN(n87901) );
  NAND2_X1 U73471 ( .A1(n87903), .A2(n87904), .ZN(n87899) );
  AOI22_X1 U73472 ( .A1(n105743), .A2(n73158), .B1(n105742), .B2(n73160), .ZN(
        n87904) );
  AOI22_X1 U73473 ( .A1(n105741), .A2(n110036), .B1(n86400), .B2(n110037), 
        .ZN(n87903) );
  NAND2_X1 U73474 ( .A1(n87905), .A2(n87906), .ZN(n87898) );
  AOI22_X1 U73475 ( .A1(n86403), .A2(n110033), .B1(n105738), .B2(n110035), 
        .ZN(n87906) );
  AOI22_X1 U73476 ( .A1(n105737), .A2(n73159), .B1(n105736), .B2(n110034), 
        .ZN(n87905) );
  NAND2_X1 U73477 ( .A1(n87907), .A2(n87908), .ZN(n87897) );
  AOI22_X1 U73478 ( .A1(n105735), .A2(n110042), .B1(n105734), .B2(n73165), 
        .ZN(n87908) );
  AOI22_X1 U73479 ( .A1(n86411), .A2(n110041), .B1(n105732), .B2(n73163), .ZN(
        n87907) );
  NOR4_X1 U73480 ( .A1(n87909), .A2(n87910), .A3(n87911), .A4(n87912), .ZN(
        n87895) );
  NAND2_X1 U73481 ( .A1(n87913), .A2(n87914), .ZN(n87912) );
  AOI22_X1 U73482 ( .A1(n105731), .A2(n110023), .B1(n105730), .B2(n110014), 
        .ZN(n87914) );
  AOI22_X1 U73483 ( .A1(n105729), .A2(n110016), .B1(n105728), .B2(n73137), 
        .ZN(n87913) );
  NAND2_X1 U73484 ( .A1(n87915), .A2(n87916), .ZN(n87911) );
  AOI22_X1 U73485 ( .A1(n105727), .A2(n110021), .B1(n86426), .B2(n110025), 
        .ZN(n87916) );
  AOI22_X1 U73486 ( .A1(n105725), .A2(n110027), .B1(n86428), .B2(n110024), 
        .ZN(n87915) );
  NAND2_X1 U73487 ( .A1(n87917), .A2(n87918), .ZN(n87910) );
  AOI22_X1 U73488 ( .A1(n105723), .A2(n73146), .B1(n105722), .B2(n110020), 
        .ZN(n87918) );
  AOI22_X1 U73489 ( .A1(n105721), .A2(n110022), .B1(n105720), .B2(n110026), 
        .ZN(n87917) );
  NAND2_X1 U73490 ( .A1(n87919), .A2(n87920), .ZN(n87909) );
  AOI22_X1 U73491 ( .A1(n105719), .A2(n110032), .B1(n105718), .B2(n73150), 
        .ZN(n87920) );
  AOI22_X1 U73492 ( .A1(n105717), .A2(n73148), .B1(n105716), .B2(n110031), 
        .ZN(n87919) );
  NAND2_X1 U73493 ( .A1(n87921), .A2(n87922), .ZN(n87866) );
  NOR4_X1 U73494 ( .A1(n87923), .A2(n87924), .A3(n87925), .A4(n87926), .ZN(
        n87922) );
  NAND2_X1 U73495 ( .A1(n87927), .A2(n87928), .ZN(n87926) );
  AOI22_X1 U73496 ( .A1(n105715), .A2(n73188), .B1(n86450), .B2(n110052), .ZN(
        n87928) );
  AOI22_X1 U73497 ( .A1(n105713), .A2(n110056), .B1(n105712), .B2(n110055), 
        .ZN(n87927) );
  NAND2_X1 U73498 ( .A1(n87929), .A2(n87930), .ZN(n87925) );
  AOI22_X1 U73499 ( .A1(n105711), .A2(n110061), .B1(n105710), .B2(n110060), 
        .ZN(n87930) );
  AOI22_X1 U73500 ( .A1(n105709), .A2(n110051), .B1(n105708), .B2(n110053), 
        .ZN(n87929) );
  NAND2_X1 U73501 ( .A1(n87931), .A2(n87932), .ZN(n87924) );
  AOI22_X1 U73502 ( .A1(n105707), .A2(n110062), .B1(n105706), .B2(n110058), 
        .ZN(n87932) );
  AOI22_X1 U73503 ( .A1(n105705), .A2(n73192), .B1(n105704), .B2(n73194), .ZN(
        n87931) );
  NAND2_X1 U73504 ( .A1(n87933), .A2(n87934), .ZN(n87923) );
  AOI22_X1 U73505 ( .A1(n86467), .A2(n110065), .B1(n105702), .B2(n73200), .ZN(
        n87934) );
  AOI22_X1 U73506 ( .A1(n105701), .A2(n110057), .B1(n105700), .B2(n110059), 
        .ZN(n87933) );
  NOR4_X1 U73507 ( .A1(n87935), .A2(n87936), .A3(n87937), .A4(n87938), .ZN(
        n87921) );
  NAND2_X1 U73508 ( .A1(n87939), .A2(n87940), .ZN(n87938) );
  AOI22_X1 U73509 ( .A1(n105699), .A2(n110040), .B1(n105698), .B2(n110045), 
        .ZN(n87940) );
  AOI22_X1 U73510 ( .A1(n105697), .A2(n110039), .B1(n105696), .B2(n73168), 
        .ZN(n87939) );
  NAND2_X1 U73511 ( .A1(n87941), .A2(n87942), .ZN(n87937) );
  AOI22_X1 U73512 ( .A1(n105695), .A2(n73177), .B1(n105694), .B2(n110047), 
        .ZN(n87942) );
  AOI22_X1 U73513 ( .A1(n105693), .A2(n110048), .B1(n105692), .B2(n110038), 
        .ZN(n87941) );
  NAND2_X1 U73514 ( .A1(n87943), .A2(n87944), .ZN(n87936) );
  AOI22_X1 U73515 ( .A1(n105691), .A2(n110046), .B1(n86490), .B2(n110050), 
        .ZN(n87944) );
  AOI22_X1 U73516 ( .A1(n105689), .A2(n110044), .B1(n105688), .B2(n110049), 
        .ZN(n87943) );
  NAND2_X1 U73517 ( .A1(n87945), .A2(n87946), .ZN(n87935) );
  AOI22_X1 U73518 ( .A1(n105687), .A2(n73182), .B1(n105686), .B2(n110054), 
        .ZN(n87946) );
  AOI22_X1 U73519 ( .A1(n105685), .A2(n73180), .B1(n105684), .B2(n110043), 
        .ZN(n87945) );
  NAND2_X1 U73520 ( .A1(n87947), .A2(n87948), .ZN(n87865) );
  NOR4_X1 U73521 ( .A1(n87949), .A2(n87950), .A3(n87951), .A4(n87952), .ZN(
        n87948) );
  NAND2_X1 U73522 ( .A1(n87953), .A2(n87954), .ZN(n87952) );
  AOI22_X1 U73523 ( .A1(n105683), .A2(n110082), .B1(n105682), .B2(n110081), 
        .ZN(n87954) );
  AOI22_X1 U73524 ( .A1(n105681), .A2(n73216), .B1(n105680), .B2(n110079), 
        .ZN(n87953) );
  NAND2_X1 U73525 ( .A1(n87955), .A2(n87956), .ZN(n87951) );
  AOI22_X1 U73526 ( .A1(n105679), .A2(n110077), .B1(n105678), .B2(n110080), 
        .ZN(n87956) );
  AOI22_X1 U73527 ( .A1(n86515), .A2(n73222), .B1(n86516), .B2(n110078), .ZN(
        n87955) );
  NAND2_X1 U73528 ( .A1(n87957), .A2(n87958), .ZN(n87950) );
  AOI22_X1 U73529 ( .A1(n86519), .A2(n110088), .B1(n86520), .B2(n73228), .ZN(
        n87958) );
  AOI22_X1 U73530 ( .A1(n86521), .A2(n110086), .B1(n86522), .B2(n110087), .ZN(
        n87957) );
  NAND2_X1 U73531 ( .A1(n87959), .A2(n87960), .ZN(n87949) );
  AOI22_X1 U73532 ( .A1(n105676), .A2(n110083), .B1(n86526), .B2(n110085), 
        .ZN(n87960) );
  AOI22_X1 U73533 ( .A1(n86527), .A2(n110089), .B1(n86528), .B2(n110084), .ZN(
        n87959) );
  NOR4_X1 U73534 ( .A1(n87961), .A2(n87962), .A3(n87963), .A4(n87964), .ZN(
        n87947) );
  NAND2_X1 U73535 ( .A1(n87965), .A2(n87966), .ZN(n87964) );
  AOI22_X1 U73536 ( .A1(n105675), .A2(n110064), .B1(n105674), .B2(n110067), 
        .ZN(n87966) );
  AOI22_X1 U73537 ( .A1(n105673), .A2(n111040), .B1(n105672), .B2(n73199), 
        .ZN(n87965) );
  NAND2_X1 U73538 ( .A1(n87967), .A2(n87968), .ZN(n87963) );
  AOI22_X1 U73539 ( .A1(n105671), .A2(n110073), .B1(n105670), .B2(n110063), 
        .ZN(n87968) );
  AOI22_X1 U73540 ( .A1(n105669), .A2(n110066), .B1(n105668), .B2(n110070), 
        .ZN(n87967) );
  NAND2_X1 U73541 ( .A1(n87969), .A2(n87970), .ZN(n87962) );
  AOI22_X1 U73542 ( .A1(n105667), .A2(n110069), .B1(n105666), .B2(n110074), 
        .ZN(n87970) );
  AOI22_X1 U73543 ( .A1(n86549), .A2(n110076), .B1(n105664), .B2(n110072), 
        .ZN(n87969) );
  NAND2_X1 U73544 ( .A1(n87971), .A2(n87972), .ZN(n87961) );
  AOI22_X1 U73545 ( .A1(n105663), .A2(n73217), .B1(n105662), .B2(n110068), 
        .ZN(n87972) );
  AOI22_X1 U73546 ( .A1(n105661), .A2(n110071), .B1(n105660), .B2(n110075), 
        .ZN(n87971) );
  AOI21_X1 U73547 ( .B1(n86302), .B2(n87974), .A(n87975), .ZN(n87973) );
  OAI21_X1 U73548 ( .B1(n87976), .B2(n105787), .A(n87977), .ZN(n87975) );
  OAI21_X1 U73549 ( .B1(n87978), .B2(n87979), .A(n105786), .ZN(n87977) );
  OAI21_X1 U73550 ( .B1(n110221), .B2(n86311), .A(n87980), .ZN(n87979) );
  AOI22_X1 U73551 ( .A1(n86313), .A2(n73398), .B1(n105784), .B2(n110219), .ZN(
        n87980) );
  NAND2_X1 U73552 ( .A1(n87981), .A2(n87982), .ZN(n87978) );
  AOI22_X1 U73553 ( .A1(n105783), .A2(n110217), .B1(n105782), .B2(n110222), 
        .ZN(n87982) );
  AOI22_X1 U73554 ( .A1(n105781), .A2(n110220), .B1(n105780), .B2(n110218), 
        .ZN(n87981) );
  NOR4_X1 U73555 ( .A1(n87983), .A2(n87984), .A3(n87985), .A4(n87986), .ZN(
        n87976) );
  NAND2_X1 U73556 ( .A1(n87987), .A2(n87988), .ZN(n87986) );
  NOR4_X1 U73557 ( .A1(n87989), .A2(n87990), .A3(n87991), .A4(n87992), .ZN(
        n87988) );
  NAND2_X1 U73558 ( .A1(n87993), .A2(n87994), .ZN(n87992) );
  AOI22_X1 U73559 ( .A1(n105779), .A2(n110198), .B1(n105778), .B2(n110199), 
        .ZN(n87994) );
  AOI22_X1 U73560 ( .A1(n105777), .A2(n110207), .B1(n105776), .B2(n110205), 
        .ZN(n87993) );
  NAND2_X1 U73561 ( .A1(n87995), .A2(n87996), .ZN(n87991) );
  AOI22_X1 U73562 ( .A1(n105775), .A2(n73267), .B1(n105774), .B2(n110202), 
        .ZN(n87996) );
  AOI22_X1 U73563 ( .A1(n105773), .A2(n73371), .B1(n105772), .B2(n110121), 
        .ZN(n87995) );
  NAND2_X1 U73564 ( .A1(n87997), .A2(n87998), .ZN(n87990) );
  AOI22_X1 U73565 ( .A1(n105771), .A2(n110124), .B1(n86346), .B2(n73271), .ZN(
        n87998) );
  AOI22_X1 U73566 ( .A1(n105769), .A2(n110203), .B1(n105768), .B2(n110200), 
        .ZN(n87997) );
  NAND2_X1 U73567 ( .A1(n87999), .A2(n88000), .ZN(n87989) );
  AOI22_X1 U73568 ( .A1(n105767), .A2(n110122), .B1(n105766), .B2(n110126), 
        .ZN(n88000) );
  AOI22_X1 U73569 ( .A1(n105765), .A2(n110125), .B1(n105764), .B2(n73273), 
        .ZN(n87999) );
  NOR4_X1 U73570 ( .A1(n88001), .A2(n88002), .A3(n88003), .A4(n88004), .ZN(
        n87987) );
  NAND2_X1 U73571 ( .A1(n88005), .A2(n88006), .ZN(n88004) );
  AOI22_X1 U73572 ( .A1(n105763), .A2(n110208), .B1(n105762), .B2(n110211), 
        .ZN(n88006) );
  AOI22_X1 U73573 ( .A1(n86363), .A2(n110212), .B1(n105760), .B2(n110214), 
        .ZN(n88005) );
  NAND2_X1 U73574 ( .A1(n88007), .A2(n88008), .ZN(n88003) );
  AOI22_X1 U73575 ( .A1(n105759), .A2(n110213), .B1(n86368), .B2(n110209), 
        .ZN(n88008) );
  AOI22_X1 U73576 ( .A1(n105757), .A2(n110215), .B1(n105756), .B2(n110210), 
        .ZN(n88007) );
  NAND2_X1 U73577 ( .A1(n88009), .A2(n88010), .ZN(n88002) );
  AOI22_X1 U73578 ( .A1(n105755), .A2(n73381), .B1(n105754), .B2(n73380), .ZN(
        n88010) );
  AOI22_X1 U73579 ( .A1(n105753), .A2(n73383), .B1(n105752), .B2(n110216), 
        .ZN(n88009) );
  NAND2_X1 U73580 ( .A1(n88011), .A2(n88012), .ZN(n88001) );
  AOI22_X1 U73581 ( .A1(n105751), .A2(n110201), .B1(n105750), .B2(n110206), 
        .ZN(n88012) );
  AOI22_X1 U73582 ( .A1(n105749), .A2(n73378), .B1(n105748), .B2(n110204), 
        .ZN(n88011) );
  NAND2_X1 U73583 ( .A1(n88013), .A2(n88014), .ZN(n87985) );
  NOR4_X1 U73584 ( .A1(n88015), .A2(n88016), .A3(n88017), .A4(n88018), .ZN(
        n88014) );
  NAND2_X1 U73585 ( .A1(n88019), .A2(n88020), .ZN(n88018) );
  AOI22_X1 U73586 ( .A1(n105747), .A2(n110135), .B1(n105746), .B2(n110137), 
        .ZN(n88020) );
  AOI22_X1 U73587 ( .A1(n105745), .A2(n73296), .B1(n105744), .B2(n110136), 
        .ZN(n88019) );
  NAND2_X1 U73588 ( .A1(n88021), .A2(n88022), .ZN(n88017) );
  AOI22_X1 U73589 ( .A1(n105743), .A2(n73300), .B1(n105742), .B2(n73302), .ZN(
        n88022) );
  AOI22_X1 U73590 ( .A1(n105741), .A2(n110143), .B1(n86400), .B2(n110144), 
        .ZN(n88021) );
  NAND2_X1 U73591 ( .A1(n88023), .A2(n88024), .ZN(n88016) );
  AOI22_X1 U73592 ( .A1(n86403), .A2(n110140), .B1(n105738), .B2(n110142), 
        .ZN(n88024) );
  AOI22_X1 U73593 ( .A1(n105737), .A2(n73301), .B1(n105736), .B2(n110141), 
        .ZN(n88023) );
  NAND2_X1 U73594 ( .A1(n88025), .A2(n88026), .ZN(n88015) );
  AOI22_X1 U73595 ( .A1(n105735), .A2(n110149), .B1(n105734), .B2(n73307), 
        .ZN(n88026) );
  AOI22_X1 U73596 ( .A1(n86411), .A2(n110148), .B1(n105732), .B2(n73305), .ZN(
        n88025) );
  NOR4_X1 U73597 ( .A1(n88027), .A2(n88028), .A3(n88029), .A4(n88030), .ZN(
        n88013) );
  NAND2_X1 U73598 ( .A1(n88031), .A2(n88032), .ZN(n88030) );
  AOI22_X1 U73599 ( .A1(n105731), .A2(n110130), .B1(n105730), .B2(n111021), 
        .ZN(n88032) );
  AOI22_X1 U73600 ( .A1(n105729), .A2(n110123), .B1(n105728), .B2(n73279), 
        .ZN(n88031) );
  NAND2_X1 U73601 ( .A1(n88033), .A2(n88034), .ZN(n88029) );
  AOI22_X1 U73602 ( .A1(n105727), .A2(n110128), .B1(n86426), .B2(n110132), 
        .ZN(n88034) );
  AOI22_X1 U73603 ( .A1(n105725), .A2(n110134), .B1(n86428), .B2(n110131), 
        .ZN(n88033) );
  NAND2_X1 U73604 ( .A1(n88035), .A2(n88036), .ZN(n88028) );
  AOI22_X1 U73605 ( .A1(n105723), .A2(n73288), .B1(n105722), .B2(n110127), 
        .ZN(n88036) );
  AOI22_X1 U73606 ( .A1(n105721), .A2(n110129), .B1(n105720), .B2(n110133), 
        .ZN(n88035) );
  NAND2_X1 U73607 ( .A1(n88037), .A2(n88038), .ZN(n88027) );
  AOI22_X1 U73608 ( .A1(n105719), .A2(n110139), .B1(n105718), .B2(n73292), 
        .ZN(n88038) );
  AOI22_X1 U73609 ( .A1(n105717), .A2(n73290), .B1(n105716), .B2(n110138), 
        .ZN(n88037) );
  NAND2_X1 U73610 ( .A1(n88039), .A2(n88040), .ZN(n87984) );
  NOR4_X1 U73611 ( .A1(n88041), .A2(n88042), .A3(n88043), .A4(n88044), .ZN(
        n88040) );
  NAND2_X1 U73612 ( .A1(n88045), .A2(n88046), .ZN(n88044) );
  AOI22_X1 U73613 ( .A1(n105715), .A2(n73330), .B1(n86450), .B2(n110159), .ZN(
        n88046) );
  AOI22_X1 U73614 ( .A1(n105713), .A2(n110163), .B1(n105712), .B2(n110162), 
        .ZN(n88045) );
  NAND2_X1 U73615 ( .A1(n88047), .A2(n88048), .ZN(n88043) );
  AOI22_X1 U73616 ( .A1(n105711), .A2(n110168), .B1(n105710), .B2(n110167), 
        .ZN(n88048) );
  AOI22_X1 U73617 ( .A1(n105709), .A2(n110158), .B1(n86458), .B2(n110160), 
        .ZN(n88047) );
  NAND2_X1 U73618 ( .A1(n88049), .A2(n88050), .ZN(n88042) );
  AOI22_X1 U73619 ( .A1(n105707), .A2(n110169), .B1(n105706), .B2(n110165), 
        .ZN(n88050) );
  AOI22_X1 U73620 ( .A1(n105705), .A2(n73334), .B1(n105704), .B2(n73336), .ZN(
        n88049) );
  NAND2_X1 U73621 ( .A1(n88051), .A2(n88052), .ZN(n88041) );
  AOI22_X1 U73622 ( .A1(n86467), .A2(n110172), .B1(n105702), .B2(n73342), .ZN(
        n88052) );
  AOI22_X1 U73623 ( .A1(n105701), .A2(n110164), .B1(n105700), .B2(n110166), 
        .ZN(n88051) );
  NOR4_X1 U73624 ( .A1(n88053), .A2(n88054), .A3(n88055), .A4(n88056), .ZN(
        n88039) );
  NAND2_X1 U73625 ( .A1(n88057), .A2(n88058), .ZN(n88056) );
  AOI22_X1 U73626 ( .A1(n105699), .A2(n110147), .B1(n105698), .B2(n110152), 
        .ZN(n88058) );
  AOI22_X1 U73627 ( .A1(n105697), .A2(n110146), .B1(n105696), .B2(n73310), 
        .ZN(n88057) );
  NAND2_X1 U73628 ( .A1(n88059), .A2(n88060), .ZN(n88055) );
  AOI22_X1 U73629 ( .A1(n105695), .A2(n73319), .B1(n105694), .B2(n110154), 
        .ZN(n88060) );
  AOI22_X1 U73630 ( .A1(n105693), .A2(n110155), .B1(n105692), .B2(n110145), 
        .ZN(n88059) );
  NAND2_X1 U73631 ( .A1(n88061), .A2(n88062), .ZN(n88054) );
  AOI22_X1 U73632 ( .A1(n105691), .A2(n110153), .B1(n86490), .B2(n110157), 
        .ZN(n88062) );
  AOI22_X1 U73633 ( .A1(n105689), .A2(n110151), .B1(n105688), .B2(n110156), 
        .ZN(n88061) );
  NAND2_X1 U73634 ( .A1(n88063), .A2(n88064), .ZN(n88053) );
  AOI22_X1 U73635 ( .A1(n105687), .A2(n73324), .B1(n105686), .B2(n110161), 
        .ZN(n88064) );
  AOI22_X1 U73636 ( .A1(n105685), .A2(n73322), .B1(n105684), .B2(n110150), 
        .ZN(n88063) );
  NAND2_X1 U73637 ( .A1(n88065), .A2(n88066), .ZN(n87983) );
  NOR4_X1 U73638 ( .A1(n88067), .A2(n88068), .A3(n88069), .A4(n88070), .ZN(
        n88066) );
  NAND2_X1 U73639 ( .A1(n88071), .A2(n88072), .ZN(n88070) );
  AOI22_X1 U73640 ( .A1(n105683), .A2(n110189), .B1(n105682), .B2(n110188), 
        .ZN(n88072) );
  AOI22_X1 U73641 ( .A1(n105681), .A2(n73358), .B1(n105680), .B2(n110186), 
        .ZN(n88071) );
  NAND2_X1 U73642 ( .A1(n88073), .A2(n88074), .ZN(n88069) );
  AOI22_X1 U73643 ( .A1(n105679), .A2(n110184), .B1(n105678), .B2(n110187), 
        .ZN(n88074) );
  AOI22_X1 U73644 ( .A1(n86515), .A2(n73364), .B1(n86516), .B2(n110185), .ZN(
        n88073) );
  NAND2_X1 U73645 ( .A1(n88075), .A2(n88076), .ZN(n88068) );
  AOI22_X1 U73646 ( .A1(n86519), .A2(n110195), .B1(n86520), .B2(n73370), .ZN(
        n88076) );
  AOI22_X1 U73647 ( .A1(n86521), .A2(n110193), .B1(n86522), .B2(n110194), .ZN(
        n88075) );
  NAND2_X1 U73648 ( .A1(n88077), .A2(n88078), .ZN(n88067) );
  AOI22_X1 U73649 ( .A1(n105676), .A2(n110190), .B1(n86526), .B2(n110192), 
        .ZN(n88078) );
  AOI22_X1 U73650 ( .A1(n86527), .A2(n110196), .B1(n86528), .B2(n110191), .ZN(
        n88077) );
  NOR4_X1 U73651 ( .A1(n88079), .A2(n88080), .A3(n88081), .A4(n88082), .ZN(
        n88065) );
  NAND2_X1 U73652 ( .A1(n88083), .A2(n88084), .ZN(n88082) );
  AOI22_X1 U73653 ( .A1(n105675), .A2(n110171), .B1(n105674), .B2(n110174), 
        .ZN(n88084) );
  AOI22_X1 U73654 ( .A1(n105673), .A2(n111035), .B1(n105672), .B2(n73341), 
        .ZN(n88083) );
  NAND2_X1 U73655 ( .A1(n88085), .A2(n88086), .ZN(n88081) );
  AOI22_X1 U73656 ( .A1(n105671), .A2(n110180), .B1(n105670), .B2(n110170), 
        .ZN(n88086) );
  AOI22_X1 U73657 ( .A1(n105669), .A2(n110173), .B1(n105668), .B2(n110177), 
        .ZN(n88085) );
  NAND2_X1 U73658 ( .A1(n88087), .A2(n88088), .ZN(n88080) );
  AOI22_X1 U73659 ( .A1(n105667), .A2(n110176), .B1(n105666), .B2(n110181), 
        .ZN(n88088) );
  AOI22_X1 U73660 ( .A1(n86549), .A2(n110183), .B1(n105664), .B2(n110179), 
        .ZN(n88087) );
  NAND2_X1 U73661 ( .A1(n88089), .A2(n88090), .ZN(n88079) );
  AOI22_X1 U73662 ( .A1(n105663), .A2(n73359), .B1(n105662), .B2(n110175), 
        .ZN(n88090) );
  AOI22_X1 U73663 ( .A1(n105661), .A2(n110178), .B1(n105660), .B2(n110182), 
        .ZN(n88089) );
  AOI21_X1 U73664 ( .B1(n86302), .B2(n88092), .A(n88093), .ZN(n88091) );
  OAI21_X1 U73665 ( .B1(n88094), .B2(n105787), .A(n88095), .ZN(n88093) );
  OAI21_X1 U73666 ( .B1(n88096), .B2(n88097), .A(n105786), .ZN(n88095) );
  OAI21_X1 U73667 ( .B1(n110006), .B2(n105785), .A(n88098), .ZN(n88097) );
  AOI22_X1 U73668 ( .A1(n86313), .A2(n73114), .B1(n105784), .B2(n110004), .ZN(
        n88098) );
  NAND2_X1 U73669 ( .A1(n88099), .A2(n88100), .ZN(n88096) );
  AOI22_X1 U73670 ( .A1(n105783), .A2(n110002), .B1(n105782), .B2(n110007), 
        .ZN(n88100) );
  AOI22_X1 U73671 ( .A1(n105781), .A2(n110005), .B1(n105780), .B2(n110003), 
        .ZN(n88099) );
  NOR4_X1 U73672 ( .A1(n88101), .A2(n88102), .A3(n88103), .A4(n88104), .ZN(
        n88094) );
  NAND2_X1 U73673 ( .A1(n88105), .A2(n88106), .ZN(n88104) );
  NOR4_X1 U73674 ( .A1(n88107), .A2(n88108), .A3(n88109), .A4(n88110), .ZN(
        n88106) );
  NAND2_X1 U73675 ( .A1(n88111), .A2(n88112), .ZN(n88110) );
  AOI22_X1 U73676 ( .A1(n105779), .A2(n109983), .B1(n105778), .B2(n109984), 
        .ZN(n88112) );
  AOI22_X1 U73677 ( .A1(n105777), .A2(n109992), .B1(n105776), .B2(n109990), 
        .ZN(n88111) );
  NAND2_X1 U73678 ( .A1(n88113), .A2(n88114), .ZN(n88109) );
  AOI22_X1 U73679 ( .A1(n105775), .A2(n72983), .B1(n105774), .B2(n109987), 
        .ZN(n88114) );
  AOI22_X1 U73680 ( .A1(n105773), .A2(n73087), .B1(n105772), .B2(n109904), 
        .ZN(n88113) );
  NAND2_X1 U73681 ( .A1(n88115), .A2(n88116), .ZN(n88108) );
  AOI22_X1 U73682 ( .A1(n105771), .A2(n109908), .B1(n86346), .B2(n72987), .ZN(
        n88116) );
  AOI22_X1 U73683 ( .A1(n105769), .A2(n109988), .B1(n105768), .B2(n109985), 
        .ZN(n88115) );
  NAND2_X1 U73684 ( .A1(n88117), .A2(n88118), .ZN(n88107) );
  AOI22_X1 U73685 ( .A1(n105767), .A2(n109906), .B1(n105766), .B2(n109910), 
        .ZN(n88118) );
  AOI22_X1 U73686 ( .A1(n105765), .A2(n109909), .B1(n105764), .B2(n72989), 
        .ZN(n88117) );
  NOR4_X1 U73687 ( .A1(n88119), .A2(n88120), .A3(n88121), .A4(n88122), .ZN(
        n88105) );
  NAND2_X1 U73688 ( .A1(n88123), .A2(n88124), .ZN(n88122) );
  AOI22_X1 U73689 ( .A1(n105763), .A2(n109993), .B1(n105762), .B2(n109996), 
        .ZN(n88124) );
  AOI22_X1 U73690 ( .A1(n86363), .A2(n109997), .B1(n105760), .B2(n109999), 
        .ZN(n88123) );
  NAND2_X1 U73691 ( .A1(n88125), .A2(n88126), .ZN(n88121) );
  AOI22_X1 U73692 ( .A1(n105759), .A2(n109998), .B1(n86368), .B2(n109994), 
        .ZN(n88126) );
  AOI22_X1 U73693 ( .A1(n105757), .A2(n110000), .B1(n105756), .B2(n109995), 
        .ZN(n88125) );
  NAND2_X1 U73694 ( .A1(n88127), .A2(n88128), .ZN(n88120) );
  AOI22_X1 U73695 ( .A1(n105755), .A2(n73097), .B1(n105754), .B2(n73096), .ZN(
        n88128) );
  AOI22_X1 U73696 ( .A1(n105753), .A2(n73099), .B1(n105752), .B2(n110001), 
        .ZN(n88127) );
  NAND2_X1 U73697 ( .A1(n88129), .A2(n88130), .ZN(n88119) );
  AOI22_X1 U73698 ( .A1(n105751), .A2(n109986), .B1(n105750), .B2(n109991), 
        .ZN(n88130) );
  AOI22_X1 U73699 ( .A1(n105749), .A2(n73094), .B1(n105748), .B2(n109989), 
        .ZN(n88129) );
  NAND2_X1 U73700 ( .A1(n88131), .A2(n88132), .ZN(n88103) );
  NOR4_X1 U73701 ( .A1(n88133), .A2(n88134), .A3(n88135), .A4(n88136), .ZN(
        n88132) );
  NAND2_X1 U73702 ( .A1(n88137), .A2(n88138), .ZN(n88136) );
  AOI22_X1 U73703 ( .A1(n105747), .A2(n109919), .B1(n105746), .B2(n109921), 
        .ZN(n88138) );
  AOI22_X1 U73704 ( .A1(n105745), .A2(n73012), .B1(n105744), .B2(n109920), 
        .ZN(n88137) );
  NAND2_X1 U73705 ( .A1(n88139), .A2(n88140), .ZN(n88135) );
  AOI22_X1 U73706 ( .A1(n105743), .A2(n73016), .B1(n105742), .B2(n73018), .ZN(
        n88140) );
  AOI22_X1 U73707 ( .A1(n105741), .A2(n109927), .B1(n86400), .B2(n109928), 
        .ZN(n88139) );
  NAND2_X1 U73708 ( .A1(n88141), .A2(n88142), .ZN(n88134) );
  AOI22_X1 U73709 ( .A1(n86403), .A2(n109924), .B1(n105738), .B2(n109926), 
        .ZN(n88142) );
  AOI22_X1 U73710 ( .A1(n105737), .A2(n73017), .B1(n105736), .B2(n109925), 
        .ZN(n88141) );
  NAND2_X1 U73711 ( .A1(n88143), .A2(n88144), .ZN(n88133) );
  AOI22_X1 U73712 ( .A1(n105735), .A2(n109933), .B1(n105734), .B2(n73023), 
        .ZN(n88144) );
  AOI22_X1 U73713 ( .A1(n86411), .A2(n109932), .B1(n105732), .B2(n73021), .ZN(
        n88143) );
  NOR4_X1 U73714 ( .A1(n88145), .A2(n88146), .A3(n88147), .A4(n88148), .ZN(
        n88131) );
  NAND2_X1 U73715 ( .A1(n88149), .A2(n88150), .ZN(n88148) );
  AOI22_X1 U73716 ( .A1(n105731), .A2(n109914), .B1(n105730), .B2(n109905), 
        .ZN(n88150) );
  AOI22_X1 U73717 ( .A1(n105729), .A2(n109907), .B1(n105728), .B2(n72995), 
        .ZN(n88149) );
  NAND2_X1 U73718 ( .A1(n88151), .A2(n88152), .ZN(n88147) );
  AOI22_X1 U73719 ( .A1(n105727), .A2(n109912), .B1(n86426), .B2(n109916), 
        .ZN(n88152) );
  AOI22_X1 U73720 ( .A1(n105725), .A2(n109918), .B1(n86428), .B2(n109915), 
        .ZN(n88151) );
  NAND2_X1 U73721 ( .A1(n88153), .A2(n88154), .ZN(n88146) );
  AOI22_X1 U73722 ( .A1(n105723), .A2(n73004), .B1(n105722), .B2(n109911), 
        .ZN(n88154) );
  AOI22_X1 U73723 ( .A1(n105721), .A2(n109913), .B1(n105720), .B2(n109917), 
        .ZN(n88153) );
  NAND2_X1 U73724 ( .A1(n88155), .A2(n88156), .ZN(n88145) );
  AOI22_X1 U73725 ( .A1(n105719), .A2(n109923), .B1(n105718), .B2(n73008), 
        .ZN(n88156) );
  AOI22_X1 U73726 ( .A1(n105717), .A2(n73006), .B1(n105716), .B2(n109922), 
        .ZN(n88155) );
  NAND2_X1 U73727 ( .A1(n88157), .A2(n88158), .ZN(n88102) );
  NOR4_X1 U73728 ( .A1(n88159), .A2(n88160), .A3(n88161), .A4(n88162), .ZN(
        n88158) );
  NAND2_X1 U73729 ( .A1(n88163), .A2(n88164), .ZN(n88162) );
  AOI22_X1 U73730 ( .A1(n105715), .A2(n73046), .B1(n86450), .B2(n109943), .ZN(
        n88164) );
  AOI22_X1 U73731 ( .A1(n105713), .A2(n109947), .B1(n105712), .B2(n109946), 
        .ZN(n88163) );
  NAND2_X1 U73732 ( .A1(n88165), .A2(n88166), .ZN(n88161) );
  AOI22_X1 U73733 ( .A1(n105711), .A2(n109952), .B1(n105710), .B2(n109951), 
        .ZN(n88166) );
  AOI22_X1 U73734 ( .A1(n105709), .A2(n109942), .B1(n86458), .B2(n109944), 
        .ZN(n88165) );
  NAND2_X1 U73735 ( .A1(n88167), .A2(n88168), .ZN(n88160) );
  AOI22_X1 U73736 ( .A1(n105707), .A2(n109953), .B1(n105706), .B2(n109949), 
        .ZN(n88168) );
  AOI22_X1 U73737 ( .A1(n105705), .A2(n73050), .B1(n105704), .B2(n73052), .ZN(
        n88167) );
  NAND2_X1 U73738 ( .A1(n88169), .A2(n88170), .ZN(n88159) );
  AOI22_X1 U73739 ( .A1(n86467), .A2(n109956), .B1(n105702), .B2(n73058), .ZN(
        n88170) );
  AOI22_X1 U73740 ( .A1(n105701), .A2(n109948), .B1(n105700), .B2(n109950), 
        .ZN(n88169) );
  NOR4_X1 U73741 ( .A1(n88171), .A2(n88172), .A3(n88173), .A4(n88174), .ZN(
        n88157) );
  NAND2_X1 U73742 ( .A1(n88175), .A2(n88176), .ZN(n88174) );
  AOI22_X1 U73743 ( .A1(n105699), .A2(n109931), .B1(n105698), .B2(n109936), 
        .ZN(n88176) );
  AOI22_X1 U73744 ( .A1(n105697), .A2(n109930), .B1(n105696), .B2(n73026), 
        .ZN(n88175) );
  NAND2_X1 U73745 ( .A1(n88177), .A2(n88178), .ZN(n88173) );
  AOI22_X1 U73746 ( .A1(n105695), .A2(n73035), .B1(n105694), .B2(n109938), 
        .ZN(n88178) );
  AOI22_X1 U73747 ( .A1(n105693), .A2(n109939), .B1(n105692), .B2(n109929), 
        .ZN(n88177) );
  NAND2_X1 U73748 ( .A1(n88179), .A2(n88180), .ZN(n88172) );
  AOI22_X1 U73749 ( .A1(n105691), .A2(n109937), .B1(n86490), .B2(n109941), 
        .ZN(n88180) );
  AOI22_X1 U73750 ( .A1(n105689), .A2(n109935), .B1(n105688), .B2(n109940), 
        .ZN(n88179) );
  NAND2_X1 U73751 ( .A1(n88181), .A2(n88182), .ZN(n88171) );
  AOI22_X1 U73752 ( .A1(n105687), .A2(n73040), .B1(n105686), .B2(n109945), 
        .ZN(n88182) );
  AOI22_X1 U73753 ( .A1(n105685), .A2(n73038), .B1(n105684), .B2(n109934), 
        .ZN(n88181) );
  NAND2_X1 U73754 ( .A1(n88183), .A2(n88184), .ZN(n88101) );
  NOR4_X1 U73755 ( .A1(n88185), .A2(n88186), .A3(n88187), .A4(n88188), .ZN(
        n88184) );
  NAND2_X1 U73756 ( .A1(n88189), .A2(n88190), .ZN(n88188) );
  AOI22_X1 U73757 ( .A1(n105683), .A2(n109974), .B1(n105682), .B2(n109973), 
        .ZN(n88190) );
  AOI22_X1 U73758 ( .A1(n105681), .A2(n73074), .B1(n105680), .B2(n109971), 
        .ZN(n88189) );
  NAND2_X1 U73759 ( .A1(n88191), .A2(n88192), .ZN(n88187) );
  AOI22_X1 U73760 ( .A1(n105679), .A2(n109969), .B1(n105678), .B2(n109972), 
        .ZN(n88192) );
  AOI22_X1 U73761 ( .A1(n86515), .A2(n73080), .B1(n86516), .B2(n109970), .ZN(
        n88191) );
  NAND2_X1 U73762 ( .A1(n88193), .A2(n88194), .ZN(n88186) );
  AOI22_X1 U73763 ( .A1(n86519), .A2(n109980), .B1(n86520), .B2(n73086), .ZN(
        n88194) );
  AOI22_X1 U73764 ( .A1(n86521), .A2(n109978), .B1(n86522), .B2(n109979), .ZN(
        n88193) );
  NAND2_X1 U73765 ( .A1(n88195), .A2(n88196), .ZN(n88185) );
  AOI22_X1 U73766 ( .A1(n105676), .A2(n109975), .B1(n86526), .B2(n109977), 
        .ZN(n88196) );
  AOI22_X1 U73767 ( .A1(n86527), .A2(n109981), .B1(n86528), .B2(n109976), .ZN(
        n88195) );
  NOR4_X1 U73768 ( .A1(n88197), .A2(n88198), .A3(n88199), .A4(n88200), .ZN(
        n88183) );
  NAND2_X1 U73769 ( .A1(n88201), .A2(n88202), .ZN(n88200) );
  AOI22_X1 U73770 ( .A1(n105675), .A2(n109955), .B1(n105674), .B2(n109959), 
        .ZN(n88202) );
  AOI22_X1 U73771 ( .A1(n105673), .A2(n109958), .B1(n105672), .B2(n73057), 
        .ZN(n88201) );
  NAND2_X1 U73772 ( .A1(n88203), .A2(n88204), .ZN(n88199) );
  AOI22_X1 U73773 ( .A1(n105671), .A2(n109965), .B1(n105670), .B2(n109954), 
        .ZN(n88204) );
  AOI22_X1 U73774 ( .A1(n105669), .A2(n109957), .B1(n105668), .B2(n109962), 
        .ZN(n88203) );
  NAND2_X1 U73775 ( .A1(n88205), .A2(n88206), .ZN(n88198) );
  AOI22_X1 U73776 ( .A1(n105667), .A2(n109961), .B1(n105666), .B2(n109966), 
        .ZN(n88206) );
  AOI22_X1 U73777 ( .A1(n86549), .A2(n109968), .B1(n105664), .B2(n109964), 
        .ZN(n88205) );
  NAND2_X1 U73778 ( .A1(n88207), .A2(n88208), .ZN(n88197) );
  AOI22_X1 U73779 ( .A1(n105663), .A2(n73075), .B1(n105662), .B2(n109960), 
        .ZN(n88208) );
  AOI22_X1 U73780 ( .A1(n105661), .A2(n109963), .B1(n105660), .B2(n109967), 
        .ZN(n88207) );
  AOI21_X1 U73781 ( .B1(n86302), .B2(n88210), .A(n88211), .ZN(n88209) );
  OAI21_X1 U73782 ( .B1(n88212), .B2(n105787), .A(n88213), .ZN(n88211) );
  OAI21_X1 U73783 ( .B1(n88214), .B2(n88215), .A(n105786), .ZN(n88213) );
  OAI21_X1 U73784 ( .B1(n109889), .B2(n86311), .A(n88216), .ZN(n88215) );
  AOI22_X1 U73785 ( .A1(n86313), .A2(n72964), .B1(n105784), .B2(n109887), .ZN(
        n88216) );
  NAND2_X1 U73786 ( .A1(n88217), .A2(n88218), .ZN(n88214) );
  AOI22_X1 U73787 ( .A1(n105783), .A2(n109885), .B1(n105782), .B2(n109890), 
        .ZN(n88218) );
  AOI22_X1 U73788 ( .A1(n105781), .A2(n109888), .B1(n105780), .B2(n109886), 
        .ZN(n88217) );
  NOR4_X1 U73789 ( .A1(n88219), .A2(n88220), .A3(n88221), .A4(n88222), .ZN(
        n88212) );
  NAND2_X1 U73790 ( .A1(n88223), .A2(n88224), .ZN(n88222) );
  NOR4_X1 U73791 ( .A1(n88225), .A2(n88226), .A3(n88227), .A4(n88228), .ZN(
        n88224) );
  NAND2_X1 U73792 ( .A1(n88229), .A2(n88230), .ZN(n88228) );
  AOI22_X1 U73793 ( .A1(n105779), .A2(n109866), .B1(n105778), .B2(n109867), 
        .ZN(n88230) );
  AOI22_X1 U73794 ( .A1(n105777), .A2(n109875), .B1(n105776), .B2(n109873), 
        .ZN(n88229) );
  NAND2_X1 U73795 ( .A1(n88231), .A2(n88232), .ZN(n88227) );
  AOI22_X1 U73796 ( .A1(n105775), .A2(n72833), .B1(n105774), .B2(n109870), 
        .ZN(n88232) );
  AOI22_X1 U73797 ( .A1(n105773), .A2(n72937), .B1(n105772), .B2(n109786), 
        .ZN(n88231) );
  NAND2_X1 U73798 ( .A1(n88233), .A2(n88234), .ZN(n88226) );
  AOI22_X1 U73799 ( .A1(n105771), .A2(n109790), .B1(n105770), .B2(n72837), 
        .ZN(n88234) );
  AOI22_X1 U73800 ( .A1(n105769), .A2(n109871), .B1(n105768), .B2(n109868), 
        .ZN(n88233) );
  NAND2_X1 U73801 ( .A1(n88235), .A2(n88236), .ZN(n88225) );
  AOI22_X1 U73802 ( .A1(n105767), .A2(n109788), .B1(n105766), .B2(n109792), 
        .ZN(n88236) );
  AOI22_X1 U73803 ( .A1(n105765), .A2(n109791), .B1(n105764), .B2(n72839), 
        .ZN(n88235) );
  NOR4_X1 U73804 ( .A1(n88237), .A2(n88238), .A3(n88239), .A4(n88240), .ZN(
        n88223) );
  NAND2_X1 U73805 ( .A1(n88241), .A2(n88242), .ZN(n88240) );
  AOI22_X1 U73806 ( .A1(n105763), .A2(n109876), .B1(n105762), .B2(n109879), 
        .ZN(n88242) );
  AOI22_X1 U73807 ( .A1(n105761), .A2(n109880), .B1(n105760), .B2(n109882), 
        .ZN(n88241) );
  NAND2_X1 U73808 ( .A1(n88243), .A2(n88244), .ZN(n88239) );
  AOI22_X1 U73809 ( .A1(n105759), .A2(n109881), .B1(n105758), .B2(n109877), 
        .ZN(n88244) );
  AOI22_X1 U73810 ( .A1(n105757), .A2(n109883), .B1(n105756), .B2(n109878), 
        .ZN(n88243) );
  NAND2_X1 U73811 ( .A1(n88245), .A2(n88246), .ZN(n88238) );
  AOI22_X1 U73812 ( .A1(n105755), .A2(n72947), .B1(n105754), .B2(n72946), .ZN(
        n88246) );
  AOI22_X1 U73813 ( .A1(n105753), .A2(n72949), .B1(n105752), .B2(n109884), 
        .ZN(n88245) );
  NAND2_X1 U73814 ( .A1(n88247), .A2(n88248), .ZN(n88237) );
  AOI22_X1 U73815 ( .A1(n105751), .A2(n109869), .B1(n105750), .B2(n109874), 
        .ZN(n88248) );
  AOI22_X1 U73816 ( .A1(n105749), .A2(n72944), .B1(n105748), .B2(n109872), 
        .ZN(n88247) );
  NAND2_X1 U73817 ( .A1(n88249), .A2(n88250), .ZN(n88221) );
  NOR4_X1 U73818 ( .A1(n88251), .A2(n88252), .A3(n88253), .A4(n88254), .ZN(
        n88250) );
  NAND2_X1 U73819 ( .A1(n88255), .A2(n88256), .ZN(n88254) );
  AOI22_X1 U73820 ( .A1(n105747), .A2(n109801), .B1(n105746), .B2(n109803), 
        .ZN(n88256) );
  AOI22_X1 U73821 ( .A1(n105745), .A2(n72862), .B1(n105744), .B2(n109802), 
        .ZN(n88255) );
  NAND2_X1 U73822 ( .A1(n88257), .A2(n88258), .ZN(n88253) );
  AOI22_X1 U73823 ( .A1(n105743), .A2(n72866), .B1(n105742), .B2(n72868), .ZN(
        n88258) );
  AOI22_X1 U73824 ( .A1(n105741), .A2(n109809), .B1(n105740), .B2(n109810), 
        .ZN(n88257) );
  NAND2_X1 U73825 ( .A1(n88259), .A2(n88260), .ZN(n88252) );
  AOI22_X1 U73826 ( .A1(n105739), .A2(n109806), .B1(n105738), .B2(n109808), 
        .ZN(n88260) );
  AOI22_X1 U73827 ( .A1(n105737), .A2(n109811), .B1(n105736), .B2(n109807), 
        .ZN(n88259) );
  NAND2_X1 U73828 ( .A1(n88261), .A2(n88262), .ZN(n88251) );
  AOI22_X1 U73829 ( .A1(n105735), .A2(n109816), .B1(n105734), .B2(n72873), 
        .ZN(n88262) );
  AOI22_X1 U73830 ( .A1(n105733), .A2(n109815), .B1(n105732), .B2(n72871), 
        .ZN(n88261) );
  NOR4_X1 U73831 ( .A1(n88263), .A2(n88264), .A3(n88265), .A4(n88266), .ZN(
        n88249) );
  NAND2_X1 U73832 ( .A1(n88267), .A2(n88268), .ZN(n88266) );
  AOI22_X1 U73833 ( .A1(n105731), .A2(n109796), .B1(n105730), .B2(n109787), 
        .ZN(n88268) );
  AOI22_X1 U73834 ( .A1(n105729), .A2(n109789), .B1(n105728), .B2(n72845), 
        .ZN(n88267) );
  NAND2_X1 U73835 ( .A1(n88269), .A2(n88270), .ZN(n88265) );
  AOI22_X1 U73836 ( .A1(n105727), .A2(n109794), .B1(n105726), .B2(n109798), 
        .ZN(n88270) );
  AOI22_X1 U73837 ( .A1(n105725), .A2(n109800), .B1(n105724), .B2(n109797), 
        .ZN(n88269) );
  NAND2_X1 U73838 ( .A1(n88271), .A2(n88272), .ZN(n88264) );
  AOI22_X1 U73839 ( .A1(n105723), .A2(n72854), .B1(n105722), .B2(n109793), 
        .ZN(n88272) );
  AOI22_X1 U73840 ( .A1(n105721), .A2(n109795), .B1(n105720), .B2(n109799), 
        .ZN(n88271) );
  NAND2_X1 U73841 ( .A1(n88273), .A2(n88274), .ZN(n88263) );
  AOI22_X1 U73842 ( .A1(n105719), .A2(n109805), .B1(n105718), .B2(n72858), 
        .ZN(n88274) );
  AOI22_X1 U73843 ( .A1(n105717), .A2(n72856), .B1(n105716), .B2(n109804), 
        .ZN(n88273) );
  NAND2_X1 U73844 ( .A1(n88275), .A2(n88276), .ZN(n88220) );
  NOR4_X1 U73845 ( .A1(n88277), .A2(n88278), .A3(n88279), .A4(n88280), .ZN(
        n88276) );
  NAND2_X1 U73846 ( .A1(n88281), .A2(n88282), .ZN(n88280) );
  AOI22_X1 U73847 ( .A1(n105715), .A2(n72896), .B1(n105714), .B2(n109826), 
        .ZN(n88282) );
  AOI22_X1 U73848 ( .A1(n105713), .A2(n109830), .B1(n105712), .B2(n109829), 
        .ZN(n88281) );
  NAND2_X1 U73849 ( .A1(n88283), .A2(n88284), .ZN(n88279) );
  AOI22_X1 U73850 ( .A1(n105711), .A2(n109835), .B1(n105710), .B2(n109834), 
        .ZN(n88284) );
  AOI22_X1 U73851 ( .A1(n105709), .A2(n109825), .B1(n86458), .B2(n109827), 
        .ZN(n88283) );
  NAND2_X1 U73852 ( .A1(n88285), .A2(n88286), .ZN(n88278) );
  AOI22_X1 U73853 ( .A1(n105707), .A2(n109836), .B1(n105706), .B2(n109832), 
        .ZN(n88286) );
  AOI22_X1 U73854 ( .A1(n105705), .A2(n72900), .B1(n105704), .B2(n72902), .ZN(
        n88285) );
  NAND2_X1 U73855 ( .A1(n88287), .A2(n88288), .ZN(n88277) );
  AOI22_X1 U73856 ( .A1(n105703), .A2(n109839), .B1(n105702), .B2(n72908), 
        .ZN(n88288) );
  AOI22_X1 U73857 ( .A1(n105701), .A2(n109831), .B1(n105700), .B2(n109833), 
        .ZN(n88287) );
  NOR4_X1 U73858 ( .A1(n88289), .A2(n88290), .A3(n88291), .A4(n88292), .ZN(
        n88275) );
  NAND2_X1 U73859 ( .A1(n88293), .A2(n88294), .ZN(n88292) );
  AOI22_X1 U73860 ( .A1(n105699), .A2(n109814), .B1(n105698), .B2(n109819), 
        .ZN(n88294) );
  AOI22_X1 U73861 ( .A1(n105697), .A2(n109813), .B1(n105696), .B2(n72876), 
        .ZN(n88293) );
  NAND2_X1 U73862 ( .A1(n88295), .A2(n88296), .ZN(n88291) );
  AOI22_X1 U73863 ( .A1(n105695), .A2(n72885), .B1(n105694), .B2(n109821), 
        .ZN(n88296) );
  AOI22_X1 U73864 ( .A1(n105693), .A2(n109822), .B1(n105692), .B2(n109812), 
        .ZN(n88295) );
  NAND2_X1 U73865 ( .A1(n88297), .A2(n88298), .ZN(n88290) );
  AOI22_X1 U73866 ( .A1(n105691), .A2(n109820), .B1(n105690), .B2(n109824), 
        .ZN(n88298) );
  AOI22_X1 U73867 ( .A1(n105689), .A2(n109818), .B1(n105688), .B2(n109823), 
        .ZN(n88297) );
  NAND2_X1 U73868 ( .A1(n88299), .A2(n88300), .ZN(n88289) );
  AOI22_X1 U73869 ( .A1(n105687), .A2(n72890), .B1(n105686), .B2(n109828), 
        .ZN(n88300) );
  AOI22_X1 U73870 ( .A1(n105685), .A2(n72888), .B1(n105684), .B2(n109817), 
        .ZN(n88299) );
  NAND2_X1 U73871 ( .A1(n88301), .A2(n88302), .ZN(n88219) );
  NOR4_X1 U73872 ( .A1(n88303), .A2(n88304), .A3(n88305), .A4(n88306), .ZN(
        n88302) );
  NAND2_X1 U73873 ( .A1(n88307), .A2(n88308), .ZN(n88306) );
  AOI22_X1 U73874 ( .A1(n105683), .A2(n109857), .B1(n105682), .B2(n109856), 
        .ZN(n88308) );
  AOI22_X1 U73875 ( .A1(n105681), .A2(n72924), .B1(n105680), .B2(n109854), 
        .ZN(n88307) );
  NAND2_X1 U73876 ( .A1(n88309), .A2(n88310), .ZN(n88305) );
  AOI22_X1 U73877 ( .A1(n105679), .A2(n109852), .B1(n105678), .B2(n109855), 
        .ZN(n88310) );
  AOI22_X1 U73878 ( .A1(n86515), .A2(n72930), .B1(n105677), .B2(n109853), .ZN(
        n88309) );
  NAND2_X1 U73879 ( .A1(n88311), .A2(n88312), .ZN(n88304) );
  AOI22_X1 U73880 ( .A1(n86519), .A2(n109863), .B1(n86520), .B2(n72936), .ZN(
        n88312) );
  AOI22_X1 U73881 ( .A1(n86521), .A2(n109861), .B1(n86522), .B2(n109862), .ZN(
        n88311) );
  NAND2_X1 U73882 ( .A1(n88313), .A2(n88314), .ZN(n88303) );
  AOI22_X1 U73883 ( .A1(n105676), .A2(n109858), .B1(n86526), .B2(n109860), 
        .ZN(n88314) );
  AOI22_X1 U73884 ( .A1(n86527), .A2(n109864), .B1(n86528), .B2(n109859), .ZN(
        n88313) );
  NOR4_X1 U73885 ( .A1(n88315), .A2(n88316), .A3(n88317), .A4(n88318), .ZN(
        n88301) );
  NAND2_X1 U73886 ( .A1(n88319), .A2(n88320), .ZN(n88318) );
  AOI22_X1 U73887 ( .A1(n105675), .A2(n109838), .B1(n105674), .B2(n109842), 
        .ZN(n88320) );
  AOI22_X1 U73888 ( .A1(n105673), .A2(n109841), .B1(n105672), .B2(n72907), 
        .ZN(n88319) );
  NAND2_X1 U73889 ( .A1(n88321), .A2(n88322), .ZN(n88317) );
  AOI22_X1 U73890 ( .A1(n105671), .A2(n109848), .B1(n105670), .B2(n109837), 
        .ZN(n88322) );
  AOI22_X1 U73891 ( .A1(n105669), .A2(n109840), .B1(n105668), .B2(n109845), 
        .ZN(n88321) );
  NAND2_X1 U73892 ( .A1(n88323), .A2(n88324), .ZN(n88316) );
  AOI22_X1 U73893 ( .A1(n105667), .A2(n109844), .B1(n105666), .B2(n109849), 
        .ZN(n88324) );
  AOI22_X1 U73894 ( .A1(n105665), .A2(n109851), .B1(n86550), .B2(n109847), 
        .ZN(n88323) );
  NAND2_X1 U73895 ( .A1(n88325), .A2(n88326), .ZN(n88315) );
  AOI22_X1 U73896 ( .A1(n105663), .A2(n72925), .B1(n105662), .B2(n109843), 
        .ZN(n88326) );
  AOI22_X1 U73897 ( .A1(n105661), .A2(n109846), .B1(n105660), .B2(n109850), 
        .ZN(n88325) );
  AOI21_X1 U73898 ( .B1(n86302), .B2(n88328), .A(n88329), .ZN(n88327) );
  OAI21_X1 U73899 ( .B1(n88330), .B2(n105787), .A(n88331), .ZN(n88329) );
  OAI21_X1 U73900 ( .B1(n88332), .B2(n88333), .A(n105786), .ZN(n88331) );
  OAI21_X1 U73901 ( .B1(n108263), .B2(n105785), .A(n88334), .ZN(n88333) );
  AOI22_X1 U73902 ( .A1(n86313), .A2(n70860), .B1(n105784), .B2(n108261), .ZN(
        n88334) );
  NAND2_X1 U73903 ( .A1(n88335), .A2(n88336), .ZN(n88332) );
  AOI22_X1 U73904 ( .A1(n105783), .A2(n108259), .B1(n105782), .B2(n108264), 
        .ZN(n88336) );
  AOI22_X1 U73905 ( .A1(n105781), .A2(n108262), .B1(n105780), .B2(n108260), 
        .ZN(n88335) );
  NOR4_X1 U73906 ( .A1(n88337), .A2(n88338), .A3(n88339), .A4(n88340), .ZN(
        n88330) );
  NAND2_X1 U73907 ( .A1(n88341), .A2(n88342), .ZN(n88340) );
  NOR4_X1 U73908 ( .A1(n88343), .A2(n88344), .A3(n88345), .A4(n88346), .ZN(
        n88342) );
  NAND2_X1 U73909 ( .A1(n88347), .A2(n88348), .ZN(n88346) );
  AOI22_X1 U73910 ( .A1(n105779), .A2(n108240), .B1(n105778), .B2(n108241), 
        .ZN(n88348) );
  AOI22_X1 U73911 ( .A1(n105777), .A2(n108249), .B1(n105776), .B2(n108247), 
        .ZN(n88347) );
  NAND2_X1 U73912 ( .A1(n88349), .A2(n88350), .ZN(n88345) );
  AOI22_X1 U73913 ( .A1(n105775), .A2(n70729), .B1(n105774), .B2(n108244), 
        .ZN(n88350) );
  AOI22_X1 U73914 ( .A1(n105773), .A2(n70833), .B1(n105772), .B2(n108160), 
        .ZN(n88349) );
  NAND2_X1 U73915 ( .A1(n88351), .A2(n88352), .ZN(n88344) );
  AOI22_X1 U73916 ( .A1(n105771), .A2(n108164), .B1(n86346), .B2(n70733), .ZN(
        n88352) );
  AOI22_X1 U73917 ( .A1(n105769), .A2(n108245), .B1(n105768), .B2(n108242), 
        .ZN(n88351) );
  NAND2_X1 U73918 ( .A1(n88353), .A2(n88354), .ZN(n88343) );
  AOI22_X1 U73919 ( .A1(n105767), .A2(n108162), .B1(n105766), .B2(n108166), 
        .ZN(n88354) );
  AOI22_X1 U73920 ( .A1(n105765), .A2(n108165), .B1(n105764), .B2(n70735), 
        .ZN(n88353) );
  NOR4_X1 U73921 ( .A1(n88355), .A2(n88356), .A3(n88357), .A4(n88358), .ZN(
        n88341) );
  NAND2_X1 U73922 ( .A1(n88359), .A2(n88360), .ZN(n88358) );
  AOI22_X1 U73923 ( .A1(n105763), .A2(n108250), .B1(n105762), .B2(n108253), 
        .ZN(n88360) );
  AOI22_X1 U73924 ( .A1(n86363), .A2(n108254), .B1(n105760), .B2(n108256), 
        .ZN(n88359) );
  NAND2_X1 U73925 ( .A1(n88361), .A2(n88362), .ZN(n88357) );
  AOI22_X1 U73926 ( .A1(n105759), .A2(n108255), .B1(n86368), .B2(n108251), 
        .ZN(n88362) );
  AOI22_X1 U73927 ( .A1(n105757), .A2(n108257), .B1(n105756), .B2(n108252), 
        .ZN(n88361) );
  NAND2_X1 U73928 ( .A1(n88363), .A2(n88364), .ZN(n88356) );
  AOI22_X1 U73929 ( .A1(n105755), .A2(n70843), .B1(n105754), .B2(n70842), .ZN(
        n88364) );
  AOI22_X1 U73930 ( .A1(n105753), .A2(n70845), .B1(n105752), .B2(n108258), 
        .ZN(n88363) );
  NAND2_X1 U73931 ( .A1(n88365), .A2(n88366), .ZN(n88355) );
  AOI22_X1 U73932 ( .A1(n105751), .A2(n108243), .B1(n105750), .B2(n108248), 
        .ZN(n88366) );
  AOI22_X1 U73933 ( .A1(n105749), .A2(n70840), .B1(n105748), .B2(n108246), 
        .ZN(n88365) );
  NAND2_X1 U73934 ( .A1(n88367), .A2(n88368), .ZN(n88339) );
  NOR4_X1 U73935 ( .A1(n88369), .A2(n88370), .A3(n88371), .A4(n88372), .ZN(
        n88368) );
  NAND2_X1 U73936 ( .A1(n88373), .A2(n88374), .ZN(n88372) );
  AOI22_X1 U73937 ( .A1(n105747), .A2(n108175), .B1(n105746), .B2(n108177), 
        .ZN(n88374) );
  AOI22_X1 U73938 ( .A1(n105745), .A2(n70758), .B1(n105744), .B2(n108176), 
        .ZN(n88373) );
  NAND2_X1 U73939 ( .A1(n88375), .A2(n88376), .ZN(n88371) );
  AOI22_X1 U73940 ( .A1(n105743), .A2(n70762), .B1(n105742), .B2(n70764), .ZN(
        n88376) );
  AOI22_X1 U73941 ( .A1(n105741), .A2(n108183), .B1(n86400), .B2(n108184), 
        .ZN(n88375) );
  NAND2_X1 U73942 ( .A1(n88377), .A2(n88378), .ZN(n88370) );
  AOI22_X1 U73943 ( .A1(n86403), .A2(n108180), .B1(n105738), .B2(n108182), 
        .ZN(n88378) );
  AOI22_X1 U73944 ( .A1(n105737), .A2(n108185), .B1(n105736), .B2(n108181), 
        .ZN(n88377) );
  NAND2_X1 U73945 ( .A1(n88379), .A2(n88380), .ZN(n88369) );
  AOI22_X1 U73946 ( .A1(n105735), .A2(n108190), .B1(n105734), .B2(n70769), 
        .ZN(n88380) );
  AOI22_X1 U73947 ( .A1(n86411), .A2(n108189), .B1(n105732), .B2(n70767), .ZN(
        n88379) );
  NOR4_X1 U73948 ( .A1(n88381), .A2(n88382), .A3(n88383), .A4(n88384), .ZN(
        n88367) );
  NAND2_X1 U73949 ( .A1(n88385), .A2(n88386), .ZN(n88384) );
  AOI22_X1 U73950 ( .A1(n105731), .A2(n108170), .B1(n105730), .B2(n108161), 
        .ZN(n88386) );
  AOI22_X1 U73951 ( .A1(n105729), .A2(n108163), .B1(n105728), .B2(n70741), 
        .ZN(n88385) );
  NAND2_X1 U73952 ( .A1(n88387), .A2(n88388), .ZN(n88383) );
  AOI22_X1 U73953 ( .A1(n105727), .A2(n108168), .B1(n86426), .B2(n108172), 
        .ZN(n88388) );
  AOI22_X1 U73954 ( .A1(n105725), .A2(n108174), .B1(n86428), .B2(n108171), 
        .ZN(n88387) );
  NAND2_X1 U73955 ( .A1(n88389), .A2(n88390), .ZN(n88382) );
  AOI22_X1 U73956 ( .A1(n105723), .A2(n70750), .B1(n105722), .B2(n108167), 
        .ZN(n88390) );
  AOI22_X1 U73957 ( .A1(n105721), .A2(n108169), .B1(n105720), .B2(n108173), 
        .ZN(n88389) );
  NAND2_X1 U73958 ( .A1(n88391), .A2(n88392), .ZN(n88381) );
  AOI22_X1 U73959 ( .A1(n105719), .A2(n108179), .B1(n105718), .B2(n70754), 
        .ZN(n88392) );
  AOI22_X1 U73960 ( .A1(n105717), .A2(n70752), .B1(n105716), .B2(n108178), 
        .ZN(n88391) );
  NAND2_X1 U73961 ( .A1(n88393), .A2(n88394), .ZN(n88338) );
  NOR4_X1 U73962 ( .A1(n88395), .A2(n88396), .A3(n88397), .A4(n88398), .ZN(
        n88394) );
  NAND2_X1 U73963 ( .A1(n88399), .A2(n88400), .ZN(n88398) );
  AOI22_X1 U73964 ( .A1(n105715), .A2(n70792), .B1(n86450), .B2(n108200), .ZN(
        n88400) );
  AOI22_X1 U73965 ( .A1(n105713), .A2(n108204), .B1(n105712), .B2(n108203), 
        .ZN(n88399) );
  NAND2_X1 U73966 ( .A1(n88401), .A2(n88402), .ZN(n88397) );
  AOI22_X1 U73967 ( .A1(n105711), .A2(n108209), .B1(n105710), .B2(n108208), 
        .ZN(n88402) );
  AOI22_X1 U73968 ( .A1(n105709), .A2(n108199), .B1(n86458), .B2(n108201), 
        .ZN(n88401) );
  NAND2_X1 U73969 ( .A1(n88403), .A2(n88404), .ZN(n88396) );
  AOI22_X1 U73970 ( .A1(n105707), .A2(n108210), .B1(n105706), .B2(n108206), 
        .ZN(n88404) );
  AOI22_X1 U73971 ( .A1(n105705), .A2(n70796), .B1(n105704), .B2(n70798), .ZN(
        n88403) );
  NAND2_X1 U73972 ( .A1(n88405), .A2(n88406), .ZN(n88395) );
  AOI22_X1 U73973 ( .A1(n86467), .A2(n108213), .B1(n105702), .B2(n70804), .ZN(
        n88406) );
  AOI22_X1 U73974 ( .A1(n105701), .A2(n108205), .B1(n105700), .B2(n108207), 
        .ZN(n88405) );
  NOR4_X1 U73975 ( .A1(n88407), .A2(n88408), .A3(n88409), .A4(n88410), .ZN(
        n88393) );
  NAND2_X1 U73976 ( .A1(n88411), .A2(n88412), .ZN(n88410) );
  AOI22_X1 U73977 ( .A1(n105699), .A2(n108188), .B1(n105698), .B2(n108193), 
        .ZN(n88412) );
  AOI22_X1 U73978 ( .A1(n105697), .A2(n108187), .B1(n105696), .B2(n70772), 
        .ZN(n88411) );
  NAND2_X1 U73979 ( .A1(n88413), .A2(n88414), .ZN(n88409) );
  AOI22_X1 U73980 ( .A1(n105695), .A2(n70781), .B1(n86484), .B2(n108195), .ZN(
        n88414) );
  AOI22_X1 U73981 ( .A1(n105693), .A2(n108196), .B1(n105692), .B2(n108186), 
        .ZN(n88413) );
  NAND2_X1 U73982 ( .A1(n88415), .A2(n88416), .ZN(n88408) );
  AOI22_X1 U73983 ( .A1(n105691), .A2(n108194), .B1(n86490), .B2(n108198), 
        .ZN(n88416) );
  AOI22_X1 U73984 ( .A1(n105689), .A2(n108192), .B1(n105688), .B2(n108197), 
        .ZN(n88415) );
  NAND2_X1 U73985 ( .A1(n88417), .A2(n88418), .ZN(n88407) );
  AOI22_X1 U73986 ( .A1(n105687), .A2(n70786), .B1(n105686), .B2(n108202), 
        .ZN(n88418) );
  AOI22_X1 U73987 ( .A1(n105685), .A2(n70784), .B1(n105684), .B2(n108191), 
        .ZN(n88417) );
  NAND2_X1 U73988 ( .A1(n88419), .A2(n88420), .ZN(n88337) );
  NOR4_X1 U73989 ( .A1(n88421), .A2(n88422), .A3(n88423), .A4(n88424), .ZN(
        n88420) );
  NAND2_X1 U73990 ( .A1(n88425), .A2(n88426), .ZN(n88424) );
  AOI22_X1 U73991 ( .A1(n105683), .A2(n108231), .B1(n105682), .B2(n108230), 
        .ZN(n88426) );
  AOI22_X1 U73992 ( .A1(n105681), .A2(n70820), .B1(n105680), .B2(n108228), 
        .ZN(n88425) );
  NAND2_X1 U73993 ( .A1(n88427), .A2(n88428), .ZN(n88423) );
  AOI22_X1 U73994 ( .A1(n105679), .A2(n108226), .B1(n105678), .B2(n108229), 
        .ZN(n88428) );
  AOI22_X1 U73995 ( .A1(n86515), .A2(n70826), .B1(n86516), .B2(n108227), .ZN(
        n88427) );
  NAND2_X1 U73996 ( .A1(n88429), .A2(n88430), .ZN(n88422) );
  AOI22_X1 U73997 ( .A1(n86519), .A2(n108237), .B1(n86520), .B2(n70832), .ZN(
        n88430) );
  AOI22_X1 U73998 ( .A1(n86521), .A2(n108235), .B1(n86522), .B2(n108236), .ZN(
        n88429) );
  NAND2_X1 U73999 ( .A1(n88431), .A2(n88432), .ZN(n88421) );
  AOI22_X1 U74000 ( .A1(n105676), .A2(n108232), .B1(n86526), .B2(n108234), 
        .ZN(n88432) );
  AOI22_X1 U74001 ( .A1(n86527), .A2(n108238), .B1(n86528), .B2(n108233), .ZN(
        n88431) );
  NOR4_X1 U74002 ( .A1(n88433), .A2(n88434), .A3(n88435), .A4(n88436), .ZN(
        n88419) );
  NAND2_X1 U74003 ( .A1(n88437), .A2(n88438), .ZN(n88436) );
  AOI22_X1 U74004 ( .A1(n105675), .A2(n108212), .B1(n105674), .B2(n108216), 
        .ZN(n88438) );
  AOI22_X1 U74005 ( .A1(n105673), .A2(n108215), .B1(n105672), .B2(n70803), 
        .ZN(n88437) );
  NAND2_X1 U74006 ( .A1(n88439), .A2(n88440), .ZN(n88435) );
  AOI22_X1 U74007 ( .A1(n105671), .A2(n108222), .B1(n105670), .B2(n108211), 
        .ZN(n88440) );
  AOI22_X1 U74008 ( .A1(n105669), .A2(n108214), .B1(n105668), .B2(n108219), 
        .ZN(n88439) );
  NAND2_X1 U74009 ( .A1(n88441), .A2(n88442), .ZN(n88434) );
  AOI22_X1 U74010 ( .A1(n105667), .A2(n108218), .B1(n105666), .B2(n108223), 
        .ZN(n88442) );
  AOI22_X1 U74011 ( .A1(n86549), .A2(n108225), .B1(n105664), .B2(n108221), 
        .ZN(n88441) );
  NAND2_X1 U74012 ( .A1(n88443), .A2(n88444), .ZN(n88433) );
  AOI22_X1 U74013 ( .A1(n105663), .A2(n70821), .B1(n105662), .B2(n108217), 
        .ZN(n88444) );
  AOI22_X1 U74014 ( .A1(n105661), .A2(n108220), .B1(n105660), .B2(n108224), 
        .ZN(n88443) );
  AOI21_X1 U74015 ( .B1(n86302), .B2(n88446), .A(n88447), .ZN(n88445) );
  OAI21_X1 U74016 ( .B1(n88448), .B2(n105787), .A(n88449), .ZN(n88447) );
  OAI21_X1 U74017 ( .B1(n88450), .B2(n88451), .A(n105786), .ZN(n88449) );
  OAI21_X1 U74018 ( .B1(n108386), .B2(n86311), .A(n88452), .ZN(n88451) );
  AOI22_X1 U74019 ( .A1(n86313), .A2(n71019), .B1(n105784), .B2(n108384), .ZN(
        n88452) );
  NAND2_X1 U74020 ( .A1(n88453), .A2(n88454), .ZN(n88450) );
  AOI22_X1 U74021 ( .A1(n105783), .A2(n108382), .B1(n105782), .B2(n108387), 
        .ZN(n88454) );
  AOI22_X1 U74022 ( .A1(n105781), .A2(n108385), .B1(n105780), .B2(n108383), 
        .ZN(n88453) );
  NOR4_X1 U74023 ( .A1(n88455), .A2(n88456), .A3(n88457), .A4(n88458), .ZN(
        n88448) );
  NAND2_X1 U74024 ( .A1(n88459), .A2(n88460), .ZN(n88458) );
  NOR4_X1 U74025 ( .A1(n88461), .A2(n88462), .A3(n88463), .A4(n88464), .ZN(
        n88460) );
  NAND2_X1 U74026 ( .A1(n88465), .A2(n88466), .ZN(n88464) );
  AOI22_X1 U74027 ( .A1(n105779), .A2(n108363), .B1(n105778), .B2(n108364), 
        .ZN(n88466) );
  AOI22_X1 U74028 ( .A1(n105777), .A2(n108372), .B1(n105776), .B2(n108370), 
        .ZN(n88465) );
  NAND2_X1 U74029 ( .A1(n88467), .A2(n88468), .ZN(n88463) );
  AOI22_X1 U74030 ( .A1(n105775), .A2(n70888), .B1(n105774), .B2(n108367), 
        .ZN(n88468) );
  AOI22_X1 U74031 ( .A1(n105773), .A2(n70992), .B1(n105772), .B2(n108283), 
        .ZN(n88467) );
  NAND2_X1 U74032 ( .A1(n88469), .A2(n88470), .ZN(n88462) );
  AOI22_X1 U74033 ( .A1(n105771), .A2(n108287), .B1(n105770), .B2(n70892), 
        .ZN(n88470) );
  AOI22_X1 U74034 ( .A1(n105769), .A2(n108368), .B1(n105768), .B2(n108365), 
        .ZN(n88469) );
  NAND2_X1 U74035 ( .A1(n88471), .A2(n88472), .ZN(n88461) );
  AOI22_X1 U74036 ( .A1(n105767), .A2(n108285), .B1(n105766), .B2(n108289), 
        .ZN(n88472) );
  AOI22_X1 U74037 ( .A1(n105765), .A2(n108288), .B1(n105764), .B2(n70894), 
        .ZN(n88471) );
  NOR4_X1 U74038 ( .A1(n88473), .A2(n88474), .A3(n88475), .A4(n88476), .ZN(
        n88459) );
  NAND2_X1 U74039 ( .A1(n88477), .A2(n88478), .ZN(n88476) );
  AOI22_X1 U74040 ( .A1(n105763), .A2(n108373), .B1(n105762), .B2(n108376), 
        .ZN(n88478) );
  AOI22_X1 U74041 ( .A1(n105761), .A2(n108377), .B1(n105760), .B2(n108379), 
        .ZN(n88477) );
  NAND2_X1 U74042 ( .A1(n88479), .A2(n88480), .ZN(n88475) );
  AOI22_X1 U74043 ( .A1(n105759), .A2(n108378), .B1(n105758), .B2(n108374), 
        .ZN(n88480) );
  AOI22_X1 U74044 ( .A1(n105757), .A2(n108380), .B1(n105756), .B2(n108375), 
        .ZN(n88479) );
  NAND2_X1 U74045 ( .A1(n88481), .A2(n88482), .ZN(n88474) );
  AOI22_X1 U74046 ( .A1(n105755), .A2(n71002), .B1(n105754), .B2(n71001), .ZN(
        n88482) );
  AOI22_X1 U74047 ( .A1(n105753), .A2(n71004), .B1(n105752), .B2(n108381), 
        .ZN(n88481) );
  NAND2_X1 U74048 ( .A1(n88483), .A2(n88484), .ZN(n88473) );
  AOI22_X1 U74049 ( .A1(n105751), .A2(n108366), .B1(n105750), .B2(n108371), 
        .ZN(n88484) );
  AOI22_X1 U74050 ( .A1(n105749), .A2(n70999), .B1(n105748), .B2(n108369), 
        .ZN(n88483) );
  NAND2_X1 U74051 ( .A1(n88485), .A2(n88486), .ZN(n88457) );
  NOR4_X1 U74052 ( .A1(n88487), .A2(n88488), .A3(n88489), .A4(n88490), .ZN(
        n88486) );
  NAND2_X1 U74053 ( .A1(n88491), .A2(n88492), .ZN(n88490) );
  AOI22_X1 U74054 ( .A1(n105747), .A2(n108298), .B1(n105746), .B2(n108300), 
        .ZN(n88492) );
  AOI22_X1 U74055 ( .A1(n105745), .A2(n70917), .B1(n105744), .B2(n108299), 
        .ZN(n88491) );
  NAND2_X1 U74056 ( .A1(n88493), .A2(n88494), .ZN(n88489) );
  AOI22_X1 U74057 ( .A1(n105743), .A2(n70921), .B1(n105742), .B2(n70923), .ZN(
        n88494) );
  AOI22_X1 U74058 ( .A1(n105741), .A2(n108306), .B1(n105740), .B2(n108307), 
        .ZN(n88493) );
  NAND2_X1 U74059 ( .A1(n88495), .A2(n88496), .ZN(n88488) );
  AOI22_X1 U74060 ( .A1(n105739), .A2(n108303), .B1(n105738), .B2(n108305), 
        .ZN(n88496) );
  AOI22_X1 U74061 ( .A1(n105737), .A2(n108308), .B1(n105736), .B2(n108304), 
        .ZN(n88495) );
  NAND2_X1 U74062 ( .A1(n88497), .A2(n88498), .ZN(n88487) );
  AOI22_X1 U74063 ( .A1(n105735), .A2(n108313), .B1(n105734), .B2(n70928), 
        .ZN(n88498) );
  AOI22_X1 U74064 ( .A1(n105733), .A2(n108312), .B1(n105732), .B2(n70926), 
        .ZN(n88497) );
  NOR4_X1 U74065 ( .A1(n88499), .A2(n88500), .A3(n88501), .A4(n88502), .ZN(
        n88485) );
  NAND2_X1 U74066 ( .A1(n88503), .A2(n88504), .ZN(n88502) );
  AOI22_X1 U74067 ( .A1(n105731), .A2(n108293), .B1(n105730), .B2(n108284), 
        .ZN(n88504) );
  AOI22_X1 U74068 ( .A1(n105729), .A2(n108286), .B1(n105728), .B2(n70900), 
        .ZN(n88503) );
  NAND2_X1 U74069 ( .A1(n88505), .A2(n88506), .ZN(n88501) );
  AOI22_X1 U74070 ( .A1(n105727), .A2(n108291), .B1(n105726), .B2(n108295), 
        .ZN(n88506) );
  AOI22_X1 U74071 ( .A1(n105725), .A2(n108297), .B1(n105724), .B2(n108294), 
        .ZN(n88505) );
  NAND2_X1 U74072 ( .A1(n88507), .A2(n88508), .ZN(n88500) );
  AOI22_X1 U74073 ( .A1(n105723), .A2(n70909), .B1(n105722), .B2(n108290), 
        .ZN(n88508) );
  AOI22_X1 U74074 ( .A1(n105721), .A2(n108292), .B1(n105720), .B2(n108296), 
        .ZN(n88507) );
  NAND2_X1 U74075 ( .A1(n88509), .A2(n88510), .ZN(n88499) );
  AOI22_X1 U74076 ( .A1(n105719), .A2(n108302), .B1(n105718), .B2(n70913), 
        .ZN(n88510) );
  AOI22_X1 U74077 ( .A1(n105717), .A2(n70911), .B1(n105716), .B2(n108301), 
        .ZN(n88509) );
  NAND2_X1 U74078 ( .A1(n88511), .A2(n88512), .ZN(n88456) );
  NOR4_X1 U74079 ( .A1(n88513), .A2(n88514), .A3(n88515), .A4(n88516), .ZN(
        n88512) );
  NAND2_X1 U74080 ( .A1(n88517), .A2(n88518), .ZN(n88516) );
  AOI22_X1 U74081 ( .A1(n105715), .A2(n70951), .B1(n105714), .B2(n108323), 
        .ZN(n88518) );
  AOI22_X1 U74082 ( .A1(n105713), .A2(n108327), .B1(n105712), .B2(n108326), 
        .ZN(n88517) );
  NAND2_X1 U74083 ( .A1(n88519), .A2(n88520), .ZN(n88515) );
  AOI22_X1 U74084 ( .A1(n105711), .A2(n108332), .B1(n105710), .B2(n108331), 
        .ZN(n88520) );
  AOI22_X1 U74085 ( .A1(n105709), .A2(n108322), .B1(n86458), .B2(n108324), 
        .ZN(n88519) );
  NAND2_X1 U74086 ( .A1(n88521), .A2(n88522), .ZN(n88514) );
  AOI22_X1 U74087 ( .A1(n105707), .A2(n108333), .B1(n105706), .B2(n108329), 
        .ZN(n88522) );
  AOI22_X1 U74088 ( .A1(n105705), .A2(n70955), .B1(n105704), .B2(n70957), .ZN(
        n88521) );
  NAND2_X1 U74089 ( .A1(n88523), .A2(n88524), .ZN(n88513) );
  AOI22_X1 U74090 ( .A1(n105703), .A2(n108336), .B1(n105702), .B2(n70963), 
        .ZN(n88524) );
  AOI22_X1 U74091 ( .A1(n105701), .A2(n108328), .B1(n105700), .B2(n108330), 
        .ZN(n88523) );
  NOR4_X1 U74092 ( .A1(n88525), .A2(n88526), .A3(n88527), .A4(n88528), .ZN(
        n88511) );
  NAND2_X1 U74093 ( .A1(n88529), .A2(n88530), .ZN(n88528) );
  AOI22_X1 U74094 ( .A1(n105699), .A2(n108311), .B1(n105698), .B2(n108316), 
        .ZN(n88530) );
  AOI22_X1 U74095 ( .A1(n105697), .A2(n108310), .B1(n105696), .B2(n70931), 
        .ZN(n88529) );
  NAND2_X1 U74096 ( .A1(n88531), .A2(n88532), .ZN(n88527) );
  AOI22_X1 U74097 ( .A1(n105695), .A2(n70940), .B1(n105694), .B2(n108318), 
        .ZN(n88532) );
  AOI22_X1 U74098 ( .A1(n105693), .A2(n108319), .B1(n105692), .B2(n108309), 
        .ZN(n88531) );
  NAND2_X1 U74099 ( .A1(n88533), .A2(n88534), .ZN(n88526) );
  AOI22_X1 U74100 ( .A1(n105691), .A2(n108317), .B1(n105690), .B2(n108321), 
        .ZN(n88534) );
  AOI22_X1 U74101 ( .A1(n105689), .A2(n108315), .B1(n105688), .B2(n108320), 
        .ZN(n88533) );
  NAND2_X1 U74102 ( .A1(n88535), .A2(n88536), .ZN(n88525) );
  AOI22_X1 U74103 ( .A1(n105687), .A2(n70945), .B1(n105686), .B2(n108325), 
        .ZN(n88536) );
  AOI22_X1 U74104 ( .A1(n105685), .A2(n70943), .B1(n105684), .B2(n108314), 
        .ZN(n88535) );
  NAND2_X1 U74105 ( .A1(n88537), .A2(n88538), .ZN(n88455) );
  NOR4_X1 U74106 ( .A1(n88539), .A2(n88540), .A3(n88541), .A4(n88542), .ZN(
        n88538) );
  NAND2_X1 U74107 ( .A1(n88543), .A2(n88544), .ZN(n88542) );
  AOI22_X1 U74108 ( .A1(n105683), .A2(n108354), .B1(n105682), .B2(n108353), 
        .ZN(n88544) );
  AOI22_X1 U74109 ( .A1(n105681), .A2(n70979), .B1(n105680), .B2(n108351), 
        .ZN(n88543) );
  NAND2_X1 U74110 ( .A1(n88545), .A2(n88546), .ZN(n88541) );
  AOI22_X1 U74111 ( .A1(n105679), .A2(n108349), .B1(n105678), .B2(n108352), 
        .ZN(n88546) );
  AOI22_X1 U74112 ( .A1(n86515), .A2(n70985), .B1(n105677), .B2(n108350), .ZN(
        n88545) );
  NAND2_X1 U74113 ( .A1(n88547), .A2(n88548), .ZN(n88540) );
  AOI22_X1 U74114 ( .A1(n86519), .A2(n108360), .B1(n86520), .B2(n70991), .ZN(
        n88548) );
  AOI22_X1 U74115 ( .A1(n86521), .A2(n108358), .B1(n86522), .B2(n108359), .ZN(
        n88547) );
  NAND2_X1 U74116 ( .A1(n88549), .A2(n88550), .ZN(n88539) );
  AOI22_X1 U74117 ( .A1(n105676), .A2(n108355), .B1(n86526), .B2(n108357), 
        .ZN(n88550) );
  AOI22_X1 U74118 ( .A1(n86527), .A2(n108361), .B1(n86528), .B2(n108356), .ZN(
        n88549) );
  NOR4_X1 U74119 ( .A1(n88551), .A2(n88552), .A3(n88553), .A4(n88554), .ZN(
        n88537) );
  NAND2_X1 U74120 ( .A1(n88555), .A2(n88556), .ZN(n88554) );
  AOI22_X1 U74121 ( .A1(n105675), .A2(n108335), .B1(n105674), .B2(n108339), 
        .ZN(n88556) );
  AOI22_X1 U74122 ( .A1(n105673), .A2(n108338), .B1(n105672), .B2(n70962), 
        .ZN(n88555) );
  NAND2_X1 U74123 ( .A1(n88557), .A2(n88558), .ZN(n88553) );
  AOI22_X1 U74124 ( .A1(n105671), .A2(n108345), .B1(n105670), .B2(n108334), 
        .ZN(n88558) );
  AOI22_X1 U74125 ( .A1(n105669), .A2(n108337), .B1(n105668), .B2(n108342), 
        .ZN(n88557) );
  NAND2_X1 U74126 ( .A1(n88559), .A2(n88560), .ZN(n88552) );
  AOI22_X1 U74127 ( .A1(n105667), .A2(n108341), .B1(n105666), .B2(n108346), 
        .ZN(n88560) );
  AOI22_X1 U74128 ( .A1(n105665), .A2(n108348), .B1(n86550), .B2(n108344), 
        .ZN(n88559) );
  NAND2_X1 U74129 ( .A1(n88561), .A2(n88562), .ZN(n88551) );
  AOI22_X1 U74130 ( .A1(n105663), .A2(n70980), .B1(n105662), .B2(n108340), 
        .ZN(n88562) );
  AOI22_X1 U74131 ( .A1(n105661), .A2(n108343), .B1(n105660), .B2(n108347), 
        .ZN(n88561) );
  AOI21_X1 U74132 ( .B1(n86302), .B2(n88564), .A(n88565), .ZN(n88563) );
  OAI21_X1 U74133 ( .B1(n88566), .B2(n105787), .A(n88567), .ZN(n88565) );
  OAI21_X1 U74134 ( .B1(n88568), .B2(n88569), .A(n105786), .ZN(n88567) );
  OAI21_X1 U74135 ( .B1(n108497), .B2(n105785), .A(n88570), .ZN(n88569) );
  AOI22_X1 U74136 ( .A1(n86313), .A2(n71164), .B1(n105784), .B2(n108495), .ZN(
        n88570) );
  NAND2_X1 U74137 ( .A1(n88571), .A2(n88572), .ZN(n88568) );
  AOI22_X1 U74138 ( .A1(n105783), .A2(n108493), .B1(n105782), .B2(n108498), 
        .ZN(n88572) );
  AOI22_X1 U74139 ( .A1(n105781), .A2(n108496), .B1(n105780), .B2(n108494), 
        .ZN(n88571) );
  NOR4_X1 U74140 ( .A1(n88573), .A2(n88574), .A3(n88575), .A4(n88576), .ZN(
        n88566) );
  NAND2_X1 U74141 ( .A1(n88577), .A2(n88578), .ZN(n88576) );
  NOR4_X1 U74142 ( .A1(n88579), .A2(n88580), .A3(n88581), .A4(n88582), .ZN(
        n88578) );
  NAND2_X1 U74143 ( .A1(n88583), .A2(n88584), .ZN(n88582) );
  AOI22_X1 U74144 ( .A1(n105779), .A2(n108474), .B1(n105778), .B2(n108475), 
        .ZN(n88584) );
  AOI22_X1 U74145 ( .A1(n105777), .A2(n108483), .B1(n105776), .B2(n108481), 
        .ZN(n88583) );
  NAND2_X1 U74146 ( .A1(n88585), .A2(n88586), .ZN(n88581) );
  AOI22_X1 U74147 ( .A1(n105775), .A2(n71033), .B1(n105774), .B2(n108478), 
        .ZN(n88586) );
  AOI22_X1 U74148 ( .A1(n105773), .A2(n71137), .B1(n105772), .B2(n108394), 
        .ZN(n88585) );
  NAND2_X1 U74149 ( .A1(n88587), .A2(n88588), .ZN(n88580) );
  AOI22_X1 U74150 ( .A1(n105771), .A2(n108398), .B1(n86346), .B2(n71037), .ZN(
        n88588) );
  AOI22_X1 U74151 ( .A1(n105769), .A2(n108479), .B1(n105768), .B2(n108476), 
        .ZN(n88587) );
  NAND2_X1 U74152 ( .A1(n88589), .A2(n88590), .ZN(n88579) );
  AOI22_X1 U74153 ( .A1(n105767), .A2(n108396), .B1(n105766), .B2(n108400), 
        .ZN(n88590) );
  AOI22_X1 U74154 ( .A1(n105765), .A2(n108399), .B1(n105764), .B2(n71039), 
        .ZN(n88589) );
  NOR4_X1 U74155 ( .A1(n88591), .A2(n88592), .A3(n88593), .A4(n88594), .ZN(
        n88577) );
  NAND2_X1 U74156 ( .A1(n88595), .A2(n88596), .ZN(n88594) );
  AOI22_X1 U74157 ( .A1(n105763), .A2(n108484), .B1(n105762), .B2(n108487), 
        .ZN(n88596) );
  AOI22_X1 U74158 ( .A1(n86363), .A2(n108488), .B1(n105760), .B2(n108490), 
        .ZN(n88595) );
  NAND2_X1 U74159 ( .A1(n88597), .A2(n88598), .ZN(n88593) );
  AOI22_X1 U74160 ( .A1(n105759), .A2(n108489), .B1(n86368), .B2(n108485), 
        .ZN(n88598) );
  AOI22_X1 U74161 ( .A1(n105757), .A2(n108491), .B1(n105756), .B2(n108486), 
        .ZN(n88597) );
  NAND2_X1 U74162 ( .A1(n88599), .A2(n88600), .ZN(n88592) );
  AOI22_X1 U74163 ( .A1(n105755), .A2(n71147), .B1(n105754), .B2(n71146), .ZN(
        n88600) );
  AOI22_X1 U74164 ( .A1(n105753), .A2(n71149), .B1(n105752), .B2(n108492), 
        .ZN(n88599) );
  NAND2_X1 U74165 ( .A1(n88601), .A2(n88602), .ZN(n88591) );
  AOI22_X1 U74166 ( .A1(n105751), .A2(n108477), .B1(n105750), .B2(n108482), 
        .ZN(n88602) );
  AOI22_X1 U74167 ( .A1(n105749), .A2(n71144), .B1(n105748), .B2(n108480), 
        .ZN(n88601) );
  NAND2_X1 U74168 ( .A1(n88603), .A2(n88604), .ZN(n88575) );
  NOR4_X1 U74169 ( .A1(n88605), .A2(n88606), .A3(n88607), .A4(n88608), .ZN(
        n88604) );
  NAND2_X1 U74170 ( .A1(n88609), .A2(n88610), .ZN(n88608) );
  AOI22_X1 U74171 ( .A1(n105747), .A2(n108409), .B1(n105746), .B2(n108411), 
        .ZN(n88610) );
  AOI22_X1 U74172 ( .A1(n105745), .A2(n71062), .B1(n105744), .B2(n108410), 
        .ZN(n88609) );
  NAND2_X1 U74173 ( .A1(n88611), .A2(n88612), .ZN(n88607) );
  AOI22_X1 U74174 ( .A1(n105743), .A2(n71066), .B1(n105742), .B2(n71068), .ZN(
        n88612) );
  AOI22_X1 U74175 ( .A1(n105741), .A2(n108417), .B1(n86400), .B2(n108418), 
        .ZN(n88611) );
  NAND2_X1 U74176 ( .A1(n88613), .A2(n88614), .ZN(n88606) );
  AOI22_X1 U74177 ( .A1(n86403), .A2(n108414), .B1(n105738), .B2(n108416), 
        .ZN(n88614) );
  AOI22_X1 U74178 ( .A1(n105737), .A2(n108419), .B1(n105736), .B2(n108415), 
        .ZN(n88613) );
  NAND2_X1 U74179 ( .A1(n88615), .A2(n88616), .ZN(n88605) );
  AOI22_X1 U74180 ( .A1(n105735), .A2(n108424), .B1(n105734), .B2(n71073), 
        .ZN(n88616) );
  AOI22_X1 U74181 ( .A1(n86411), .A2(n108423), .B1(n105732), .B2(n71071), .ZN(
        n88615) );
  NOR4_X1 U74182 ( .A1(n88617), .A2(n88618), .A3(n88619), .A4(n88620), .ZN(
        n88603) );
  NAND2_X1 U74183 ( .A1(n88621), .A2(n88622), .ZN(n88620) );
  AOI22_X1 U74184 ( .A1(n105731), .A2(n108404), .B1(n105730), .B2(n108395), 
        .ZN(n88622) );
  AOI22_X1 U74185 ( .A1(n105729), .A2(n108397), .B1(n105728), .B2(n71045), 
        .ZN(n88621) );
  NAND2_X1 U74186 ( .A1(n88623), .A2(n88624), .ZN(n88619) );
  AOI22_X1 U74187 ( .A1(n105727), .A2(n108402), .B1(n86426), .B2(n108406), 
        .ZN(n88624) );
  AOI22_X1 U74188 ( .A1(n105725), .A2(n108408), .B1(n86428), .B2(n108405), 
        .ZN(n88623) );
  NAND2_X1 U74189 ( .A1(n88625), .A2(n88626), .ZN(n88618) );
  AOI22_X1 U74190 ( .A1(n105723), .A2(n71054), .B1(n105722), .B2(n108401), 
        .ZN(n88626) );
  AOI22_X1 U74191 ( .A1(n105721), .A2(n108403), .B1(n105720), .B2(n108407), 
        .ZN(n88625) );
  NAND2_X1 U74192 ( .A1(n88627), .A2(n88628), .ZN(n88617) );
  AOI22_X1 U74193 ( .A1(n105719), .A2(n108413), .B1(n105718), .B2(n71058), 
        .ZN(n88628) );
  AOI22_X1 U74194 ( .A1(n105717), .A2(n71056), .B1(n105716), .B2(n108412), 
        .ZN(n88627) );
  NAND2_X1 U74195 ( .A1(n88629), .A2(n88630), .ZN(n88574) );
  NOR4_X1 U74196 ( .A1(n88631), .A2(n88632), .A3(n88633), .A4(n88634), .ZN(
        n88630) );
  NAND2_X1 U74197 ( .A1(n88635), .A2(n88636), .ZN(n88634) );
  AOI22_X1 U74198 ( .A1(n105715), .A2(n71096), .B1(n86450), .B2(n108434), .ZN(
        n88636) );
  AOI22_X1 U74199 ( .A1(n105713), .A2(n108438), .B1(n105712), .B2(n108437), 
        .ZN(n88635) );
  NAND2_X1 U74200 ( .A1(n88637), .A2(n88638), .ZN(n88633) );
  AOI22_X1 U74201 ( .A1(n105711), .A2(n108443), .B1(n105710), .B2(n108442), 
        .ZN(n88638) );
  AOI22_X1 U74202 ( .A1(n105709), .A2(n108433), .B1(n86458), .B2(n108435), 
        .ZN(n88637) );
  NAND2_X1 U74203 ( .A1(n88639), .A2(n88640), .ZN(n88632) );
  AOI22_X1 U74204 ( .A1(n105707), .A2(n108444), .B1(n105706), .B2(n108440), 
        .ZN(n88640) );
  AOI22_X1 U74205 ( .A1(n105705), .A2(n71100), .B1(n105704), .B2(n71102), .ZN(
        n88639) );
  NAND2_X1 U74206 ( .A1(n88641), .A2(n88642), .ZN(n88631) );
  AOI22_X1 U74207 ( .A1(n86467), .A2(n108447), .B1(n105702), .B2(n71108), .ZN(
        n88642) );
  AOI22_X1 U74208 ( .A1(n105701), .A2(n108439), .B1(n105700), .B2(n108441), 
        .ZN(n88641) );
  NOR4_X1 U74209 ( .A1(n88643), .A2(n88644), .A3(n88645), .A4(n88646), .ZN(
        n88629) );
  NAND2_X1 U74210 ( .A1(n88647), .A2(n88648), .ZN(n88646) );
  AOI22_X1 U74211 ( .A1(n105699), .A2(n108422), .B1(n105698), .B2(n108427), 
        .ZN(n88648) );
  AOI22_X1 U74212 ( .A1(n105697), .A2(n108421), .B1(n105696), .B2(n71076), 
        .ZN(n88647) );
  NAND2_X1 U74213 ( .A1(n88649), .A2(n88650), .ZN(n88645) );
  AOI22_X1 U74214 ( .A1(n105695), .A2(n71085), .B1(n86484), .B2(n108429), .ZN(
        n88650) );
  AOI22_X1 U74215 ( .A1(n105693), .A2(n108430), .B1(n105692), .B2(n108420), 
        .ZN(n88649) );
  NAND2_X1 U74216 ( .A1(n88651), .A2(n88652), .ZN(n88644) );
  AOI22_X1 U74217 ( .A1(n105691), .A2(n108428), .B1(n86490), .B2(n108432), 
        .ZN(n88652) );
  AOI22_X1 U74218 ( .A1(n105689), .A2(n108426), .B1(n105688), .B2(n108431), 
        .ZN(n88651) );
  NAND2_X1 U74219 ( .A1(n88653), .A2(n88654), .ZN(n88643) );
  AOI22_X1 U74220 ( .A1(n105687), .A2(n71090), .B1(n105686), .B2(n108436), 
        .ZN(n88654) );
  AOI22_X1 U74221 ( .A1(n105685), .A2(n71088), .B1(n105684), .B2(n108425), 
        .ZN(n88653) );
  NAND2_X1 U74222 ( .A1(n88655), .A2(n88656), .ZN(n88573) );
  NOR4_X1 U74223 ( .A1(n88657), .A2(n88658), .A3(n88659), .A4(n88660), .ZN(
        n88656) );
  NAND2_X1 U74224 ( .A1(n88661), .A2(n88662), .ZN(n88660) );
  AOI22_X1 U74225 ( .A1(n105683), .A2(n108465), .B1(n105682), .B2(n108464), 
        .ZN(n88662) );
  AOI22_X1 U74226 ( .A1(n105681), .A2(n71124), .B1(n105680), .B2(n108462), 
        .ZN(n88661) );
  NAND2_X1 U74227 ( .A1(n88663), .A2(n88664), .ZN(n88659) );
  AOI22_X1 U74228 ( .A1(n105679), .A2(n108460), .B1(n105678), .B2(n108463), 
        .ZN(n88664) );
  AOI22_X1 U74229 ( .A1(n86515), .A2(n71130), .B1(n86516), .B2(n108461), .ZN(
        n88663) );
  NAND2_X1 U74230 ( .A1(n88665), .A2(n88666), .ZN(n88658) );
  AOI22_X1 U74231 ( .A1(n86519), .A2(n108471), .B1(n86520), .B2(n71136), .ZN(
        n88666) );
  AOI22_X1 U74232 ( .A1(n86521), .A2(n108469), .B1(n86522), .B2(n108470), .ZN(
        n88665) );
  NAND2_X1 U74233 ( .A1(n88667), .A2(n88668), .ZN(n88657) );
  AOI22_X1 U74234 ( .A1(n105676), .A2(n108466), .B1(n86526), .B2(n108468), 
        .ZN(n88668) );
  AOI22_X1 U74235 ( .A1(n86527), .A2(n108472), .B1(n86528), .B2(n108467), .ZN(
        n88667) );
  NOR4_X1 U74236 ( .A1(n88669), .A2(n88670), .A3(n88671), .A4(n88672), .ZN(
        n88655) );
  NAND2_X1 U74237 ( .A1(n88673), .A2(n88674), .ZN(n88672) );
  AOI22_X1 U74238 ( .A1(n105675), .A2(n108446), .B1(n105674), .B2(n108450), 
        .ZN(n88674) );
  AOI22_X1 U74239 ( .A1(n105673), .A2(n108449), .B1(n105672), .B2(n71107), 
        .ZN(n88673) );
  NAND2_X1 U74240 ( .A1(n88675), .A2(n88676), .ZN(n88671) );
  AOI22_X1 U74241 ( .A1(n105671), .A2(n108456), .B1(n105670), .B2(n108445), 
        .ZN(n88676) );
  AOI22_X1 U74242 ( .A1(n105669), .A2(n108448), .B1(n105668), .B2(n108453), 
        .ZN(n88675) );
  NAND2_X1 U74243 ( .A1(n88677), .A2(n88678), .ZN(n88670) );
  AOI22_X1 U74244 ( .A1(n105667), .A2(n108452), .B1(n105666), .B2(n108457), 
        .ZN(n88678) );
  AOI22_X1 U74245 ( .A1(n86549), .A2(n108459), .B1(n105664), .B2(n108455), 
        .ZN(n88677) );
  NAND2_X1 U74246 ( .A1(n88679), .A2(n88680), .ZN(n88669) );
  AOI22_X1 U74247 ( .A1(n105663), .A2(n71125), .B1(n105662), .B2(n108451), 
        .ZN(n88680) );
  AOI22_X1 U74248 ( .A1(n86555), .A2(n108454), .B1(n105660), .B2(n108458), 
        .ZN(n88679) );
  AOI21_X1 U74249 ( .B1(n86302), .B2(n88682), .A(n88683), .ZN(n88681) );
  OAI21_X1 U74250 ( .B1(n88684), .B2(n105787), .A(n88685), .ZN(n88683) );
  OAI21_X1 U74251 ( .B1(n88686), .B2(n88687), .A(n105786), .ZN(n88685) );
  OAI21_X1 U74252 ( .B1(n107734), .B2(n86311), .A(n88688), .ZN(n88687) );
  AOI22_X1 U74253 ( .A1(n86313), .A2(n70125), .B1(n105784), .B2(n107732), .ZN(
        n88688) );
  NAND2_X1 U74254 ( .A1(n88689), .A2(n88690), .ZN(n88686) );
  AOI22_X1 U74255 ( .A1(n105783), .A2(n107730), .B1(n105782), .B2(n107735), 
        .ZN(n88690) );
  AOI22_X1 U74256 ( .A1(n105781), .A2(n107733), .B1(n105780), .B2(n107731), 
        .ZN(n88689) );
  NOR4_X1 U74257 ( .A1(n88691), .A2(n88692), .A3(n88693), .A4(n88694), .ZN(
        n88684) );
  NAND2_X1 U74258 ( .A1(n88695), .A2(n88696), .ZN(n88694) );
  NOR4_X1 U74259 ( .A1(n88697), .A2(n88698), .A3(n88699), .A4(n88700), .ZN(
        n88696) );
  NAND2_X1 U74260 ( .A1(n88701), .A2(n88702), .ZN(n88700) );
  AOI22_X1 U74261 ( .A1(n105779), .A2(n107711), .B1(n105778), .B2(n107712), 
        .ZN(n88702) );
  AOI22_X1 U74262 ( .A1(n105777), .A2(n107720), .B1(n105776), .B2(n107718), 
        .ZN(n88701) );
  NAND2_X1 U74263 ( .A1(n88703), .A2(n88704), .ZN(n88699) );
  AOI22_X1 U74264 ( .A1(n105775), .A2(n69994), .B1(n105774), .B2(n107715), 
        .ZN(n88704) );
  AOI22_X1 U74265 ( .A1(n105773), .A2(n70098), .B1(n105772), .B2(n107632), 
        .ZN(n88703) );
  NAND2_X1 U74266 ( .A1(n88705), .A2(n88706), .ZN(n88698) );
  AOI22_X1 U74267 ( .A1(n105771), .A2(n107636), .B1(n105770), .B2(n69998), 
        .ZN(n88706) );
  AOI22_X1 U74268 ( .A1(n105769), .A2(n107716), .B1(n105768), .B2(n107713), 
        .ZN(n88705) );
  NAND2_X1 U74269 ( .A1(n88707), .A2(n88708), .ZN(n88697) );
  AOI22_X1 U74270 ( .A1(n105767), .A2(n107634), .B1(n105766), .B2(n107638), 
        .ZN(n88708) );
  AOI22_X1 U74271 ( .A1(n105765), .A2(n107637), .B1(n105764), .B2(n70000), 
        .ZN(n88707) );
  NOR4_X1 U74272 ( .A1(n88709), .A2(n88710), .A3(n88711), .A4(n88712), .ZN(
        n88695) );
  NAND2_X1 U74273 ( .A1(n88713), .A2(n88714), .ZN(n88712) );
  AOI22_X1 U74274 ( .A1(n105763), .A2(n107721), .B1(n105762), .B2(n107724), 
        .ZN(n88714) );
  AOI22_X1 U74275 ( .A1(n105761), .A2(n107725), .B1(n105760), .B2(n107727), 
        .ZN(n88713) );
  NAND2_X1 U74276 ( .A1(n88715), .A2(n88716), .ZN(n88711) );
  AOI22_X1 U74277 ( .A1(n105759), .A2(n107726), .B1(n105758), .B2(n107722), 
        .ZN(n88716) );
  AOI22_X1 U74278 ( .A1(n105757), .A2(n107728), .B1(n105756), .B2(n107723), 
        .ZN(n88715) );
  NAND2_X1 U74279 ( .A1(n88717), .A2(n88718), .ZN(n88710) );
  AOI22_X1 U74280 ( .A1(n105755), .A2(n70108), .B1(n105754), .B2(n70107), .ZN(
        n88718) );
  AOI22_X1 U74281 ( .A1(n105753), .A2(n70110), .B1(n105752), .B2(n107729), 
        .ZN(n88717) );
  NAND2_X1 U74282 ( .A1(n88719), .A2(n88720), .ZN(n88709) );
  AOI22_X1 U74283 ( .A1(n105751), .A2(n107714), .B1(n105750), .B2(n107719), 
        .ZN(n88720) );
  AOI22_X1 U74284 ( .A1(n105749), .A2(n70105), .B1(n105748), .B2(n107717), 
        .ZN(n88719) );
  NAND2_X1 U74285 ( .A1(n88721), .A2(n88722), .ZN(n88693) );
  NOR4_X1 U74286 ( .A1(n88723), .A2(n88724), .A3(n88725), .A4(n88726), .ZN(
        n88722) );
  NAND2_X1 U74287 ( .A1(n88727), .A2(n88728), .ZN(n88726) );
  AOI22_X1 U74288 ( .A1(n105747), .A2(n107647), .B1(n105746), .B2(n107649), 
        .ZN(n88728) );
  AOI22_X1 U74289 ( .A1(n105745), .A2(n70023), .B1(n105744), .B2(n107648), 
        .ZN(n88727) );
  NAND2_X1 U74290 ( .A1(n88729), .A2(n88730), .ZN(n88725) );
  AOI22_X1 U74291 ( .A1(n105743), .A2(n70027), .B1(n105742), .B2(n70029), .ZN(
        n88730) );
  AOI22_X1 U74292 ( .A1(n105741), .A2(n107655), .B1(n105740), .B2(n107656), 
        .ZN(n88729) );
  NAND2_X1 U74293 ( .A1(n88731), .A2(n88732), .ZN(n88724) );
  AOI22_X1 U74294 ( .A1(n105739), .A2(n107652), .B1(n105738), .B2(n107654), 
        .ZN(n88732) );
  AOI22_X1 U74295 ( .A1(n105737), .A2(n107657), .B1(n105736), .B2(n107653), 
        .ZN(n88731) );
  NAND2_X1 U74296 ( .A1(n88733), .A2(n88734), .ZN(n88723) );
  AOI22_X1 U74297 ( .A1(n105735), .A2(n107662), .B1(n105734), .B2(n70034), 
        .ZN(n88734) );
  AOI22_X1 U74298 ( .A1(n105733), .A2(n107661), .B1(n105732), .B2(n70032), 
        .ZN(n88733) );
  NOR4_X1 U74299 ( .A1(n88735), .A2(n88736), .A3(n88737), .A4(n88738), .ZN(
        n88721) );
  NAND2_X1 U74300 ( .A1(n88739), .A2(n88740), .ZN(n88738) );
  AOI22_X1 U74301 ( .A1(n105731), .A2(n107642), .B1(n105730), .B2(n107633), 
        .ZN(n88740) );
  AOI22_X1 U74302 ( .A1(n105729), .A2(n107635), .B1(n105728), .B2(n70006), 
        .ZN(n88739) );
  NAND2_X1 U74303 ( .A1(n88741), .A2(n88742), .ZN(n88737) );
  AOI22_X1 U74304 ( .A1(n105727), .A2(n107640), .B1(n105726), .B2(n107644), 
        .ZN(n88742) );
  AOI22_X1 U74305 ( .A1(n105725), .A2(n107646), .B1(n105724), .B2(n107643), 
        .ZN(n88741) );
  NAND2_X1 U74306 ( .A1(n88743), .A2(n88744), .ZN(n88736) );
  AOI22_X1 U74307 ( .A1(n105723), .A2(n70015), .B1(n105722), .B2(n107639), 
        .ZN(n88744) );
  AOI22_X1 U74308 ( .A1(n105721), .A2(n107641), .B1(n105720), .B2(n107645), 
        .ZN(n88743) );
  NAND2_X1 U74309 ( .A1(n88745), .A2(n88746), .ZN(n88735) );
  AOI22_X1 U74310 ( .A1(n105719), .A2(n107651), .B1(n105718), .B2(n70019), 
        .ZN(n88746) );
  AOI22_X1 U74311 ( .A1(n105717), .A2(n70017), .B1(n105716), .B2(n107650), 
        .ZN(n88745) );
  NAND2_X1 U74312 ( .A1(n88747), .A2(n88748), .ZN(n88692) );
  NOR4_X1 U74313 ( .A1(n88749), .A2(n88750), .A3(n88751), .A4(n88752), .ZN(
        n88748) );
  NAND2_X1 U74314 ( .A1(n88753), .A2(n88754), .ZN(n88752) );
  AOI22_X1 U74315 ( .A1(n105715), .A2(n70057), .B1(n105714), .B2(n107672), 
        .ZN(n88754) );
  AOI22_X1 U74316 ( .A1(n105713), .A2(n107676), .B1(n105712), .B2(n107675), 
        .ZN(n88753) );
  NAND2_X1 U74317 ( .A1(n88755), .A2(n88756), .ZN(n88751) );
  AOI22_X1 U74318 ( .A1(n105711), .A2(n107681), .B1(n105710), .B2(n107680), 
        .ZN(n88756) );
  AOI22_X1 U74319 ( .A1(n105709), .A2(n107671), .B1(n86458), .B2(n107673), 
        .ZN(n88755) );
  NAND2_X1 U74320 ( .A1(n88757), .A2(n88758), .ZN(n88750) );
  AOI22_X1 U74321 ( .A1(n105707), .A2(n107682), .B1(n105706), .B2(n107678), 
        .ZN(n88758) );
  AOI22_X1 U74322 ( .A1(n105705), .A2(n70061), .B1(n105704), .B2(n70063), .ZN(
        n88757) );
  NAND2_X1 U74323 ( .A1(n88759), .A2(n88760), .ZN(n88749) );
  AOI22_X1 U74324 ( .A1(n105703), .A2(n107685), .B1(n105702), .B2(n70069), 
        .ZN(n88760) );
  AOI22_X1 U74325 ( .A1(n105701), .A2(n107677), .B1(n105700), .B2(n107679), 
        .ZN(n88759) );
  NOR4_X1 U74326 ( .A1(n88761), .A2(n88762), .A3(n88763), .A4(n88764), .ZN(
        n88747) );
  NAND2_X1 U74327 ( .A1(n88765), .A2(n88766), .ZN(n88764) );
  AOI22_X1 U74328 ( .A1(n105699), .A2(n107660), .B1(n105698), .B2(n107665), 
        .ZN(n88766) );
  AOI22_X1 U74329 ( .A1(n105697), .A2(n107659), .B1(n105696), .B2(n70037), 
        .ZN(n88765) );
  NAND2_X1 U74330 ( .A1(n88767), .A2(n88768), .ZN(n88763) );
  AOI22_X1 U74331 ( .A1(n105695), .A2(n70046), .B1(n86484), .B2(n107667), .ZN(
        n88768) );
  AOI22_X1 U74332 ( .A1(n105693), .A2(n107668), .B1(n105692), .B2(n107658), 
        .ZN(n88767) );
  NAND2_X1 U74333 ( .A1(n88769), .A2(n88770), .ZN(n88762) );
  AOI22_X1 U74334 ( .A1(n105691), .A2(n107666), .B1(n105690), .B2(n107670), 
        .ZN(n88770) );
  AOI22_X1 U74335 ( .A1(n105689), .A2(n107664), .B1(n105688), .B2(n107669), 
        .ZN(n88769) );
  NAND2_X1 U74336 ( .A1(n88771), .A2(n88772), .ZN(n88761) );
  AOI22_X1 U74337 ( .A1(n105687), .A2(n70051), .B1(n105686), .B2(n107674), 
        .ZN(n88772) );
  AOI22_X1 U74338 ( .A1(n105685), .A2(n70049), .B1(n105684), .B2(n107663), 
        .ZN(n88771) );
  NAND2_X1 U74339 ( .A1(n88773), .A2(n88774), .ZN(n88691) );
  NOR4_X1 U74340 ( .A1(n88775), .A2(n88776), .A3(n88777), .A4(n88778), .ZN(
        n88774) );
  NAND2_X1 U74341 ( .A1(n88779), .A2(n88780), .ZN(n88778) );
  AOI22_X1 U74342 ( .A1(n105683), .A2(n107703), .B1(n105682), .B2(n107702), 
        .ZN(n88780) );
  AOI22_X1 U74343 ( .A1(n105681), .A2(n70085), .B1(n105680), .B2(n107700), 
        .ZN(n88779) );
  NAND2_X1 U74344 ( .A1(n88781), .A2(n88782), .ZN(n88777) );
  AOI22_X1 U74345 ( .A1(n105679), .A2(n107698), .B1(n105678), .B2(n107701), 
        .ZN(n88782) );
  AOI22_X1 U74346 ( .A1(n86515), .A2(n70091), .B1(n105677), .B2(n107699), .ZN(
        n88781) );
  NAND2_X1 U74347 ( .A1(n88783), .A2(n88784), .ZN(n88776) );
  AOI22_X1 U74348 ( .A1(n86519), .A2(n107709), .B1(n86520), .B2(n70097), .ZN(
        n88784) );
  AOI22_X1 U74349 ( .A1(n86521), .A2(n107707), .B1(n86522), .B2(n107708), .ZN(
        n88783) );
  NAND2_X1 U74350 ( .A1(n88785), .A2(n88786), .ZN(n88775) );
  AOI22_X1 U74351 ( .A1(n105676), .A2(n107704), .B1(n86526), .B2(n107706), 
        .ZN(n88786) );
  AOI22_X1 U74352 ( .A1(n86527), .A2(n107710), .B1(n86528), .B2(n107705), .ZN(
        n88785) );
  NOR4_X1 U74353 ( .A1(n88787), .A2(n88788), .A3(n88789), .A4(n88790), .ZN(
        n88773) );
  NAND2_X1 U74354 ( .A1(n88791), .A2(n88792), .ZN(n88790) );
  AOI22_X1 U74355 ( .A1(n105675), .A2(n107684), .B1(n105674), .B2(n107688), 
        .ZN(n88792) );
  AOI22_X1 U74356 ( .A1(n105673), .A2(n107687), .B1(n105672), .B2(n70068), 
        .ZN(n88791) );
  NAND2_X1 U74357 ( .A1(n88793), .A2(n88794), .ZN(n88789) );
  AOI22_X1 U74358 ( .A1(n105671), .A2(n107694), .B1(n105670), .B2(n107683), 
        .ZN(n88794) );
  AOI22_X1 U74359 ( .A1(n105669), .A2(n107686), .B1(n105668), .B2(n107691), 
        .ZN(n88793) );
  NAND2_X1 U74360 ( .A1(n88795), .A2(n88796), .ZN(n88788) );
  AOI22_X1 U74361 ( .A1(n105667), .A2(n107690), .B1(n105666), .B2(n107695), 
        .ZN(n88796) );
  AOI22_X1 U74362 ( .A1(n105665), .A2(n107697), .B1(n86550), .B2(n107693), 
        .ZN(n88795) );
  NAND2_X1 U74363 ( .A1(n88797), .A2(n88798), .ZN(n88787) );
  AOI22_X1 U74364 ( .A1(n105663), .A2(n70086), .B1(n105662), .B2(n107689), 
        .ZN(n88798) );
  AOI22_X1 U74365 ( .A1(n86555), .A2(n107692), .B1(n105660), .B2(n107696), 
        .ZN(n88797) );
  AOI21_X1 U74366 ( .B1(n86302), .B2(n88800), .A(n88801), .ZN(n88799) );
  OAI21_X1 U74367 ( .B1(n88802), .B2(n105787), .A(n88803), .ZN(n88801) );
  OAI21_X1 U74368 ( .B1(n88804), .B2(n88805), .A(n105786), .ZN(n88803) );
  OAI21_X1 U74369 ( .B1(n109649), .B2(n105785), .A(n88806), .ZN(n88805) );
  AOI22_X1 U74370 ( .A1(n86313), .A2(n72654), .B1(n86314), .B2(n109647), .ZN(
        n88806) );
  NAND2_X1 U74371 ( .A1(n88807), .A2(n88808), .ZN(n88804) );
  AOI22_X1 U74372 ( .A1(n105783), .A2(n109645), .B1(n105782), .B2(n109650), 
        .ZN(n88808) );
  AOI22_X1 U74373 ( .A1(n105781), .A2(n109648), .B1(n105780), .B2(n109646), 
        .ZN(n88807) );
  NOR4_X1 U74374 ( .A1(n88809), .A2(n88810), .A3(n88811), .A4(n88812), .ZN(
        n88802) );
  NAND2_X1 U74375 ( .A1(n88813), .A2(n88814), .ZN(n88812) );
  NOR4_X1 U74376 ( .A1(n88815), .A2(n88816), .A3(n88817), .A4(n88818), .ZN(
        n88814) );
  NAND2_X1 U74377 ( .A1(n88819), .A2(n88820), .ZN(n88818) );
  AOI22_X1 U74378 ( .A1(n105779), .A2(n109626), .B1(n105778), .B2(n109627), 
        .ZN(n88820) );
  AOI22_X1 U74379 ( .A1(n105777), .A2(n109635), .B1(n105776), .B2(n109633), 
        .ZN(n88819) );
  NAND2_X1 U74380 ( .A1(n88821), .A2(n88822), .ZN(n88817) );
  AOI22_X1 U74381 ( .A1(n105775), .A2(n72523), .B1(n105774), .B2(n109630), 
        .ZN(n88822) );
  AOI22_X1 U74382 ( .A1(n105773), .A2(n72627), .B1(n105772), .B2(n109550), 
        .ZN(n88821) );
  NAND2_X1 U74383 ( .A1(n88823), .A2(n88824), .ZN(n88816) );
  AOI22_X1 U74384 ( .A1(n105771), .A2(n109554), .B1(n86346), .B2(n72527), .ZN(
        n88824) );
  AOI22_X1 U74385 ( .A1(n105769), .A2(n109631), .B1(n105768), .B2(n109628), 
        .ZN(n88823) );
  NAND2_X1 U74386 ( .A1(n88825), .A2(n88826), .ZN(n88815) );
  AOI22_X1 U74387 ( .A1(n105767), .A2(n109552), .B1(n105766), .B2(n109556), 
        .ZN(n88826) );
  AOI22_X1 U74388 ( .A1(n105765), .A2(n109555), .B1(n105764), .B2(n72529), 
        .ZN(n88825) );
  NOR4_X1 U74389 ( .A1(n88827), .A2(n88828), .A3(n88829), .A4(n88830), .ZN(
        n88813) );
  NAND2_X1 U74390 ( .A1(n88831), .A2(n88832), .ZN(n88830) );
  AOI22_X1 U74391 ( .A1(n105763), .A2(n109636), .B1(n105762), .B2(n109639), 
        .ZN(n88832) );
  AOI22_X1 U74392 ( .A1(n105761), .A2(n109640), .B1(n86364), .B2(n109642), 
        .ZN(n88831) );
  NAND2_X1 U74393 ( .A1(n88833), .A2(n88834), .ZN(n88829) );
  AOI22_X1 U74394 ( .A1(n105759), .A2(n109641), .B1(n86368), .B2(n109637), 
        .ZN(n88834) );
  AOI22_X1 U74395 ( .A1(n105757), .A2(n109643), .B1(n105756), .B2(n109638), 
        .ZN(n88833) );
  NAND2_X1 U74396 ( .A1(n88835), .A2(n88836), .ZN(n88828) );
  AOI22_X1 U74397 ( .A1(n105755), .A2(n72637), .B1(n105754), .B2(n72636), .ZN(
        n88836) );
  AOI22_X1 U74398 ( .A1(n105753), .A2(n72639), .B1(n105752), .B2(n109644), 
        .ZN(n88835) );
  NAND2_X1 U74399 ( .A1(n88837), .A2(n88838), .ZN(n88827) );
  AOI22_X1 U74400 ( .A1(n105751), .A2(n109629), .B1(n105750), .B2(n109634), 
        .ZN(n88838) );
  AOI22_X1 U74401 ( .A1(n105749), .A2(n72634), .B1(n86382), .B2(n109632), .ZN(
        n88837) );
  NAND2_X1 U74402 ( .A1(n88839), .A2(n88840), .ZN(n88811) );
  NOR4_X1 U74403 ( .A1(n88841), .A2(n88842), .A3(n88843), .A4(n88844), .ZN(
        n88840) );
  NAND2_X1 U74404 ( .A1(n88845), .A2(n88846), .ZN(n88844) );
  AOI22_X1 U74405 ( .A1(n105747), .A2(n109565), .B1(n105746), .B2(n109567), 
        .ZN(n88846) );
  AOI22_X1 U74406 ( .A1(n105745), .A2(n72552), .B1(n105744), .B2(n109566), 
        .ZN(n88845) );
  NAND2_X1 U74407 ( .A1(n88847), .A2(n88848), .ZN(n88843) );
  AOI22_X1 U74408 ( .A1(n105743), .A2(n72556), .B1(n105742), .B2(n72558), .ZN(
        n88848) );
  AOI22_X1 U74409 ( .A1(n105741), .A2(n109573), .B1(n86400), .B2(n109574), 
        .ZN(n88847) );
  NAND2_X1 U74410 ( .A1(n88849), .A2(n88850), .ZN(n88842) );
  AOI22_X1 U74411 ( .A1(n86403), .A2(n109570), .B1(n105738), .B2(n109572), 
        .ZN(n88850) );
  AOI22_X1 U74412 ( .A1(n105737), .A2(n109575), .B1(n86406), .B2(n109571), 
        .ZN(n88849) );
  NAND2_X1 U74413 ( .A1(n88851), .A2(n88852), .ZN(n88841) );
  AOI22_X1 U74414 ( .A1(n105735), .A2(n109580), .B1(n105734), .B2(n72563), 
        .ZN(n88852) );
  AOI22_X1 U74415 ( .A1(n86411), .A2(n109579), .B1(n105732), .B2(n72561), .ZN(
        n88851) );
  NOR4_X1 U74416 ( .A1(n88853), .A2(n88854), .A3(n88855), .A4(n88856), .ZN(
        n88839) );
  NAND2_X1 U74417 ( .A1(n88857), .A2(n88858), .ZN(n88856) );
  AOI22_X1 U74418 ( .A1(n105731), .A2(n109560), .B1(n105730), .B2(n109551), 
        .ZN(n88858) );
  AOI22_X1 U74419 ( .A1(n105729), .A2(n109553), .B1(n105728), .B2(n72535), 
        .ZN(n88857) );
  NAND2_X1 U74420 ( .A1(n88859), .A2(n88860), .ZN(n88855) );
  AOI22_X1 U74421 ( .A1(n105727), .A2(n109558), .B1(n86426), .B2(n109562), 
        .ZN(n88860) );
  AOI22_X1 U74422 ( .A1(n86427), .A2(n109564), .B1(n86428), .B2(n109561), .ZN(
        n88859) );
  NAND2_X1 U74423 ( .A1(n88861), .A2(n88862), .ZN(n88854) );
  AOI22_X1 U74424 ( .A1(n105723), .A2(n72544), .B1(n105722), .B2(n109557), 
        .ZN(n88862) );
  AOI22_X1 U74425 ( .A1(n105721), .A2(n109559), .B1(n105720), .B2(n109563), 
        .ZN(n88861) );
  NAND2_X1 U74426 ( .A1(n88863), .A2(n88864), .ZN(n88853) );
  AOI22_X1 U74427 ( .A1(n105719), .A2(n109569), .B1(n105718), .B2(n72548), 
        .ZN(n88864) );
  AOI22_X1 U74428 ( .A1(n105717), .A2(n72546), .B1(n86440), .B2(n109568), .ZN(
        n88863) );
  NAND2_X1 U74429 ( .A1(n88865), .A2(n88866), .ZN(n88810) );
  NOR4_X1 U74430 ( .A1(n88867), .A2(n88868), .A3(n88869), .A4(n88870), .ZN(
        n88866) );
  NAND2_X1 U74431 ( .A1(n88871), .A2(n88872), .ZN(n88870) );
  AOI22_X1 U74432 ( .A1(n105715), .A2(n72586), .B1(n86450), .B2(n109590), .ZN(
        n88872) );
  AOI22_X1 U74433 ( .A1(n105713), .A2(n109594), .B1(n105712), .B2(n109593), 
        .ZN(n88871) );
  NAND2_X1 U74434 ( .A1(n88873), .A2(n88874), .ZN(n88869) );
  AOI22_X1 U74435 ( .A1(n86455), .A2(n109599), .B1(n105710), .B2(n109598), 
        .ZN(n88874) );
  AOI22_X1 U74436 ( .A1(n86457), .A2(n109589), .B1(n105708), .B2(n109591), 
        .ZN(n88873) );
  NAND2_X1 U74437 ( .A1(n88875), .A2(n88876), .ZN(n88868) );
  AOI22_X1 U74438 ( .A1(n105707), .A2(n109600), .B1(n105706), .B2(n109596), 
        .ZN(n88876) );
  AOI22_X1 U74439 ( .A1(n105705), .A2(n72590), .B1(n105704), .B2(n72592), .ZN(
        n88875) );
  NAND2_X1 U74440 ( .A1(n88877), .A2(n88878), .ZN(n88867) );
  AOI22_X1 U74441 ( .A1(n86467), .A2(n109603), .B1(n105702), .B2(n72598), .ZN(
        n88878) );
  AOI22_X1 U74442 ( .A1(n105701), .A2(n109595), .B1(n105700), .B2(n109597), 
        .ZN(n88877) );
  NOR4_X1 U74443 ( .A1(n88879), .A2(n88880), .A3(n88881), .A4(n88882), .ZN(
        n88865) );
  NAND2_X1 U74444 ( .A1(n88883), .A2(n88884), .ZN(n88882) );
  AOI22_X1 U74445 ( .A1(n105699), .A2(n109578), .B1(n105698), .B2(n109583), 
        .ZN(n88884) );
  AOI22_X1 U74446 ( .A1(n86479), .A2(n109577), .B1(n105696), .B2(n72566), .ZN(
        n88883) );
  NAND2_X1 U74447 ( .A1(n88885), .A2(n88886), .ZN(n88881) );
  AOI22_X1 U74448 ( .A1(n105695), .A2(n72575), .B1(n86484), .B2(n109585), .ZN(
        n88886) );
  AOI22_X1 U74449 ( .A1(n105693), .A2(n109586), .B1(n105692), .B2(n109576), 
        .ZN(n88885) );
  NAND2_X1 U74450 ( .A1(n88887), .A2(n88888), .ZN(n88880) );
  AOI22_X1 U74451 ( .A1(n105691), .A2(n109584), .B1(n86490), .B2(n109588), 
        .ZN(n88888) );
  AOI22_X1 U74452 ( .A1(n105689), .A2(n109582), .B1(n105688), .B2(n109587), 
        .ZN(n88887) );
  NAND2_X1 U74453 ( .A1(n88889), .A2(n88890), .ZN(n88879) );
  AOI22_X1 U74454 ( .A1(n86495), .A2(n72580), .B1(n105686), .B2(n109592), .ZN(
        n88890) );
  AOI22_X1 U74455 ( .A1(n105685), .A2(n72578), .B1(n105684), .B2(n109581), 
        .ZN(n88889) );
  NAND2_X1 U74456 ( .A1(n88891), .A2(n88892), .ZN(n88809) );
  NOR4_X1 U74457 ( .A1(n88893), .A2(n88894), .A3(n88895), .A4(n88896), .ZN(
        n88892) );
  NAND2_X1 U74458 ( .A1(n88897), .A2(n88898), .ZN(n88896) );
  AOI22_X1 U74459 ( .A1(n105683), .A2(n109618), .B1(n105682), .B2(n109617), 
        .ZN(n88898) );
  AOI22_X1 U74460 ( .A1(n105681), .A2(n72614), .B1(n105680), .B2(n109615), 
        .ZN(n88897) );
  NAND2_X1 U74461 ( .A1(n88899), .A2(n88900), .ZN(n88895) );
  AOI22_X1 U74462 ( .A1(n105679), .A2(n109613), .B1(n86514), .B2(n109616), 
        .ZN(n88900) );
  AOI22_X1 U74463 ( .A1(n86515), .A2(n72620), .B1(n86516), .B2(n109614), .ZN(
        n88899) );
  NAND2_X1 U74464 ( .A1(n88901), .A2(n88902), .ZN(n88894) );
  AOI22_X1 U74465 ( .A1(n86519), .A2(n109624), .B1(n86520), .B2(n72626), .ZN(
        n88902) );
  AOI22_X1 U74466 ( .A1(n86521), .A2(n109622), .B1(n86522), .B2(n109623), .ZN(
        n88901) );
  NAND2_X1 U74467 ( .A1(n88903), .A2(n88904), .ZN(n88893) );
  AOI22_X1 U74468 ( .A1(n105676), .A2(n109619), .B1(n86526), .B2(n109621), 
        .ZN(n88904) );
  AOI22_X1 U74469 ( .A1(n86527), .A2(n109625), .B1(n86528), .B2(n109620), .ZN(
        n88903) );
  NOR4_X1 U74470 ( .A1(n88905), .A2(n88906), .A3(n88907), .A4(n88908), .ZN(
        n88891) );
  NAND2_X1 U74471 ( .A1(n88909), .A2(n88910), .ZN(n88908) );
  AOI22_X1 U74472 ( .A1(n86535), .A2(n109602), .B1(n105674), .B2(n72600), .ZN(
        n88910) );
  AOI22_X1 U74473 ( .A1(n105673), .A2(n109605), .B1(n105672), .B2(n72597), 
        .ZN(n88909) );
  NAND2_X1 U74474 ( .A1(n88911), .A2(n88912), .ZN(n88907) );
  AOI22_X1 U74475 ( .A1(n105671), .A2(n109610), .B1(n105670), .B2(n109601), 
        .ZN(n88912) );
  AOI22_X1 U74476 ( .A1(n105669), .A2(n109604), .B1(n86544), .B2(n72603), .ZN(
        n88911) );
  NAND2_X1 U74477 ( .A1(n88913), .A2(n88914), .ZN(n88906) );
  AOI22_X1 U74478 ( .A1(n105667), .A2(n109607), .B1(n105666), .B2(n72607), 
        .ZN(n88914) );
  AOI22_X1 U74479 ( .A1(n86549), .A2(n109612), .B1(n105664), .B2(n109609), 
        .ZN(n88913) );
  NAND2_X1 U74480 ( .A1(n88915), .A2(n88916), .ZN(n88905) );
  AOI22_X1 U74481 ( .A1(n105663), .A2(n72615), .B1(n105662), .B2(n109606), 
        .ZN(n88916) );
  AOI22_X1 U74482 ( .A1(n105661), .A2(n109608), .B1(n86556), .B2(n109611), 
        .ZN(n88915) );
  AOI21_X1 U74483 ( .B1(n86302), .B2(n88918), .A(n88919), .ZN(n88917) );
  OAI21_X1 U74484 ( .B1(n88920), .B2(n105787), .A(n88921), .ZN(n88919) );
  OAI21_X1 U74485 ( .B1(n88922), .B2(n88923), .A(n105786), .ZN(n88921) );
  OAI21_X1 U74486 ( .B1(n108611), .B2(n105785), .A(n88924), .ZN(n88923) );
  AOI22_X1 U74487 ( .A1(n86313), .A2(n71313), .B1(n86314), .B2(n108609), .ZN(
        n88924) );
  NAND2_X1 U74488 ( .A1(n88925), .A2(n88926), .ZN(n88922) );
  AOI22_X1 U74489 ( .A1(n105783), .A2(n108607), .B1(n105782), .B2(n108612), 
        .ZN(n88926) );
  AOI22_X1 U74490 ( .A1(n105781), .A2(n108610), .B1(n105780), .B2(n108608), 
        .ZN(n88925) );
  NOR4_X1 U74491 ( .A1(n88927), .A2(n88928), .A3(n88929), .A4(n88930), .ZN(
        n88920) );
  NAND2_X1 U74492 ( .A1(n88931), .A2(n88932), .ZN(n88930) );
  NOR4_X1 U74493 ( .A1(n88933), .A2(n88934), .A3(n88935), .A4(n88936), .ZN(
        n88932) );
  NAND2_X1 U74494 ( .A1(n88937), .A2(n88938), .ZN(n88936) );
  AOI22_X1 U74495 ( .A1(n105779), .A2(n108588), .B1(n105778), .B2(n108589), 
        .ZN(n88938) );
  AOI22_X1 U74496 ( .A1(n105777), .A2(n108597), .B1(n105776), .B2(n108595), 
        .ZN(n88937) );
  NAND2_X1 U74497 ( .A1(n88939), .A2(n88940), .ZN(n88935) );
  AOI22_X1 U74498 ( .A1(n105775), .A2(n71182), .B1(n105774), .B2(n108592), 
        .ZN(n88940) );
  AOI22_X1 U74499 ( .A1(n105773), .A2(n71286), .B1(n105772), .B2(n108511), 
        .ZN(n88939) );
  NAND2_X1 U74500 ( .A1(n88941), .A2(n88942), .ZN(n88934) );
  AOI22_X1 U74501 ( .A1(n105771), .A2(n108515), .B1(n86346), .B2(n71186), .ZN(
        n88942) );
  AOI22_X1 U74502 ( .A1(n105769), .A2(n108593), .B1(n105768), .B2(n108590), 
        .ZN(n88941) );
  NAND2_X1 U74503 ( .A1(n88943), .A2(n88944), .ZN(n88933) );
  AOI22_X1 U74504 ( .A1(n105767), .A2(n108513), .B1(n105766), .B2(n108517), 
        .ZN(n88944) );
  AOI22_X1 U74505 ( .A1(n105765), .A2(n108516), .B1(n105764), .B2(n71188), 
        .ZN(n88943) );
  NOR4_X1 U74506 ( .A1(n88945), .A2(n88946), .A3(n88947), .A4(n88948), .ZN(
        n88931) );
  NAND2_X1 U74507 ( .A1(n88949), .A2(n88950), .ZN(n88948) );
  AOI22_X1 U74508 ( .A1(n105763), .A2(n108598), .B1(n105762), .B2(n108601), 
        .ZN(n88950) );
  AOI22_X1 U74509 ( .A1(n105761), .A2(n108602), .B1(n86364), .B2(n108604), 
        .ZN(n88949) );
  NAND2_X1 U74510 ( .A1(n88951), .A2(n88952), .ZN(n88947) );
  AOI22_X1 U74511 ( .A1(n105759), .A2(n108603), .B1(n86368), .B2(n108599), 
        .ZN(n88952) );
  AOI22_X1 U74512 ( .A1(n105757), .A2(n108605), .B1(n105756), .B2(n108600), 
        .ZN(n88951) );
  NAND2_X1 U74513 ( .A1(n88953), .A2(n88954), .ZN(n88946) );
  AOI22_X1 U74514 ( .A1(n105755), .A2(n71296), .B1(n105754), .B2(n71295), .ZN(
        n88954) );
  AOI22_X1 U74515 ( .A1(n105753), .A2(n71298), .B1(n105752), .B2(n108606), 
        .ZN(n88953) );
  NAND2_X1 U74516 ( .A1(n88955), .A2(n88956), .ZN(n88945) );
  AOI22_X1 U74517 ( .A1(n105751), .A2(n108591), .B1(n105750), .B2(n108596), 
        .ZN(n88956) );
  AOI22_X1 U74518 ( .A1(n105749), .A2(n71293), .B1(n86382), .B2(n108594), .ZN(
        n88955) );
  NAND2_X1 U74519 ( .A1(n88957), .A2(n88958), .ZN(n88929) );
  NOR4_X1 U74520 ( .A1(n88959), .A2(n88960), .A3(n88961), .A4(n88962), .ZN(
        n88958) );
  NAND2_X1 U74521 ( .A1(n88963), .A2(n88964), .ZN(n88962) );
  AOI22_X1 U74522 ( .A1(n105747), .A2(n108526), .B1(n105746), .B2(n108528), 
        .ZN(n88964) );
  AOI22_X1 U74523 ( .A1(n105745), .A2(n71211), .B1(n105744), .B2(n108527), 
        .ZN(n88963) );
  NAND2_X1 U74524 ( .A1(n88965), .A2(n88966), .ZN(n88961) );
  AOI22_X1 U74525 ( .A1(n105743), .A2(n71215), .B1(n105742), .B2(n71217), .ZN(
        n88966) );
  AOI22_X1 U74526 ( .A1(n105741), .A2(n108534), .B1(n86400), .B2(n108535), 
        .ZN(n88965) );
  NAND2_X1 U74527 ( .A1(n88967), .A2(n88968), .ZN(n88960) );
  AOI22_X1 U74528 ( .A1(n86403), .A2(n108531), .B1(n105738), .B2(n108533), 
        .ZN(n88968) );
  AOI22_X1 U74529 ( .A1(n105737), .A2(n108536), .B1(n86406), .B2(n108532), 
        .ZN(n88967) );
  NAND2_X1 U74530 ( .A1(n88969), .A2(n88970), .ZN(n88959) );
  AOI22_X1 U74531 ( .A1(n105735), .A2(n108541), .B1(n105734), .B2(n71222), 
        .ZN(n88970) );
  AOI22_X1 U74532 ( .A1(n86411), .A2(n108540), .B1(n105732), .B2(n71220), .ZN(
        n88969) );
  NOR4_X1 U74533 ( .A1(n88971), .A2(n88972), .A3(n88973), .A4(n88974), .ZN(
        n88957) );
  NAND2_X1 U74534 ( .A1(n88975), .A2(n88976), .ZN(n88974) );
  AOI22_X1 U74535 ( .A1(n105731), .A2(n108521), .B1(n105730), .B2(n108512), 
        .ZN(n88976) );
  AOI22_X1 U74536 ( .A1(n105729), .A2(n108514), .B1(n105728), .B2(n71194), 
        .ZN(n88975) );
  NAND2_X1 U74537 ( .A1(n88977), .A2(n88978), .ZN(n88973) );
  AOI22_X1 U74538 ( .A1(n105727), .A2(n108519), .B1(n86426), .B2(n108523), 
        .ZN(n88978) );
  AOI22_X1 U74539 ( .A1(n86427), .A2(n108525), .B1(n86428), .B2(n108522), .ZN(
        n88977) );
  NAND2_X1 U74540 ( .A1(n88979), .A2(n88980), .ZN(n88972) );
  AOI22_X1 U74541 ( .A1(n105723), .A2(n71203), .B1(n105722), .B2(n108518), 
        .ZN(n88980) );
  AOI22_X1 U74542 ( .A1(n105721), .A2(n108520), .B1(n105720), .B2(n108524), 
        .ZN(n88979) );
  NAND2_X1 U74543 ( .A1(n88981), .A2(n88982), .ZN(n88971) );
  AOI22_X1 U74544 ( .A1(n105719), .A2(n108530), .B1(n105718), .B2(n71207), 
        .ZN(n88982) );
  AOI22_X1 U74545 ( .A1(n105717), .A2(n71205), .B1(n86440), .B2(n108529), .ZN(
        n88981) );
  NAND2_X1 U74546 ( .A1(n88983), .A2(n88984), .ZN(n88928) );
  NOR4_X1 U74547 ( .A1(n88985), .A2(n88986), .A3(n88987), .A4(n88988), .ZN(
        n88984) );
  NAND2_X1 U74548 ( .A1(n88989), .A2(n88990), .ZN(n88988) );
  AOI22_X1 U74549 ( .A1(n105715), .A2(n71245), .B1(n86450), .B2(n108551), .ZN(
        n88990) );
  AOI22_X1 U74550 ( .A1(n105713), .A2(n108555), .B1(n105712), .B2(n108554), 
        .ZN(n88989) );
  NAND2_X1 U74551 ( .A1(n88991), .A2(n88992), .ZN(n88987) );
  AOI22_X1 U74552 ( .A1(n86455), .A2(n108560), .B1(n105710), .B2(n108559), 
        .ZN(n88992) );
  AOI22_X1 U74553 ( .A1(n86457), .A2(n108550), .B1(n105708), .B2(n108552), 
        .ZN(n88991) );
  NAND2_X1 U74554 ( .A1(n88993), .A2(n88994), .ZN(n88986) );
  AOI22_X1 U74555 ( .A1(n105707), .A2(n108561), .B1(n105706), .B2(n108557), 
        .ZN(n88994) );
  AOI22_X1 U74556 ( .A1(n105705), .A2(n71249), .B1(n105704), .B2(n71251), .ZN(
        n88993) );
  NAND2_X1 U74557 ( .A1(n88995), .A2(n88996), .ZN(n88985) );
  AOI22_X1 U74558 ( .A1(n86467), .A2(n108564), .B1(n105702), .B2(n71257), .ZN(
        n88996) );
  AOI22_X1 U74559 ( .A1(n105701), .A2(n108556), .B1(n105700), .B2(n108558), 
        .ZN(n88995) );
  NOR4_X1 U74560 ( .A1(n88997), .A2(n88998), .A3(n88999), .A4(n89000), .ZN(
        n88983) );
  NAND2_X1 U74561 ( .A1(n89001), .A2(n89002), .ZN(n89000) );
  AOI22_X1 U74562 ( .A1(n105699), .A2(n108539), .B1(n105698), .B2(n108544), 
        .ZN(n89002) );
  AOI22_X1 U74563 ( .A1(n86479), .A2(n108538), .B1(n105696), .B2(n71225), .ZN(
        n89001) );
  NAND2_X1 U74564 ( .A1(n89003), .A2(n89004), .ZN(n88999) );
  AOI22_X1 U74565 ( .A1(n105695), .A2(n71234), .B1(n86484), .B2(n108546), .ZN(
        n89004) );
  AOI22_X1 U74566 ( .A1(n105693), .A2(n108547), .B1(n105692), .B2(n108537), 
        .ZN(n89003) );
  NAND2_X1 U74567 ( .A1(n89005), .A2(n89006), .ZN(n88998) );
  AOI22_X1 U74568 ( .A1(n105691), .A2(n108545), .B1(n86490), .B2(n108549), 
        .ZN(n89006) );
  AOI22_X1 U74569 ( .A1(n105689), .A2(n108543), .B1(n105688), .B2(n108548), 
        .ZN(n89005) );
  NAND2_X1 U74570 ( .A1(n89007), .A2(n89008), .ZN(n88997) );
  AOI22_X1 U74571 ( .A1(n86495), .A2(n71239), .B1(n105686), .B2(n108553), .ZN(
        n89008) );
  AOI22_X1 U74572 ( .A1(n105685), .A2(n71237), .B1(n105684), .B2(n108542), 
        .ZN(n89007) );
  NAND2_X1 U74573 ( .A1(n89009), .A2(n89010), .ZN(n88927) );
  NOR4_X1 U74574 ( .A1(n89011), .A2(n89012), .A3(n89013), .A4(n89014), .ZN(
        n89010) );
  NAND2_X1 U74575 ( .A1(n89015), .A2(n89016), .ZN(n89014) );
  AOI22_X1 U74576 ( .A1(n105683), .A2(n108580), .B1(n105682), .B2(n108579), 
        .ZN(n89016) );
  AOI22_X1 U74577 ( .A1(n105681), .A2(n71273), .B1(n105680), .B2(n108577), 
        .ZN(n89015) );
  NAND2_X1 U74578 ( .A1(n89017), .A2(n89018), .ZN(n89013) );
  AOI22_X1 U74579 ( .A1(n105679), .A2(n108575), .B1(n86514), .B2(n108578), 
        .ZN(n89018) );
  AOI22_X1 U74580 ( .A1(n86515), .A2(n71279), .B1(n86516), .B2(n108576), .ZN(
        n89017) );
  NAND2_X1 U74581 ( .A1(n89019), .A2(n89020), .ZN(n89012) );
  AOI22_X1 U74582 ( .A1(n86519), .A2(n108586), .B1(n86520), .B2(n71285), .ZN(
        n89020) );
  AOI22_X1 U74583 ( .A1(n86521), .A2(n108584), .B1(n86522), .B2(n108585), .ZN(
        n89019) );
  NAND2_X1 U74584 ( .A1(n89021), .A2(n89022), .ZN(n89011) );
  AOI22_X1 U74585 ( .A1(n105676), .A2(n108581), .B1(n86526), .B2(n108583), 
        .ZN(n89022) );
  AOI22_X1 U74586 ( .A1(n86527), .A2(n108587), .B1(n86528), .B2(n108582), .ZN(
        n89021) );
  NOR4_X1 U74587 ( .A1(n89023), .A2(n89024), .A3(n89025), .A4(n89026), .ZN(
        n89009) );
  NAND2_X1 U74588 ( .A1(n89027), .A2(n89028), .ZN(n89026) );
  AOI22_X1 U74589 ( .A1(n86535), .A2(n108563), .B1(n105674), .B2(n108567), 
        .ZN(n89028) );
  AOI22_X1 U74590 ( .A1(n105673), .A2(n108566), .B1(n105672), .B2(n71256), 
        .ZN(n89027) );
  NAND2_X1 U74591 ( .A1(n89029), .A2(n89030), .ZN(n89025) );
  AOI22_X1 U74592 ( .A1(n105671), .A2(n108572), .B1(n105670), .B2(n108562), 
        .ZN(n89030) );
  AOI22_X1 U74593 ( .A1(n105669), .A2(n108565), .B1(n86544), .B2(n71262), .ZN(
        n89029) );
  NAND2_X1 U74594 ( .A1(n89031), .A2(n89032), .ZN(n89024) );
  AOI22_X1 U74595 ( .A1(n105667), .A2(n108569), .B1(n105666), .B2(n71266), 
        .ZN(n89032) );
  AOI22_X1 U74596 ( .A1(n86549), .A2(n108574), .B1(n105664), .B2(n108571), 
        .ZN(n89031) );
  NAND2_X1 U74597 ( .A1(n89033), .A2(n89034), .ZN(n89023) );
  AOI22_X1 U74598 ( .A1(n105663), .A2(n71274), .B1(n105662), .B2(n108568), 
        .ZN(n89034) );
  AOI22_X1 U74599 ( .A1(n86555), .A2(n108570), .B1(n86556), .B2(n108573), .ZN(
        n89033) );
  AOI21_X1 U74600 ( .B1(n86302), .B2(n81794), .A(n89036), .ZN(n89035) );
  OAI21_X1 U74601 ( .B1(n89037), .B2(n105787), .A(n89038), .ZN(n89036) );
  OAI21_X1 U74602 ( .B1(n89039), .B2(n89040), .A(n105786), .ZN(n89038) );
  OAI21_X1 U74603 ( .B1(n109756), .B2(n105785), .A(n89041), .ZN(n89040) );
  AOI22_X1 U74604 ( .A1(n86313), .A2(n72796), .B1(n86314), .B2(n109754), .ZN(
        n89041) );
  NAND2_X1 U74605 ( .A1(n89042), .A2(n89043), .ZN(n89039) );
  AOI22_X1 U74606 ( .A1(n105783), .A2(n109752), .B1(n105782), .B2(n109757), 
        .ZN(n89043) );
  AOI22_X1 U74607 ( .A1(n105781), .A2(n109755), .B1(n105780), .B2(n109753), 
        .ZN(n89042) );
  NOR4_X1 U74608 ( .A1(n89044), .A2(n89045), .A3(n89046), .A4(n89047), .ZN(
        n89037) );
  NAND2_X1 U74609 ( .A1(n89048), .A2(n89049), .ZN(n89047) );
  NOR4_X1 U74610 ( .A1(n89050), .A2(n89051), .A3(n89052), .A4(n89053), .ZN(
        n89049) );
  NAND2_X1 U74611 ( .A1(n89054), .A2(n89055), .ZN(n89053) );
  AOI22_X1 U74612 ( .A1(n105779), .A2(n109733), .B1(n105778), .B2(n109734), 
        .ZN(n89055) );
  AOI22_X1 U74613 ( .A1(n105777), .A2(n109742), .B1(n105776), .B2(n109740), 
        .ZN(n89054) );
  NAND2_X1 U74614 ( .A1(n89056), .A2(n89057), .ZN(n89052) );
  AOI22_X1 U74615 ( .A1(n105775), .A2(n72665), .B1(n105774), .B2(n109737), 
        .ZN(n89057) );
  AOI22_X1 U74616 ( .A1(n105773), .A2(n72769), .B1(n105772), .B2(n109655), 
        .ZN(n89056) );
  NAND2_X1 U74617 ( .A1(n89058), .A2(n89059), .ZN(n89051) );
  AOI22_X1 U74618 ( .A1(n105771), .A2(n109659), .B1(n105770), .B2(n72669), 
        .ZN(n89059) );
  AOI22_X1 U74619 ( .A1(n105769), .A2(n109738), .B1(n105768), .B2(n109735), 
        .ZN(n89058) );
  NAND2_X1 U74620 ( .A1(n89060), .A2(n89061), .ZN(n89050) );
  AOI22_X1 U74621 ( .A1(n105767), .A2(n109657), .B1(n105766), .B2(n109661), 
        .ZN(n89061) );
  AOI22_X1 U74622 ( .A1(n105765), .A2(n109660), .B1(n105764), .B2(n72671), 
        .ZN(n89060) );
  NOR4_X1 U74623 ( .A1(n89062), .A2(n89063), .A3(n89064), .A4(n89065), .ZN(
        n89048) );
  NAND2_X1 U74624 ( .A1(n89066), .A2(n89067), .ZN(n89065) );
  AOI22_X1 U74625 ( .A1(n105763), .A2(n109743), .B1(n105762), .B2(n109746), 
        .ZN(n89067) );
  AOI22_X1 U74626 ( .A1(n105761), .A2(n109747), .B1(n86364), .B2(n109749), 
        .ZN(n89066) );
  NAND2_X1 U74627 ( .A1(n89068), .A2(n89069), .ZN(n89064) );
  AOI22_X1 U74628 ( .A1(n105759), .A2(n109748), .B1(n105758), .B2(n109744), 
        .ZN(n89069) );
  AOI22_X1 U74629 ( .A1(n105757), .A2(n109750), .B1(n105756), .B2(n109745), 
        .ZN(n89068) );
  NAND2_X1 U74630 ( .A1(n89070), .A2(n89071), .ZN(n89063) );
  AOI22_X1 U74631 ( .A1(n105755), .A2(n72779), .B1(n105754), .B2(n72778), .ZN(
        n89071) );
  AOI22_X1 U74632 ( .A1(n105753), .A2(n72781), .B1(n105752), .B2(n109751), 
        .ZN(n89070) );
  NAND2_X1 U74633 ( .A1(n89072), .A2(n89073), .ZN(n89062) );
  AOI22_X1 U74634 ( .A1(n105751), .A2(n109736), .B1(n105750), .B2(n109741), 
        .ZN(n89073) );
  AOI22_X1 U74635 ( .A1(n105749), .A2(n72776), .B1(n86382), .B2(n109739), .ZN(
        n89072) );
  NAND2_X1 U74636 ( .A1(n89074), .A2(n89075), .ZN(n89046) );
  NOR4_X1 U74637 ( .A1(n89076), .A2(n89077), .A3(n89078), .A4(n89079), .ZN(
        n89075) );
  NAND2_X1 U74638 ( .A1(n89080), .A2(n89081), .ZN(n89079) );
  AOI22_X1 U74639 ( .A1(n105747), .A2(n109670), .B1(n105746), .B2(n109672), 
        .ZN(n89081) );
  AOI22_X1 U74640 ( .A1(n105745), .A2(n72694), .B1(n105744), .B2(n109671), 
        .ZN(n89080) );
  NAND2_X1 U74641 ( .A1(n89082), .A2(n89083), .ZN(n89078) );
  AOI22_X1 U74642 ( .A1(n105743), .A2(n72698), .B1(n105742), .B2(n72700), .ZN(
        n89083) );
  AOI22_X1 U74643 ( .A1(n105741), .A2(n109678), .B1(n105740), .B2(n109679), 
        .ZN(n89082) );
  NAND2_X1 U74644 ( .A1(n89084), .A2(n89085), .ZN(n89077) );
  AOI22_X1 U74645 ( .A1(n105739), .A2(n109675), .B1(n105738), .B2(n109677), 
        .ZN(n89085) );
  AOI22_X1 U74646 ( .A1(n105737), .A2(n109680), .B1(n86406), .B2(n109676), 
        .ZN(n89084) );
  NAND2_X1 U74647 ( .A1(n89086), .A2(n89087), .ZN(n89076) );
  AOI22_X1 U74648 ( .A1(n105735), .A2(n109685), .B1(n105734), .B2(n72705), 
        .ZN(n89087) );
  AOI22_X1 U74649 ( .A1(n105733), .A2(n109684), .B1(n105732), .B2(n72703), 
        .ZN(n89086) );
  NOR4_X1 U74650 ( .A1(n89088), .A2(n89089), .A3(n89090), .A4(n89091), .ZN(
        n89074) );
  NAND2_X1 U74651 ( .A1(n89092), .A2(n89093), .ZN(n89091) );
  AOI22_X1 U74652 ( .A1(n105731), .A2(n109665), .B1(n105730), .B2(n109656), 
        .ZN(n89093) );
  AOI22_X1 U74653 ( .A1(n105729), .A2(n109658), .B1(n105728), .B2(n72677), 
        .ZN(n89092) );
  NAND2_X1 U74654 ( .A1(n89094), .A2(n89095), .ZN(n89090) );
  AOI22_X1 U74655 ( .A1(n105727), .A2(n109663), .B1(n105726), .B2(n109667), 
        .ZN(n89095) );
  AOI22_X1 U74656 ( .A1(n86427), .A2(n109669), .B1(n105724), .B2(n109666), 
        .ZN(n89094) );
  NAND2_X1 U74657 ( .A1(n89096), .A2(n89097), .ZN(n89089) );
  AOI22_X1 U74658 ( .A1(n105723), .A2(n72686), .B1(n105722), .B2(n109662), 
        .ZN(n89097) );
  AOI22_X1 U74659 ( .A1(n105721), .A2(n109664), .B1(n105720), .B2(n109668), 
        .ZN(n89096) );
  NAND2_X1 U74660 ( .A1(n89098), .A2(n89099), .ZN(n89088) );
  AOI22_X1 U74661 ( .A1(n105719), .A2(n109674), .B1(n105718), .B2(n72690), 
        .ZN(n89099) );
  AOI22_X1 U74662 ( .A1(n105717), .A2(n72688), .B1(n86440), .B2(n109673), .ZN(
        n89098) );
  NAND2_X1 U74663 ( .A1(n89100), .A2(n89101), .ZN(n89045) );
  NOR4_X1 U74664 ( .A1(n89102), .A2(n89103), .A3(n89104), .A4(n89105), .ZN(
        n89101) );
  NAND2_X1 U74665 ( .A1(n89106), .A2(n89107), .ZN(n89105) );
  AOI22_X1 U74666 ( .A1(n105715), .A2(n72728), .B1(n105714), .B2(n109695), 
        .ZN(n89107) );
  AOI22_X1 U74667 ( .A1(n105713), .A2(n109699), .B1(n105712), .B2(n109698), 
        .ZN(n89106) );
  NAND2_X1 U74668 ( .A1(n89108), .A2(n89109), .ZN(n89104) );
  AOI22_X1 U74669 ( .A1(n86455), .A2(n109704), .B1(n105710), .B2(n109703), 
        .ZN(n89109) );
  AOI22_X1 U74670 ( .A1(n86457), .A2(n109694), .B1(n105708), .B2(n109696), 
        .ZN(n89108) );
  NAND2_X1 U74671 ( .A1(n89110), .A2(n89111), .ZN(n89103) );
  AOI22_X1 U74672 ( .A1(n105707), .A2(n109705), .B1(n105706), .B2(n109701), 
        .ZN(n89111) );
  AOI22_X1 U74673 ( .A1(n105705), .A2(n72732), .B1(n105704), .B2(n72734), .ZN(
        n89110) );
  NAND2_X1 U74674 ( .A1(n89112), .A2(n89113), .ZN(n89102) );
  AOI22_X1 U74675 ( .A1(n105703), .A2(n109708), .B1(n105702), .B2(n72740), 
        .ZN(n89113) );
  AOI22_X1 U74676 ( .A1(n105701), .A2(n109700), .B1(n105700), .B2(n109702), 
        .ZN(n89112) );
  NOR4_X1 U74677 ( .A1(n89114), .A2(n89115), .A3(n89116), .A4(n89117), .ZN(
        n89100) );
  NAND2_X1 U74678 ( .A1(n89118), .A2(n89119), .ZN(n89117) );
  AOI22_X1 U74679 ( .A1(n105699), .A2(n109683), .B1(n105698), .B2(n109688), 
        .ZN(n89119) );
  AOI22_X1 U74680 ( .A1(n86479), .A2(n109682), .B1(n105696), .B2(n72708), .ZN(
        n89118) );
  NAND2_X1 U74681 ( .A1(n89120), .A2(n89121), .ZN(n89116) );
  AOI22_X1 U74682 ( .A1(n105695), .A2(n72717), .B1(n86484), .B2(n109690), .ZN(
        n89121) );
  AOI22_X1 U74683 ( .A1(n105693), .A2(n109691), .B1(n105692), .B2(n109681), 
        .ZN(n89120) );
  NAND2_X1 U74684 ( .A1(n89122), .A2(n89123), .ZN(n89115) );
  AOI22_X1 U74685 ( .A1(n105691), .A2(n109689), .B1(n105690), .B2(n109693), 
        .ZN(n89123) );
  AOI22_X1 U74686 ( .A1(n105689), .A2(n109687), .B1(n105688), .B2(n109692), 
        .ZN(n89122) );
  NAND2_X1 U74687 ( .A1(n89124), .A2(n89125), .ZN(n89114) );
  AOI22_X1 U74688 ( .A1(n86495), .A2(n72722), .B1(n105686), .B2(n109697), .ZN(
        n89125) );
  AOI22_X1 U74689 ( .A1(n105685), .A2(n72720), .B1(n105684), .B2(n109686), 
        .ZN(n89124) );
  NAND2_X1 U74690 ( .A1(n89126), .A2(n89127), .ZN(n89044) );
  NOR4_X1 U74691 ( .A1(n89128), .A2(n89129), .A3(n89130), .A4(n89131), .ZN(
        n89127) );
  NAND2_X1 U74692 ( .A1(n89132), .A2(n89133), .ZN(n89131) );
  AOI22_X1 U74693 ( .A1(n105683), .A2(n109725), .B1(n105682), .B2(n109724), 
        .ZN(n89133) );
  AOI22_X1 U74694 ( .A1(n105681), .A2(n72756), .B1(n105680), .B2(n109722), 
        .ZN(n89132) );
  NAND2_X1 U74695 ( .A1(n89134), .A2(n89135), .ZN(n89130) );
  AOI22_X1 U74696 ( .A1(n105679), .A2(n109720), .B1(n86514), .B2(n109723), 
        .ZN(n89135) );
  AOI22_X1 U74697 ( .A1(n86515), .A2(n72762), .B1(n105677), .B2(n109721), .ZN(
        n89134) );
  NAND2_X1 U74698 ( .A1(n89136), .A2(n89137), .ZN(n89129) );
  AOI22_X1 U74699 ( .A1(n86519), .A2(n109731), .B1(n86520), .B2(n72768), .ZN(
        n89137) );
  AOI22_X1 U74700 ( .A1(n86521), .A2(n109729), .B1(n86522), .B2(n109730), .ZN(
        n89136) );
  NAND2_X1 U74701 ( .A1(n89138), .A2(n89139), .ZN(n89128) );
  AOI22_X1 U74702 ( .A1(n105676), .A2(n109726), .B1(n86526), .B2(n109728), 
        .ZN(n89139) );
  AOI22_X1 U74703 ( .A1(n86527), .A2(n109732), .B1(n86528), .B2(n109727), .ZN(
        n89138) );
  NOR4_X1 U74704 ( .A1(n89140), .A2(n89141), .A3(n89142), .A4(n89143), .ZN(
        n89126) );
  NAND2_X1 U74705 ( .A1(n89144), .A2(n89145), .ZN(n89143) );
  AOI22_X1 U74706 ( .A1(n86535), .A2(n109707), .B1(n105674), .B2(n109711), 
        .ZN(n89145) );
  AOI22_X1 U74707 ( .A1(n105673), .A2(n109710), .B1(n105672), .B2(n72739), 
        .ZN(n89144) );
  NAND2_X1 U74708 ( .A1(n89146), .A2(n89147), .ZN(n89142) );
  AOI22_X1 U74709 ( .A1(n105671), .A2(n109716), .B1(n105670), .B2(n109706), 
        .ZN(n89147) );
  AOI22_X1 U74710 ( .A1(n105669), .A2(n109709), .B1(n86544), .B2(n72745), .ZN(
        n89146) );
  NAND2_X1 U74711 ( .A1(n89148), .A2(n89149), .ZN(n89141) );
  AOI22_X1 U74712 ( .A1(n105667), .A2(n109713), .B1(n105666), .B2(n109717), 
        .ZN(n89149) );
  AOI22_X1 U74713 ( .A1(n105665), .A2(n109719), .B1(n105664), .B2(n109715), 
        .ZN(n89148) );
  NAND2_X1 U74714 ( .A1(n89150), .A2(n89151), .ZN(n89140) );
  AOI22_X1 U74715 ( .A1(n105663), .A2(n72757), .B1(n105662), .B2(n109712), 
        .ZN(n89151) );
  AOI22_X1 U74716 ( .A1(n105661), .A2(n109714), .B1(n86556), .B2(n109718), 
        .ZN(n89150) );
  AOI21_X1 U74717 ( .B1(n86302), .B2(n89153), .A(n89154), .ZN(n89152) );
  OAI21_X1 U74718 ( .B1(n89155), .B2(n105787), .A(n89156), .ZN(n89154) );
  OAI21_X1 U74719 ( .B1(n89157), .B2(n89158), .A(n105786), .ZN(n89156) );
  OAI21_X1 U74720 ( .B1(n109541), .B2(n105785), .A(n89159), .ZN(n89158) );
  AOI22_X1 U74721 ( .A1(n86313), .A2(n72506), .B1(n86314), .B2(n109539), .ZN(
        n89159) );
  NAND2_X1 U74722 ( .A1(n89160), .A2(n89161), .ZN(n89157) );
  AOI22_X1 U74723 ( .A1(n105783), .A2(n109537), .B1(n105782), .B2(n109542), 
        .ZN(n89161) );
  AOI22_X1 U74724 ( .A1(n105781), .A2(n109540), .B1(n105780), .B2(n109538), 
        .ZN(n89160) );
  NOR4_X1 U74725 ( .A1(n89162), .A2(n89163), .A3(n89164), .A4(n89165), .ZN(
        n89155) );
  NAND2_X1 U74726 ( .A1(n89166), .A2(n89167), .ZN(n89165) );
  NOR4_X1 U74727 ( .A1(n89168), .A2(n89169), .A3(n89170), .A4(n89171), .ZN(
        n89167) );
  NAND2_X1 U74728 ( .A1(n89172), .A2(n89173), .ZN(n89171) );
  AOI22_X1 U74729 ( .A1(n105779), .A2(n109518), .B1(n105778), .B2(n109519), 
        .ZN(n89173) );
  AOI22_X1 U74730 ( .A1(n105777), .A2(n109527), .B1(n105776), .B2(n109525), 
        .ZN(n89172) );
  NAND2_X1 U74731 ( .A1(n89174), .A2(n89175), .ZN(n89170) );
  AOI22_X1 U74732 ( .A1(n105775), .A2(n72375), .B1(n105774), .B2(n109522), 
        .ZN(n89175) );
  AOI22_X1 U74733 ( .A1(n105773), .A2(n72479), .B1(n105772), .B2(n109439), 
        .ZN(n89174) );
  NAND2_X1 U74734 ( .A1(n89176), .A2(n89177), .ZN(n89169) );
  AOI22_X1 U74735 ( .A1(n105771), .A2(n109443), .B1(n86346), .B2(n72379), .ZN(
        n89177) );
  AOI22_X1 U74736 ( .A1(n105769), .A2(n109523), .B1(n105768), .B2(n109520), 
        .ZN(n89176) );
  NAND2_X1 U74737 ( .A1(n89178), .A2(n89179), .ZN(n89168) );
  AOI22_X1 U74738 ( .A1(n105767), .A2(n109441), .B1(n105766), .B2(n109445), 
        .ZN(n89179) );
  AOI22_X1 U74739 ( .A1(n105765), .A2(n109444), .B1(n105764), .B2(n72381), 
        .ZN(n89178) );
  NOR4_X1 U74740 ( .A1(n89180), .A2(n89181), .A3(n89182), .A4(n89183), .ZN(
        n89166) );
  NAND2_X1 U74741 ( .A1(n89184), .A2(n89185), .ZN(n89183) );
  AOI22_X1 U74742 ( .A1(n105763), .A2(n109528), .B1(n105762), .B2(n109531), 
        .ZN(n89185) );
  AOI22_X1 U74743 ( .A1(n105761), .A2(n109532), .B1(n86364), .B2(n109534), 
        .ZN(n89184) );
  NAND2_X1 U74744 ( .A1(n89186), .A2(n89187), .ZN(n89182) );
  AOI22_X1 U74745 ( .A1(n105759), .A2(n109533), .B1(n86368), .B2(n109529), 
        .ZN(n89187) );
  AOI22_X1 U74746 ( .A1(n105757), .A2(n109535), .B1(n105756), .B2(n109530), 
        .ZN(n89186) );
  NAND2_X1 U74747 ( .A1(n89188), .A2(n89189), .ZN(n89181) );
  AOI22_X1 U74748 ( .A1(n105755), .A2(n72489), .B1(n105754), .B2(n72488), .ZN(
        n89189) );
  AOI22_X1 U74749 ( .A1(n105753), .A2(n72491), .B1(n105752), .B2(n109536), 
        .ZN(n89188) );
  NAND2_X1 U74750 ( .A1(n89190), .A2(n89191), .ZN(n89180) );
  AOI22_X1 U74751 ( .A1(n105751), .A2(n109521), .B1(n105750), .B2(n109526), 
        .ZN(n89191) );
  AOI22_X1 U74752 ( .A1(n105749), .A2(n72486), .B1(n86382), .B2(n109524), .ZN(
        n89190) );
  NAND2_X1 U74753 ( .A1(n89192), .A2(n89193), .ZN(n89164) );
  NOR4_X1 U74754 ( .A1(n89194), .A2(n89195), .A3(n89196), .A4(n89197), .ZN(
        n89193) );
  NAND2_X1 U74755 ( .A1(n89198), .A2(n89199), .ZN(n89197) );
  AOI22_X1 U74756 ( .A1(n105747), .A2(n109454), .B1(n105746), .B2(n109456), 
        .ZN(n89199) );
  AOI22_X1 U74757 ( .A1(n105745), .A2(n72404), .B1(n105744), .B2(n109455), 
        .ZN(n89198) );
  NAND2_X1 U74758 ( .A1(n89200), .A2(n89201), .ZN(n89196) );
  AOI22_X1 U74759 ( .A1(n105743), .A2(n72408), .B1(n105742), .B2(n72410), .ZN(
        n89201) );
  AOI22_X1 U74760 ( .A1(n105741), .A2(n109462), .B1(n86400), .B2(n109463), 
        .ZN(n89200) );
  NAND2_X1 U74761 ( .A1(n89202), .A2(n89203), .ZN(n89195) );
  AOI22_X1 U74762 ( .A1(n105739), .A2(n109459), .B1(n105738), .B2(n109461), 
        .ZN(n89203) );
  AOI22_X1 U74763 ( .A1(n105737), .A2(n109464), .B1(n86406), .B2(n109460), 
        .ZN(n89202) );
  NAND2_X1 U74764 ( .A1(n89204), .A2(n89205), .ZN(n89194) );
  AOI22_X1 U74765 ( .A1(n105735), .A2(n109469), .B1(n105734), .B2(n72415), 
        .ZN(n89205) );
  AOI22_X1 U74766 ( .A1(n105733), .A2(n109468), .B1(n105732), .B2(n72413), 
        .ZN(n89204) );
  NOR4_X1 U74767 ( .A1(n89206), .A2(n89207), .A3(n89208), .A4(n89209), .ZN(
        n89192) );
  NAND2_X1 U74768 ( .A1(n89210), .A2(n89211), .ZN(n89209) );
  AOI22_X1 U74769 ( .A1(n105731), .A2(n109449), .B1(n105730), .B2(n109440), 
        .ZN(n89211) );
  AOI22_X1 U74770 ( .A1(n105729), .A2(n109442), .B1(n105728), .B2(n72387), 
        .ZN(n89210) );
  NAND2_X1 U74771 ( .A1(n89212), .A2(n89213), .ZN(n89208) );
  AOI22_X1 U74772 ( .A1(n105727), .A2(n109447), .B1(n86426), .B2(n109451), 
        .ZN(n89213) );
  AOI22_X1 U74773 ( .A1(n86427), .A2(n109453), .B1(n86428), .B2(n109450), .ZN(
        n89212) );
  NAND2_X1 U74774 ( .A1(n89214), .A2(n89215), .ZN(n89207) );
  AOI22_X1 U74775 ( .A1(n105723), .A2(n72396), .B1(n105722), .B2(n109446), 
        .ZN(n89215) );
  AOI22_X1 U74776 ( .A1(n105721), .A2(n109448), .B1(n105720), .B2(n109452), 
        .ZN(n89214) );
  NAND2_X1 U74777 ( .A1(n89216), .A2(n89217), .ZN(n89206) );
  AOI22_X1 U74778 ( .A1(n105719), .A2(n109458), .B1(n105718), .B2(n72400), 
        .ZN(n89217) );
  AOI22_X1 U74779 ( .A1(n105717), .A2(n72398), .B1(n86440), .B2(n109457), .ZN(
        n89216) );
  NAND2_X1 U74780 ( .A1(n89218), .A2(n89219), .ZN(n89163) );
  NOR4_X1 U74781 ( .A1(n89220), .A2(n89221), .A3(n89222), .A4(n89223), .ZN(
        n89219) );
  NAND2_X1 U74782 ( .A1(n89224), .A2(n89225), .ZN(n89223) );
  AOI22_X1 U74783 ( .A1(n105715), .A2(n72438), .B1(n86450), .B2(n109479), .ZN(
        n89225) );
  AOI22_X1 U74784 ( .A1(n105713), .A2(n109483), .B1(n105712), .B2(n109482), 
        .ZN(n89224) );
  NAND2_X1 U74785 ( .A1(n89226), .A2(n89227), .ZN(n89222) );
  AOI22_X1 U74786 ( .A1(n86455), .A2(n109488), .B1(n105710), .B2(n109487), 
        .ZN(n89227) );
  AOI22_X1 U74787 ( .A1(n86457), .A2(n109478), .B1(n105708), .B2(n109480), 
        .ZN(n89226) );
  NAND2_X1 U74788 ( .A1(n89228), .A2(n89229), .ZN(n89221) );
  AOI22_X1 U74789 ( .A1(n105707), .A2(n109489), .B1(n105706), .B2(n109485), 
        .ZN(n89229) );
  AOI22_X1 U74790 ( .A1(n105705), .A2(n72442), .B1(n105704), .B2(n72444), .ZN(
        n89228) );
  NAND2_X1 U74791 ( .A1(n89230), .A2(n89231), .ZN(n89220) );
  AOI22_X1 U74792 ( .A1(n105703), .A2(n109492), .B1(n105702), .B2(n72450), 
        .ZN(n89231) );
  AOI22_X1 U74793 ( .A1(n105701), .A2(n109484), .B1(n105700), .B2(n109486), 
        .ZN(n89230) );
  NOR4_X1 U74794 ( .A1(n89232), .A2(n89233), .A3(n89234), .A4(n89235), .ZN(
        n89218) );
  NAND2_X1 U74795 ( .A1(n89236), .A2(n89237), .ZN(n89235) );
  AOI22_X1 U74796 ( .A1(n105699), .A2(n109467), .B1(n105698), .B2(n109472), 
        .ZN(n89237) );
  AOI22_X1 U74797 ( .A1(n86479), .A2(n109466), .B1(n105696), .B2(n72418), .ZN(
        n89236) );
  NAND2_X1 U74798 ( .A1(n89238), .A2(n89239), .ZN(n89234) );
  AOI22_X1 U74799 ( .A1(n105695), .A2(n72427), .B1(n86484), .B2(n109474), .ZN(
        n89239) );
  AOI22_X1 U74800 ( .A1(n105693), .A2(n109475), .B1(n105692), .B2(n109465), 
        .ZN(n89238) );
  NAND2_X1 U74801 ( .A1(n89240), .A2(n89241), .ZN(n89233) );
  AOI22_X1 U74802 ( .A1(n105691), .A2(n109473), .B1(n86490), .B2(n109477), 
        .ZN(n89241) );
  AOI22_X1 U74803 ( .A1(n105689), .A2(n109471), .B1(n105688), .B2(n109476), 
        .ZN(n89240) );
  NAND2_X1 U74804 ( .A1(n89242), .A2(n89243), .ZN(n89232) );
  AOI22_X1 U74805 ( .A1(n86495), .A2(n72432), .B1(n105686), .B2(n109481), .ZN(
        n89243) );
  AOI22_X1 U74806 ( .A1(n105685), .A2(n72430), .B1(n105684), .B2(n109470), 
        .ZN(n89242) );
  NAND2_X1 U74807 ( .A1(n89244), .A2(n89245), .ZN(n89162) );
  NOR4_X1 U74808 ( .A1(n89246), .A2(n89247), .A3(n89248), .A4(n89249), .ZN(
        n89245) );
  NAND2_X1 U74809 ( .A1(n89250), .A2(n89251), .ZN(n89249) );
  AOI22_X1 U74810 ( .A1(n105683), .A2(n109510), .B1(n105682), .B2(n109509), 
        .ZN(n89251) );
  AOI22_X1 U74811 ( .A1(n105681), .A2(n72466), .B1(n105680), .B2(n109507), 
        .ZN(n89250) );
  NAND2_X1 U74812 ( .A1(n89252), .A2(n89253), .ZN(n89248) );
  AOI22_X1 U74813 ( .A1(n105679), .A2(n109505), .B1(n86514), .B2(n109508), 
        .ZN(n89253) );
  AOI22_X1 U74814 ( .A1(n86515), .A2(n72472), .B1(n86516), .B2(n109506), .ZN(
        n89252) );
  NAND2_X1 U74815 ( .A1(n89254), .A2(n89255), .ZN(n89247) );
  AOI22_X1 U74816 ( .A1(n86519), .A2(n109516), .B1(n86520), .B2(n72478), .ZN(
        n89255) );
  AOI22_X1 U74817 ( .A1(n86521), .A2(n109514), .B1(n86522), .B2(n109515), .ZN(
        n89254) );
  NAND2_X1 U74818 ( .A1(n89256), .A2(n89257), .ZN(n89246) );
  AOI22_X1 U74819 ( .A1(n105676), .A2(n109511), .B1(n86526), .B2(n109513), 
        .ZN(n89257) );
  AOI22_X1 U74820 ( .A1(n86527), .A2(n109517), .B1(n86528), .B2(n109512), .ZN(
        n89256) );
  NOR4_X1 U74821 ( .A1(n89258), .A2(n89259), .A3(n89260), .A4(n89261), .ZN(
        n89244) );
  NAND2_X1 U74822 ( .A1(n89262), .A2(n89263), .ZN(n89261) );
  AOI22_X1 U74823 ( .A1(n86535), .A2(n109491), .B1(n105674), .B2(n109495), 
        .ZN(n89263) );
  AOI22_X1 U74824 ( .A1(n105673), .A2(n109494), .B1(n105672), .B2(n72449), 
        .ZN(n89262) );
  NAND2_X1 U74825 ( .A1(n89264), .A2(n89265), .ZN(n89260) );
  AOI22_X1 U74826 ( .A1(n105671), .A2(n109501), .B1(n105670), .B2(n109490), 
        .ZN(n89265) );
  AOI22_X1 U74827 ( .A1(n105669), .A2(n109493), .B1(n86544), .B2(n109498), 
        .ZN(n89264) );
  NAND2_X1 U74828 ( .A1(n89266), .A2(n89267), .ZN(n89259) );
  AOI22_X1 U74829 ( .A1(n105667), .A2(n109497), .B1(n105666), .B2(n109502), 
        .ZN(n89267) );
  AOI22_X1 U74830 ( .A1(n105665), .A2(n109504), .B1(n105664), .B2(n109500), 
        .ZN(n89266) );
  NAND2_X1 U74831 ( .A1(n89268), .A2(n89269), .ZN(n89258) );
  AOI22_X1 U74832 ( .A1(n105663), .A2(n72467), .B1(n105662), .B2(n109496), 
        .ZN(n89269) );
  AOI22_X1 U74833 ( .A1(n86555), .A2(n109499), .B1(n86556), .B2(n109503), .ZN(
        n89268) );
  AOI21_X1 U74834 ( .B1(n86302), .B2(n89271), .A(n89272), .ZN(n89270) );
  OAI21_X1 U74835 ( .B1(n89273), .B2(n105787), .A(n89274), .ZN(n89272) );
  OAI21_X1 U74836 ( .B1(n89275), .B2(n89276), .A(n86310), .ZN(n89274) );
  OAI21_X1 U74837 ( .B1(n109079), .B2(n105785), .A(n89277), .ZN(n89276) );
  AOI22_X1 U74838 ( .A1(n86313), .A2(n71906), .B1(n86314), .B2(n109077), .ZN(
        n89277) );
  NAND2_X1 U74839 ( .A1(n89278), .A2(n89279), .ZN(n89275) );
  AOI22_X1 U74840 ( .A1(n105783), .A2(n109075), .B1(n105782), .B2(n109080), 
        .ZN(n89279) );
  AOI22_X1 U74841 ( .A1(n105781), .A2(n109078), .B1(n105780), .B2(n109076), 
        .ZN(n89278) );
  NOR4_X1 U74842 ( .A1(n89280), .A2(n89281), .A3(n89282), .A4(n89283), .ZN(
        n89273) );
  NAND2_X1 U74843 ( .A1(n89284), .A2(n89285), .ZN(n89283) );
  NOR4_X1 U74844 ( .A1(n89286), .A2(n89287), .A3(n89288), .A4(n89289), .ZN(
        n89285) );
  NAND2_X1 U74845 ( .A1(n89290), .A2(n89291), .ZN(n89289) );
  AOI22_X1 U74846 ( .A1(n105779), .A2(n109056), .B1(n105778), .B2(n109057), 
        .ZN(n89291) );
  AOI22_X1 U74847 ( .A1(n105777), .A2(n109065), .B1(n105776), .B2(n109063), 
        .ZN(n89290) );
  NAND2_X1 U74848 ( .A1(n89292), .A2(n89293), .ZN(n89288) );
  AOI22_X1 U74849 ( .A1(n105775), .A2(n71775), .B1(n105774), .B2(n109060), 
        .ZN(n89293) );
  AOI22_X1 U74850 ( .A1(n105773), .A2(n71879), .B1(n105772), .B2(n108976), 
        .ZN(n89292) );
  NAND2_X1 U74851 ( .A1(n89294), .A2(n89295), .ZN(n89287) );
  AOI22_X1 U74852 ( .A1(n105771), .A2(n108980), .B1(n105770), .B2(n71779), 
        .ZN(n89295) );
  AOI22_X1 U74853 ( .A1(n105769), .A2(n109061), .B1(n105768), .B2(n109058), 
        .ZN(n89294) );
  NAND2_X1 U74854 ( .A1(n89296), .A2(n89297), .ZN(n89286) );
  AOI22_X1 U74855 ( .A1(n105767), .A2(n108978), .B1(n105766), .B2(n108982), 
        .ZN(n89297) );
  AOI22_X1 U74856 ( .A1(n105765), .A2(n108981), .B1(n105764), .B2(n71781), 
        .ZN(n89296) );
  NOR4_X1 U74857 ( .A1(n89298), .A2(n89299), .A3(n89300), .A4(n89301), .ZN(
        n89284) );
  NAND2_X1 U74858 ( .A1(n89302), .A2(n89303), .ZN(n89301) );
  AOI22_X1 U74859 ( .A1(n105763), .A2(n109066), .B1(n105762), .B2(n109069), 
        .ZN(n89303) );
  AOI22_X1 U74860 ( .A1(n105761), .A2(n109070), .B1(n86364), .B2(n109072), 
        .ZN(n89302) );
  NAND2_X1 U74861 ( .A1(n89304), .A2(n89305), .ZN(n89300) );
  AOI22_X1 U74862 ( .A1(n105759), .A2(n109071), .B1(n105758), .B2(n109067), 
        .ZN(n89305) );
  AOI22_X1 U74863 ( .A1(n105757), .A2(n109073), .B1(n105756), .B2(n109068), 
        .ZN(n89304) );
  NAND2_X1 U74864 ( .A1(n89306), .A2(n89307), .ZN(n89299) );
  AOI22_X1 U74865 ( .A1(n105755), .A2(n71889), .B1(n105754), .B2(n71888), .ZN(
        n89307) );
  AOI22_X1 U74866 ( .A1(n105753), .A2(n71891), .B1(n105752), .B2(n109074), 
        .ZN(n89306) );
  NAND2_X1 U74867 ( .A1(n89308), .A2(n89309), .ZN(n89298) );
  AOI22_X1 U74868 ( .A1(n105751), .A2(n109059), .B1(n105750), .B2(n109064), 
        .ZN(n89309) );
  AOI22_X1 U74869 ( .A1(n105749), .A2(n71886), .B1(n86382), .B2(n109062), .ZN(
        n89308) );
  NAND2_X1 U74870 ( .A1(n89310), .A2(n89311), .ZN(n89282) );
  NOR4_X1 U74871 ( .A1(n89312), .A2(n89313), .A3(n89314), .A4(n89315), .ZN(
        n89311) );
  NAND2_X1 U74872 ( .A1(n89316), .A2(n89317), .ZN(n89315) );
  AOI22_X1 U74873 ( .A1(n105747), .A2(n108991), .B1(n105746), .B2(n108993), 
        .ZN(n89317) );
  AOI22_X1 U74874 ( .A1(n105745), .A2(n71804), .B1(n105744), .B2(n108992), 
        .ZN(n89316) );
  NAND2_X1 U74875 ( .A1(n89318), .A2(n89319), .ZN(n89314) );
  AOI22_X1 U74876 ( .A1(n105743), .A2(n71808), .B1(n105742), .B2(n71810), .ZN(
        n89319) );
  AOI22_X1 U74877 ( .A1(n105741), .A2(n108999), .B1(n105740), .B2(n109000), 
        .ZN(n89318) );
  NAND2_X1 U74878 ( .A1(n89320), .A2(n89321), .ZN(n89313) );
  AOI22_X1 U74879 ( .A1(n105739), .A2(n108996), .B1(n105738), .B2(n108998), 
        .ZN(n89321) );
  AOI22_X1 U74880 ( .A1(n105737), .A2(n109001), .B1(n86406), .B2(n108997), 
        .ZN(n89320) );
  NAND2_X1 U74881 ( .A1(n89322), .A2(n89323), .ZN(n89312) );
  AOI22_X1 U74882 ( .A1(n105735), .A2(n109006), .B1(n105734), .B2(n71815), 
        .ZN(n89323) );
  AOI22_X1 U74883 ( .A1(n105733), .A2(n109005), .B1(n105732), .B2(n71813), 
        .ZN(n89322) );
  NOR4_X1 U74884 ( .A1(n89324), .A2(n89325), .A3(n89326), .A4(n89327), .ZN(
        n89310) );
  NAND2_X1 U74885 ( .A1(n89328), .A2(n89329), .ZN(n89327) );
  AOI22_X1 U74886 ( .A1(n105731), .A2(n108986), .B1(n105730), .B2(n108977), 
        .ZN(n89329) );
  AOI22_X1 U74887 ( .A1(n105729), .A2(n108979), .B1(n105728), .B2(n71787), 
        .ZN(n89328) );
  NAND2_X1 U74888 ( .A1(n89330), .A2(n89331), .ZN(n89326) );
  AOI22_X1 U74889 ( .A1(n105727), .A2(n108984), .B1(n105726), .B2(n108988), 
        .ZN(n89331) );
  AOI22_X1 U74890 ( .A1(n86427), .A2(n108990), .B1(n105724), .B2(n108987), 
        .ZN(n89330) );
  NAND2_X1 U74891 ( .A1(n89332), .A2(n89333), .ZN(n89325) );
  AOI22_X1 U74892 ( .A1(n105723), .A2(n71796), .B1(n105722), .B2(n108983), 
        .ZN(n89333) );
  AOI22_X1 U74893 ( .A1(n105721), .A2(n108985), .B1(n105720), .B2(n108989), 
        .ZN(n89332) );
  NAND2_X1 U74894 ( .A1(n89334), .A2(n89335), .ZN(n89324) );
  AOI22_X1 U74895 ( .A1(n105719), .A2(n108995), .B1(n105718), .B2(n71800), 
        .ZN(n89335) );
  AOI22_X1 U74896 ( .A1(n105717), .A2(n71798), .B1(n86440), .B2(n108994), .ZN(
        n89334) );
  NAND2_X1 U74897 ( .A1(n89336), .A2(n89337), .ZN(n89281) );
  NOR4_X1 U74898 ( .A1(n89338), .A2(n89339), .A3(n89340), .A4(n89341), .ZN(
        n89337) );
  NAND2_X1 U74899 ( .A1(n89342), .A2(n89343), .ZN(n89341) );
  AOI22_X1 U74900 ( .A1(n105715), .A2(n71838), .B1(n105714), .B2(n109016), 
        .ZN(n89343) );
  AOI22_X1 U74901 ( .A1(n105713), .A2(n109020), .B1(n105712), .B2(n109019), 
        .ZN(n89342) );
  NAND2_X1 U74902 ( .A1(n89344), .A2(n89345), .ZN(n89340) );
  AOI22_X1 U74903 ( .A1(n86455), .A2(n109025), .B1(n105710), .B2(n109024), 
        .ZN(n89345) );
  AOI22_X1 U74904 ( .A1(n86457), .A2(n109015), .B1(n105708), .B2(n109017), 
        .ZN(n89344) );
  NAND2_X1 U74905 ( .A1(n89346), .A2(n89347), .ZN(n89339) );
  AOI22_X1 U74906 ( .A1(n105707), .A2(n109026), .B1(n105706), .B2(n109022), 
        .ZN(n89347) );
  AOI22_X1 U74907 ( .A1(n105705), .A2(n71842), .B1(n105704), .B2(n71844), .ZN(
        n89346) );
  NAND2_X1 U74908 ( .A1(n89348), .A2(n89349), .ZN(n89338) );
  AOI22_X1 U74909 ( .A1(n105703), .A2(n109029), .B1(n105702), .B2(n71850), 
        .ZN(n89349) );
  AOI22_X1 U74910 ( .A1(n105701), .A2(n109021), .B1(n105700), .B2(n109023), 
        .ZN(n89348) );
  NOR4_X1 U74911 ( .A1(n89350), .A2(n89351), .A3(n89352), .A4(n89353), .ZN(
        n89336) );
  NAND2_X1 U74912 ( .A1(n89354), .A2(n89355), .ZN(n89353) );
  AOI22_X1 U74913 ( .A1(n105699), .A2(n109004), .B1(n105698), .B2(n109009), 
        .ZN(n89355) );
  AOI22_X1 U74914 ( .A1(n86479), .A2(n109003), .B1(n105696), .B2(n71818), .ZN(
        n89354) );
  NAND2_X1 U74915 ( .A1(n89356), .A2(n89357), .ZN(n89352) );
  AOI22_X1 U74916 ( .A1(n105695), .A2(n71827), .B1(n86484), .B2(n109011), .ZN(
        n89357) );
  AOI22_X1 U74917 ( .A1(n105693), .A2(n109012), .B1(n105692), .B2(n109002), 
        .ZN(n89356) );
  NAND2_X1 U74918 ( .A1(n89358), .A2(n89359), .ZN(n89351) );
  AOI22_X1 U74919 ( .A1(n105691), .A2(n109010), .B1(n105690), .B2(n109014), 
        .ZN(n89359) );
  AOI22_X1 U74920 ( .A1(n105689), .A2(n109008), .B1(n105688), .B2(n109013), 
        .ZN(n89358) );
  NAND2_X1 U74921 ( .A1(n89360), .A2(n89361), .ZN(n89350) );
  AOI22_X1 U74922 ( .A1(n86495), .A2(n71832), .B1(n105686), .B2(n109018), .ZN(
        n89361) );
  AOI22_X1 U74923 ( .A1(n105685), .A2(n71830), .B1(n105684), .B2(n109007), 
        .ZN(n89360) );
  NAND2_X1 U74924 ( .A1(n89362), .A2(n89363), .ZN(n89280) );
  NOR4_X1 U74925 ( .A1(n89364), .A2(n89365), .A3(n89366), .A4(n89367), .ZN(
        n89363) );
  NAND2_X1 U74926 ( .A1(n89368), .A2(n89369), .ZN(n89367) );
  AOI22_X1 U74927 ( .A1(n105683), .A2(n109047), .B1(n105682), .B2(n109046), 
        .ZN(n89369) );
  AOI22_X1 U74928 ( .A1(n105681), .A2(n71866), .B1(n105680), .B2(n109044), 
        .ZN(n89368) );
  NAND2_X1 U74929 ( .A1(n89370), .A2(n89371), .ZN(n89366) );
  AOI22_X1 U74930 ( .A1(n105679), .A2(n109042), .B1(n86514), .B2(n109045), 
        .ZN(n89371) );
  AOI22_X1 U74931 ( .A1(n86515), .A2(n71872), .B1(n105677), .B2(n109043), .ZN(
        n89370) );
  NAND2_X1 U74932 ( .A1(n89372), .A2(n89373), .ZN(n89365) );
  AOI22_X1 U74933 ( .A1(n86519), .A2(n109053), .B1(n86520), .B2(n71878), .ZN(
        n89373) );
  AOI22_X1 U74934 ( .A1(n86521), .A2(n109051), .B1(n86522), .B2(n109052), .ZN(
        n89372) );
  NAND2_X1 U74935 ( .A1(n89374), .A2(n89375), .ZN(n89364) );
  AOI22_X1 U74936 ( .A1(n105676), .A2(n109048), .B1(n86526), .B2(n109050), 
        .ZN(n89375) );
  AOI22_X1 U74937 ( .A1(n86527), .A2(n109054), .B1(n86528), .B2(n109049), .ZN(
        n89374) );
  NOR4_X1 U74938 ( .A1(n89376), .A2(n89377), .A3(n89378), .A4(n89379), .ZN(
        n89362) );
  NAND2_X1 U74939 ( .A1(n89380), .A2(n89381), .ZN(n89379) );
  AOI22_X1 U74940 ( .A1(n86535), .A2(n109028), .B1(n105674), .B2(n109032), 
        .ZN(n89381) );
  AOI22_X1 U74941 ( .A1(n105673), .A2(n109031), .B1(n105672), .B2(n71849), 
        .ZN(n89380) );
  NAND2_X1 U74942 ( .A1(n89382), .A2(n89383), .ZN(n89378) );
  AOI22_X1 U74943 ( .A1(n105671), .A2(n109038), .B1(n105670), .B2(n109027), 
        .ZN(n89383) );
  AOI22_X1 U74944 ( .A1(n105669), .A2(n109030), .B1(n86544), .B2(n109035), 
        .ZN(n89382) );
  NAND2_X1 U74945 ( .A1(n89384), .A2(n89385), .ZN(n89377) );
  AOI22_X1 U74946 ( .A1(n105667), .A2(n109034), .B1(n105666), .B2(n109039), 
        .ZN(n89385) );
  AOI22_X1 U74947 ( .A1(n105665), .A2(n109041), .B1(n105664), .B2(n109037), 
        .ZN(n89384) );
  NAND2_X1 U74948 ( .A1(n89386), .A2(n89387), .ZN(n89376) );
  AOI22_X1 U74949 ( .A1(n105663), .A2(n71867), .B1(n105662), .B2(n109033), 
        .ZN(n89387) );
  AOI22_X1 U74950 ( .A1(n105661), .A2(n109036), .B1(n105660), .B2(n109040), 
        .ZN(n89386) );
  AOI21_X1 U74951 ( .B1(n86302), .B2(n81792), .A(n89389), .ZN(n89388) );
  OAI21_X1 U74952 ( .B1(n89390), .B2(n105787), .A(n89391), .ZN(n89389) );
  OAI21_X1 U74953 ( .B1(n89392), .B2(n89393), .A(n86310), .ZN(n89391) );
  OAI21_X1 U74954 ( .B1(n109426), .B2(n105785), .A(n89394), .ZN(n89393) );
  AOI22_X1 U74955 ( .A1(n86313), .A2(n72355), .B1(n86314), .B2(n109424), .ZN(
        n89394) );
  NAND2_X1 U74956 ( .A1(n89395), .A2(n89396), .ZN(n89392) );
  AOI22_X1 U74957 ( .A1(n105783), .A2(n109422), .B1(n105782), .B2(n109427), 
        .ZN(n89396) );
  AOI22_X1 U74958 ( .A1(n105781), .A2(n109425), .B1(n105780), .B2(n109423), 
        .ZN(n89395) );
  NOR4_X1 U74959 ( .A1(n89397), .A2(n89398), .A3(n89399), .A4(n89400), .ZN(
        n89390) );
  NAND2_X1 U74960 ( .A1(n89401), .A2(n89402), .ZN(n89400) );
  NOR4_X1 U74961 ( .A1(n89403), .A2(n89404), .A3(n89405), .A4(n89406), .ZN(
        n89402) );
  NAND2_X1 U74962 ( .A1(n89407), .A2(n89408), .ZN(n89406) );
  AOI22_X1 U74963 ( .A1(n105779), .A2(n109403), .B1(n105778), .B2(n109404), 
        .ZN(n89408) );
  AOI22_X1 U74964 ( .A1(n105777), .A2(n109412), .B1(n105776), .B2(n109410), 
        .ZN(n89407) );
  NAND2_X1 U74965 ( .A1(n89409), .A2(n89410), .ZN(n89405) );
  AOI22_X1 U74966 ( .A1(n105775), .A2(n72224), .B1(n105774), .B2(n109407), 
        .ZN(n89410) );
  AOI22_X1 U74967 ( .A1(n105773), .A2(n72328), .B1(n105772), .B2(n109324), 
        .ZN(n89409) );
  NAND2_X1 U74968 ( .A1(n89411), .A2(n89412), .ZN(n89404) );
  AOI22_X1 U74969 ( .A1(n105771), .A2(n109328), .B1(n105770), .B2(n72228), 
        .ZN(n89412) );
  AOI22_X1 U74970 ( .A1(n105769), .A2(n109408), .B1(n105768), .B2(n109405), 
        .ZN(n89411) );
  NAND2_X1 U74971 ( .A1(n89413), .A2(n89414), .ZN(n89403) );
  AOI22_X1 U74972 ( .A1(n105767), .A2(n109326), .B1(n105766), .B2(n109330), 
        .ZN(n89414) );
  AOI22_X1 U74973 ( .A1(n105765), .A2(n109329), .B1(n105764), .B2(n72230), 
        .ZN(n89413) );
  NOR4_X1 U74974 ( .A1(n89415), .A2(n89416), .A3(n89417), .A4(n89418), .ZN(
        n89401) );
  NAND2_X1 U74975 ( .A1(n89419), .A2(n89420), .ZN(n89418) );
  AOI22_X1 U74976 ( .A1(n105763), .A2(n109413), .B1(n105762), .B2(n109416), 
        .ZN(n89420) );
  AOI22_X1 U74977 ( .A1(n105761), .A2(n109417), .B1(n86364), .B2(n109419), 
        .ZN(n89419) );
  NAND2_X1 U74978 ( .A1(n89421), .A2(n89422), .ZN(n89417) );
  AOI22_X1 U74979 ( .A1(n105759), .A2(n109418), .B1(n105758), .B2(n109414), 
        .ZN(n89422) );
  AOI22_X1 U74980 ( .A1(n105757), .A2(n109420), .B1(n105756), .B2(n109415), 
        .ZN(n89421) );
  NAND2_X1 U74981 ( .A1(n89423), .A2(n89424), .ZN(n89416) );
  AOI22_X1 U74982 ( .A1(n105755), .A2(n72338), .B1(n105754), .B2(n72337), .ZN(
        n89424) );
  AOI22_X1 U74983 ( .A1(n105753), .A2(n72340), .B1(n105752), .B2(n109421), 
        .ZN(n89423) );
  NAND2_X1 U74984 ( .A1(n89425), .A2(n89426), .ZN(n89415) );
  AOI22_X1 U74985 ( .A1(n105751), .A2(n109406), .B1(n105750), .B2(n109411), 
        .ZN(n89426) );
  AOI22_X1 U74986 ( .A1(n105749), .A2(n72335), .B1(n86382), .B2(n109409), .ZN(
        n89425) );
  NAND2_X1 U74987 ( .A1(n89427), .A2(n89428), .ZN(n89399) );
  NOR4_X1 U74988 ( .A1(n89429), .A2(n89430), .A3(n89431), .A4(n89432), .ZN(
        n89428) );
  NAND2_X1 U74989 ( .A1(n89433), .A2(n89434), .ZN(n89432) );
  AOI22_X1 U74990 ( .A1(n105747), .A2(n109339), .B1(n105746), .B2(n109341), 
        .ZN(n89434) );
  AOI22_X1 U74991 ( .A1(n105745), .A2(n72253), .B1(n105744), .B2(n109340), 
        .ZN(n89433) );
  NAND2_X1 U74992 ( .A1(n89435), .A2(n89436), .ZN(n89431) );
  AOI22_X1 U74993 ( .A1(n105743), .A2(n72257), .B1(n105742), .B2(n72259), .ZN(
        n89436) );
  AOI22_X1 U74994 ( .A1(n105741), .A2(n109347), .B1(n105740), .B2(n109348), 
        .ZN(n89435) );
  NAND2_X1 U74995 ( .A1(n89437), .A2(n89438), .ZN(n89430) );
  AOI22_X1 U74996 ( .A1(n105739), .A2(n109344), .B1(n105738), .B2(n109346), 
        .ZN(n89438) );
  AOI22_X1 U74997 ( .A1(n105737), .A2(n109349), .B1(n86406), .B2(n109345), 
        .ZN(n89437) );
  NAND2_X1 U74998 ( .A1(n89439), .A2(n89440), .ZN(n89429) );
  AOI22_X1 U74999 ( .A1(n105735), .A2(n109354), .B1(n105734), .B2(n72264), 
        .ZN(n89440) );
  AOI22_X1 U75000 ( .A1(n105733), .A2(n109353), .B1(n105732), .B2(n72262), 
        .ZN(n89439) );
  NOR4_X1 U75001 ( .A1(n89441), .A2(n89442), .A3(n89443), .A4(n89444), .ZN(
        n89427) );
  NAND2_X1 U75002 ( .A1(n89445), .A2(n89446), .ZN(n89444) );
  AOI22_X1 U75003 ( .A1(n105731), .A2(n109334), .B1(n105730), .B2(n109325), 
        .ZN(n89446) );
  AOI22_X1 U75004 ( .A1(n105729), .A2(n109327), .B1(n105728), .B2(n72236), 
        .ZN(n89445) );
  NAND2_X1 U75005 ( .A1(n89447), .A2(n89448), .ZN(n89443) );
  AOI22_X1 U75006 ( .A1(n105727), .A2(n109332), .B1(n105726), .B2(n109336), 
        .ZN(n89448) );
  AOI22_X1 U75007 ( .A1(n86427), .A2(n109338), .B1(n105724), .B2(n109335), 
        .ZN(n89447) );
  NAND2_X1 U75008 ( .A1(n89449), .A2(n89450), .ZN(n89442) );
  AOI22_X1 U75009 ( .A1(n105723), .A2(n72245), .B1(n105722), .B2(n109331), 
        .ZN(n89450) );
  AOI22_X1 U75010 ( .A1(n105721), .A2(n109333), .B1(n105720), .B2(n109337), 
        .ZN(n89449) );
  NAND2_X1 U75011 ( .A1(n89451), .A2(n89452), .ZN(n89441) );
  AOI22_X1 U75012 ( .A1(n105719), .A2(n109343), .B1(n105718), .B2(n72249), 
        .ZN(n89452) );
  AOI22_X1 U75013 ( .A1(n105717), .A2(n72247), .B1(n86440), .B2(n109342), .ZN(
        n89451) );
  NAND2_X1 U75014 ( .A1(n89453), .A2(n89454), .ZN(n89398) );
  NOR4_X1 U75015 ( .A1(n89455), .A2(n89456), .A3(n89457), .A4(n89458), .ZN(
        n89454) );
  NAND2_X1 U75016 ( .A1(n89459), .A2(n89460), .ZN(n89458) );
  AOI22_X1 U75017 ( .A1(n105715), .A2(n72287), .B1(n105714), .B2(n109364), 
        .ZN(n89460) );
  AOI22_X1 U75018 ( .A1(n105713), .A2(n109368), .B1(n105712), .B2(n109367), 
        .ZN(n89459) );
  NAND2_X1 U75019 ( .A1(n89461), .A2(n89462), .ZN(n89457) );
  AOI22_X1 U75020 ( .A1(n86455), .A2(n109373), .B1(n105710), .B2(n109372), 
        .ZN(n89462) );
  AOI22_X1 U75021 ( .A1(n86457), .A2(n109363), .B1(n105708), .B2(n109365), 
        .ZN(n89461) );
  NAND2_X1 U75022 ( .A1(n89463), .A2(n89464), .ZN(n89456) );
  AOI22_X1 U75023 ( .A1(n105707), .A2(n109374), .B1(n105706), .B2(n109370), 
        .ZN(n89464) );
  AOI22_X1 U75024 ( .A1(n105705), .A2(n72291), .B1(n105704), .B2(n72293), .ZN(
        n89463) );
  NAND2_X1 U75025 ( .A1(n89465), .A2(n89466), .ZN(n89455) );
  AOI22_X1 U75026 ( .A1(n105703), .A2(n109377), .B1(n105702), .B2(n72299), 
        .ZN(n89466) );
  AOI22_X1 U75027 ( .A1(n105701), .A2(n109369), .B1(n105700), .B2(n109371), 
        .ZN(n89465) );
  NOR4_X1 U75028 ( .A1(n89467), .A2(n89468), .A3(n89469), .A4(n89470), .ZN(
        n89453) );
  NAND2_X1 U75029 ( .A1(n89471), .A2(n89472), .ZN(n89470) );
  AOI22_X1 U75030 ( .A1(n105699), .A2(n109352), .B1(n105698), .B2(n109357), 
        .ZN(n89472) );
  AOI22_X1 U75031 ( .A1(n86479), .A2(n109351), .B1(n105696), .B2(n72267), .ZN(
        n89471) );
  NAND2_X1 U75032 ( .A1(n89473), .A2(n89474), .ZN(n89469) );
  AOI22_X1 U75033 ( .A1(n105695), .A2(n72276), .B1(n86484), .B2(n109359), .ZN(
        n89474) );
  AOI22_X1 U75034 ( .A1(n105693), .A2(n109360), .B1(n105692), .B2(n109350), 
        .ZN(n89473) );
  NAND2_X1 U75035 ( .A1(n89475), .A2(n89476), .ZN(n89468) );
  AOI22_X1 U75036 ( .A1(n105691), .A2(n109358), .B1(n105690), .B2(n109362), 
        .ZN(n89476) );
  AOI22_X1 U75037 ( .A1(n105689), .A2(n109356), .B1(n105688), .B2(n109361), 
        .ZN(n89475) );
  NAND2_X1 U75038 ( .A1(n89477), .A2(n89478), .ZN(n89467) );
  AOI22_X1 U75039 ( .A1(n86495), .A2(n72281), .B1(n105686), .B2(n109366), .ZN(
        n89478) );
  AOI22_X1 U75040 ( .A1(n105685), .A2(n72279), .B1(n105684), .B2(n109355), 
        .ZN(n89477) );
  NAND2_X1 U75041 ( .A1(n89479), .A2(n89480), .ZN(n89397) );
  NOR4_X1 U75042 ( .A1(n89481), .A2(n89482), .A3(n89483), .A4(n89484), .ZN(
        n89480) );
  NAND2_X1 U75043 ( .A1(n89485), .A2(n89486), .ZN(n89484) );
  AOI22_X1 U75044 ( .A1(n105683), .A2(n109395), .B1(n105682), .B2(n109394), 
        .ZN(n89486) );
  AOI22_X1 U75045 ( .A1(n105681), .A2(n72315), .B1(n105680), .B2(n109392), 
        .ZN(n89485) );
  NAND2_X1 U75046 ( .A1(n89487), .A2(n89488), .ZN(n89483) );
  AOI22_X1 U75047 ( .A1(n105679), .A2(n109390), .B1(n86514), .B2(n109393), 
        .ZN(n89488) );
  AOI22_X1 U75048 ( .A1(n86515), .A2(n72321), .B1(n105677), .B2(n109391), .ZN(
        n89487) );
  NAND2_X1 U75049 ( .A1(n89489), .A2(n89490), .ZN(n89482) );
  AOI22_X1 U75050 ( .A1(n86519), .A2(n109401), .B1(n86520), .B2(n72327), .ZN(
        n89490) );
  AOI22_X1 U75051 ( .A1(n86521), .A2(n109399), .B1(n86522), .B2(n109400), .ZN(
        n89489) );
  NAND2_X1 U75052 ( .A1(n89491), .A2(n89492), .ZN(n89481) );
  AOI22_X1 U75053 ( .A1(n105676), .A2(n109396), .B1(n86526), .B2(n109398), 
        .ZN(n89492) );
  AOI22_X1 U75054 ( .A1(n86527), .A2(n109402), .B1(n86528), .B2(n109397), .ZN(
        n89491) );
  NOR4_X1 U75055 ( .A1(n89493), .A2(n89494), .A3(n89495), .A4(n89496), .ZN(
        n89479) );
  NAND2_X1 U75056 ( .A1(n89497), .A2(n89498), .ZN(n89496) );
  AOI22_X1 U75057 ( .A1(n86535), .A2(n109376), .B1(n105674), .B2(n109380), 
        .ZN(n89498) );
  AOI22_X1 U75058 ( .A1(n105673), .A2(n109379), .B1(n105672), .B2(n72298), 
        .ZN(n89497) );
  NAND2_X1 U75059 ( .A1(n89499), .A2(n89500), .ZN(n89495) );
  AOI22_X1 U75060 ( .A1(n105671), .A2(n109386), .B1(n105670), .B2(n109375), 
        .ZN(n89500) );
  AOI22_X1 U75061 ( .A1(n105669), .A2(n109378), .B1(n86544), .B2(n109383), 
        .ZN(n89499) );
  NAND2_X1 U75062 ( .A1(n89501), .A2(n89502), .ZN(n89494) );
  AOI22_X1 U75063 ( .A1(n105667), .A2(n109382), .B1(n105666), .B2(n109387), 
        .ZN(n89502) );
  AOI22_X1 U75064 ( .A1(n105665), .A2(n109389), .B1(n105664), .B2(n109385), 
        .ZN(n89501) );
  NAND2_X1 U75065 ( .A1(n89503), .A2(n89504), .ZN(n89493) );
  AOI22_X1 U75066 ( .A1(n105663), .A2(n72316), .B1(n105662), .B2(n109381), 
        .ZN(n89504) );
  AOI22_X1 U75067 ( .A1(n86555), .A2(n109384), .B1(n105660), .B2(n109388), 
        .ZN(n89503) );
  AOI21_X1 U75068 ( .B1(n86302), .B2(n89506), .A(n89507), .ZN(n89505) );
  OAI21_X1 U75069 ( .B1(n89508), .B2(n105787), .A(n89509), .ZN(n89507) );
  OAI21_X1 U75070 ( .B1(n89510), .B2(n89511), .A(n86310), .ZN(n89509) );
  OAI21_X1 U75071 ( .B1(n109307), .B2(n105785), .A(n89512), .ZN(n89511) );
  AOI22_X1 U75072 ( .A1(n86313), .A2(n72204), .B1(n86314), .B2(n109305), .ZN(
        n89512) );
  NAND2_X1 U75073 ( .A1(n89513), .A2(n89514), .ZN(n89510) );
  AOI22_X1 U75074 ( .A1(n105783), .A2(n109303), .B1(n105782), .B2(n109308), 
        .ZN(n89514) );
  AOI22_X1 U75075 ( .A1(n105781), .A2(n109306), .B1(n105780), .B2(n109304), 
        .ZN(n89513) );
  NOR4_X1 U75076 ( .A1(n89515), .A2(n89516), .A3(n89517), .A4(n89518), .ZN(
        n89508) );
  NAND2_X1 U75077 ( .A1(n89519), .A2(n89520), .ZN(n89518) );
  NOR4_X1 U75078 ( .A1(n89521), .A2(n89522), .A3(n89523), .A4(n89524), .ZN(
        n89520) );
  NAND2_X1 U75079 ( .A1(n89525), .A2(n89526), .ZN(n89524) );
  AOI22_X1 U75080 ( .A1(n105779), .A2(n109284), .B1(n105778), .B2(n109285), 
        .ZN(n89526) );
  AOI22_X1 U75081 ( .A1(n105777), .A2(n109293), .B1(n105776), .B2(n109291), 
        .ZN(n89525) );
  NAND2_X1 U75082 ( .A1(n89527), .A2(n89528), .ZN(n89523) );
  AOI22_X1 U75083 ( .A1(n105775), .A2(n72073), .B1(n105774), .B2(n109288), 
        .ZN(n89528) );
  AOI22_X1 U75084 ( .A1(n105773), .A2(n72177), .B1(n105772), .B2(n109206), 
        .ZN(n89527) );
  NAND2_X1 U75085 ( .A1(n89529), .A2(n89530), .ZN(n89522) );
  AOI22_X1 U75086 ( .A1(n105771), .A2(n109210), .B1(n105770), .B2(n72077), 
        .ZN(n89530) );
  AOI22_X1 U75087 ( .A1(n105769), .A2(n109289), .B1(n105768), .B2(n109286), 
        .ZN(n89529) );
  NAND2_X1 U75088 ( .A1(n89531), .A2(n89532), .ZN(n89521) );
  AOI22_X1 U75089 ( .A1(n105767), .A2(n109208), .B1(n105766), .B2(n109212), 
        .ZN(n89532) );
  AOI22_X1 U75090 ( .A1(n105765), .A2(n109211), .B1(n105764), .B2(n72079), 
        .ZN(n89531) );
  NOR4_X1 U75091 ( .A1(n89533), .A2(n89534), .A3(n89535), .A4(n89536), .ZN(
        n89519) );
  NAND2_X1 U75092 ( .A1(n89537), .A2(n89538), .ZN(n89536) );
  AOI22_X1 U75093 ( .A1(n105763), .A2(n109294), .B1(n105762), .B2(n109297), 
        .ZN(n89538) );
  AOI22_X1 U75094 ( .A1(n105761), .A2(n109298), .B1(n86364), .B2(n109300), 
        .ZN(n89537) );
  NAND2_X1 U75095 ( .A1(n89539), .A2(n89540), .ZN(n89535) );
  AOI22_X1 U75096 ( .A1(n105759), .A2(n109299), .B1(n105758), .B2(n109295), 
        .ZN(n89540) );
  AOI22_X1 U75097 ( .A1(n105757), .A2(n109301), .B1(n105756), .B2(n109296), 
        .ZN(n89539) );
  NAND2_X1 U75098 ( .A1(n89541), .A2(n89542), .ZN(n89534) );
  AOI22_X1 U75099 ( .A1(n105755), .A2(n72187), .B1(n105754), .B2(n72186), .ZN(
        n89542) );
  AOI22_X1 U75100 ( .A1(n105753), .A2(n72189), .B1(n105752), .B2(n109302), 
        .ZN(n89541) );
  NAND2_X1 U75101 ( .A1(n89543), .A2(n89544), .ZN(n89533) );
  AOI22_X1 U75102 ( .A1(n105751), .A2(n109287), .B1(n105750), .B2(n109292), 
        .ZN(n89544) );
  AOI22_X1 U75103 ( .A1(n105749), .A2(n72184), .B1(n86382), .B2(n109290), .ZN(
        n89543) );
  NAND2_X1 U75104 ( .A1(n89545), .A2(n89546), .ZN(n89517) );
  NOR4_X1 U75105 ( .A1(n89547), .A2(n89548), .A3(n89549), .A4(n89550), .ZN(
        n89546) );
  NAND2_X1 U75106 ( .A1(n89551), .A2(n89552), .ZN(n89550) );
  AOI22_X1 U75107 ( .A1(n105747), .A2(n109221), .B1(n105746), .B2(n109223), 
        .ZN(n89552) );
  AOI22_X1 U75108 ( .A1(n105745), .A2(n72102), .B1(n105744), .B2(n109222), 
        .ZN(n89551) );
  NAND2_X1 U75109 ( .A1(n89553), .A2(n89554), .ZN(n89549) );
  AOI22_X1 U75110 ( .A1(n105743), .A2(n72106), .B1(n105742), .B2(n72108), .ZN(
        n89554) );
  AOI22_X1 U75111 ( .A1(n105741), .A2(n109229), .B1(n105740), .B2(n109230), 
        .ZN(n89553) );
  NAND2_X1 U75112 ( .A1(n89555), .A2(n89556), .ZN(n89548) );
  AOI22_X1 U75113 ( .A1(n105739), .A2(n109226), .B1(n105738), .B2(n109228), 
        .ZN(n89556) );
  AOI22_X1 U75114 ( .A1(n105737), .A2(n109231), .B1(n86406), .B2(n109227), 
        .ZN(n89555) );
  NAND2_X1 U75115 ( .A1(n89557), .A2(n89558), .ZN(n89547) );
  AOI22_X1 U75116 ( .A1(n105735), .A2(n109236), .B1(n105734), .B2(n72113), 
        .ZN(n89558) );
  AOI22_X1 U75117 ( .A1(n105733), .A2(n109235), .B1(n105732), .B2(n72111), 
        .ZN(n89557) );
  NOR4_X1 U75118 ( .A1(n89559), .A2(n89560), .A3(n89561), .A4(n89562), .ZN(
        n89545) );
  NAND2_X1 U75119 ( .A1(n89563), .A2(n89564), .ZN(n89562) );
  AOI22_X1 U75120 ( .A1(n105731), .A2(n109216), .B1(n105730), .B2(n109207), 
        .ZN(n89564) );
  AOI22_X1 U75121 ( .A1(n105729), .A2(n109209), .B1(n105728), .B2(n72085), 
        .ZN(n89563) );
  NAND2_X1 U75122 ( .A1(n89565), .A2(n89566), .ZN(n89561) );
  AOI22_X1 U75123 ( .A1(n105727), .A2(n109214), .B1(n105726), .B2(n109218), 
        .ZN(n89566) );
  AOI22_X1 U75124 ( .A1(n86427), .A2(n109220), .B1(n105724), .B2(n109217), 
        .ZN(n89565) );
  NAND2_X1 U75125 ( .A1(n89567), .A2(n89568), .ZN(n89560) );
  AOI22_X1 U75126 ( .A1(n105723), .A2(n72094), .B1(n105722), .B2(n109213), 
        .ZN(n89568) );
  AOI22_X1 U75127 ( .A1(n105721), .A2(n109215), .B1(n105720), .B2(n109219), 
        .ZN(n89567) );
  NAND2_X1 U75128 ( .A1(n89569), .A2(n89570), .ZN(n89559) );
  AOI22_X1 U75129 ( .A1(n105719), .A2(n109225), .B1(n105718), .B2(n72098), 
        .ZN(n89570) );
  AOI22_X1 U75130 ( .A1(n105717), .A2(n72096), .B1(n86440), .B2(n109224), .ZN(
        n89569) );
  NAND2_X1 U75131 ( .A1(n89571), .A2(n89572), .ZN(n89516) );
  NOR4_X1 U75132 ( .A1(n89573), .A2(n89574), .A3(n89575), .A4(n89576), .ZN(
        n89572) );
  NAND2_X1 U75133 ( .A1(n89577), .A2(n89578), .ZN(n89576) );
  AOI22_X1 U75134 ( .A1(n105715), .A2(n72136), .B1(n105714), .B2(n109246), 
        .ZN(n89578) );
  AOI22_X1 U75135 ( .A1(n105713), .A2(n109250), .B1(n105712), .B2(n109249), 
        .ZN(n89577) );
  NAND2_X1 U75136 ( .A1(n89579), .A2(n89580), .ZN(n89575) );
  AOI22_X1 U75137 ( .A1(n86455), .A2(n109255), .B1(n105710), .B2(n109254), 
        .ZN(n89580) );
  AOI22_X1 U75138 ( .A1(n86457), .A2(n109245), .B1(n105708), .B2(n109247), 
        .ZN(n89579) );
  NAND2_X1 U75139 ( .A1(n89581), .A2(n89582), .ZN(n89574) );
  AOI22_X1 U75140 ( .A1(n105707), .A2(n109256), .B1(n105706), .B2(n109252), 
        .ZN(n89582) );
  AOI22_X1 U75141 ( .A1(n105705), .A2(n72140), .B1(n105704), .B2(n72142), .ZN(
        n89581) );
  NAND2_X1 U75142 ( .A1(n89583), .A2(n89584), .ZN(n89573) );
  AOI22_X1 U75143 ( .A1(n105703), .A2(n109259), .B1(n105702), .B2(n72148), 
        .ZN(n89584) );
  AOI22_X1 U75144 ( .A1(n105701), .A2(n109251), .B1(n105700), .B2(n109253), 
        .ZN(n89583) );
  NOR4_X1 U75145 ( .A1(n89585), .A2(n89586), .A3(n89587), .A4(n89588), .ZN(
        n89571) );
  NAND2_X1 U75146 ( .A1(n89589), .A2(n89590), .ZN(n89588) );
  AOI22_X1 U75147 ( .A1(n105699), .A2(n109234), .B1(n105698), .B2(n109239), 
        .ZN(n89590) );
  AOI22_X1 U75148 ( .A1(n86479), .A2(n109233), .B1(n105696), .B2(n72116), .ZN(
        n89589) );
  NAND2_X1 U75149 ( .A1(n89591), .A2(n89592), .ZN(n89587) );
  AOI22_X1 U75150 ( .A1(n105695), .A2(n72125), .B1(n86484), .B2(n109241), .ZN(
        n89592) );
  AOI22_X1 U75151 ( .A1(n105693), .A2(n109242), .B1(n105692), .B2(n109232), 
        .ZN(n89591) );
  NAND2_X1 U75152 ( .A1(n89593), .A2(n89594), .ZN(n89586) );
  AOI22_X1 U75153 ( .A1(n105691), .A2(n109240), .B1(n105690), .B2(n109244), 
        .ZN(n89594) );
  AOI22_X1 U75154 ( .A1(n105689), .A2(n109238), .B1(n105688), .B2(n109243), 
        .ZN(n89593) );
  NAND2_X1 U75155 ( .A1(n89595), .A2(n89596), .ZN(n89585) );
  AOI22_X1 U75156 ( .A1(n86495), .A2(n72130), .B1(n105686), .B2(n109248), .ZN(
        n89596) );
  AOI22_X1 U75157 ( .A1(n105685), .A2(n72128), .B1(n105684), .B2(n109237), 
        .ZN(n89595) );
  NAND2_X1 U75158 ( .A1(n89597), .A2(n89598), .ZN(n89515) );
  NOR4_X1 U75159 ( .A1(n89599), .A2(n89600), .A3(n89601), .A4(n89602), .ZN(
        n89598) );
  NAND2_X1 U75160 ( .A1(n89603), .A2(n89604), .ZN(n89602) );
  AOI22_X1 U75161 ( .A1(n105683), .A2(n109277), .B1(n105682), .B2(n109276), 
        .ZN(n89604) );
  AOI22_X1 U75162 ( .A1(n105681), .A2(n72164), .B1(n105680), .B2(n109274), 
        .ZN(n89603) );
  NAND2_X1 U75163 ( .A1(n89605), .A2(n89606), .ZN(n89601) );
  AOI22_X1 U75164 ( .A1(n105679), .A2(n109272), .B1(n86514), .B2(n109275), 
        .ZN(n89606) );
  AOI22_X1 U75165 ( .A1(n86515), .A2(n72170), .B1(n105677), .B2(n109273), .ZN(
        n89605) );
  NAND2_X1 U75166 ( .A1(n89607), .A2(n89608), .ZN(n89600) );
  AOI22_X1 U75167 ( .A1(n86519), .A2(n109282), .B1(n86520), .B2(n72176), .ZN(
        n89608) );
  AOI22_X1 U75168 ( .A1(n86521), .A2(n109280), .B1(n86522), .B2(n109281), .ZN(
        n89607) );
  NAND2_X1 U75169 ( .A1(n89609), .A2(n89610), .ZN(n89599) );
  AOI22_X1 U75170 ( .A1(n105676), .A2(n109278), .B1(n86526), .B2(n72171), .ZN(
        n89610) );
  AOI22_X1 U75171 ( .A1(n86527), .A2(n109283), .B1(n86528), .B2(n109279), .ZN(
        n89609) );
  NOR4_X1 U75172 ( .A1(n89611), .A2(n89612), .A3(n89613), .A4(n89614), .ZN(
        n89597) );
  NAND2_X1 U75173 ( .A1(n89615), .A2(n89616), .ZN(n89614) );
  AOI22_X1 U75174 ( .A1(n86535), .A2(n109258), .B1(n105674), .B2(n109262), 
        .ZN(n89616) );
  AOI22_X1 U75175 ( .A1(n105673), .A2(n109261), .B1(n105672), .B2(n72147), 
        .ZN(n89615) );
  NAND2_X1 U75176 ( .A1(n89617), .A2(n89618), .ZN(n89613) );
  AOI22_X1 U75177 ( .A1(n105671), .A2(n109268), .B1(n105670), .B2(n109257), 
        .ZN(n89618) );
  AOI22_X1 U75178 ( .A1(n105669), .A2(n109260), .B1(n86544), .B2(n109265), 
        .ZN(n89617) );
  NAND2_X1 U75179 ( .A1(n89619), .A2(n89620), .ZN(n89612) );
  AOI22_X1 U75180 ( .A1(n105667), .A2(n109264), .B1(n105666), .B2(n109269), 
        .ZN(n89620) );
  AOI22_X1 U75181 ( .A1(n105665), .A2(n109271), .B1(n105664), .B2(n109267), 
        .ZN(n89619) );
  NAND2_X1 U75182 ( .A1(n89621), .A2(n89622), .ZN(n89611) );
  AOI22_X1 U75183 ( .A1(n105663), .A2(n72165), .B1(n105662), .B2(n109263), 
        .ZN(n89622) );
  AOI22_X1 U75184 ( .A1(n86555), .A2(n109266), .B1(n105660), .B2(n109270), 
        .ZN(n89621) );
  AOI21_X1 U75185 ( .B1(n86302), .B2(n89624), .A(n89625), .ZN(n89623) );
  OAI21_X1 U75186 ( .B1(n89626), .B2(n105787), .A(n89627), .ZN(n89625) );
  OAI21_X1 U75187 ( .B1(n89628), .B2(n89629), .A(n86310), .ZN(n89627) );
  OAI21_X1 U75188 ( .B1(n109199), .B2(n105785), .A(n89630), .ZN(n89629) );
  AOI22_X1 U75189 ( .A1(n86313), .A2(n72060), .B1(n86314), .B2(n109197), .ZN(
        n89630) );
  NAND2_X1 U75190 ( .A1(n89631), .A2(n89632), .ZN(n89628) );
  AOI22_X1 U75191 ( .A1(n105783), .A2(n109195), .B1(n105782), .B2(n109200), 
        .ZN(n89632) );
  AOI22_X1 U75192 ( .A1(n105781), .A2(n109198), .B1(n105780), .B2(n109196), 
        .ZN(n89631) );
  NOR4_X1 U75193 ( .A1(n89633), .A2(n89634), .A3(n89635), .A4(n89636), .ZN(
        n89626) );
  NAND2_X1 U75194 ( .A1(n89637), .A2(n89638), .ZN(n89636) );
  NOR4_X1 U75195 ( .A1(n89639), .A2(n89640), .A3(n89641), .A4(n89642), .ZN(
        n89638) );
  NAND2_X1 U75196 ( .A1(n89643), .A2(n89644), .ZN(n89642) );
  AOI22_X1 U75197 ( .A1(n105779), .A2(n109176), .B1(n105778), .B2(n109177), 
        .ZN(n89644) );
  AOI22_X1 U75198 ( .A1(n105777), .A2(n109185), .B1(n105776), .B2(n109183), 
        .ZN(n89643) );
  NAND2_X1 U75199 ( .A1(n89645), .A2(n89646), .ZN(n89641) );
  AOI22_X1 U75200 ( .A1(n105775), .A2(n71929), .B1(n105774), .B2(n109180), 
        .ZN(n89646) );
  AOI22_X1 U75201 ( .A1(n105773), .A2(n72033), .B1(n105772), .B2(n109098), 
        .ZN(n89645) );
  NAND2_X1 U75202 ( .A1(n89647), .A2(n89648), .ZN(n89640) );
  AOI22_X1 U75203 ( .A1(n105771), .A2(n109102), .B1(n105770), .B2(n71933), 
        .ZN(n89648) );
  AOI22_X1 U75204 ( .A1(n105769), .A2(n109181), .B1(n105768), .B2(n109178), 
        .ZN(n89647) );
  NAND2_X1 U75205 ( .A1(n89649), .A2(n89650), .ZN(n89639) );
  AOI22_X1 U75206 ( .A1(n105767), .A2(n109100), .B1(n105766), .B2(n109104), 
        .ZN(n89650) );
  AOI22_X1 U75207 ( .A1(n105765), .A2(n109103), .B1(n105764), .B2(n71935), 
        .ZN(n89649) );
  NOR4_X1 U75208 ( .A1(n89651), .A2(n89652), .A3(n89653), .A4(n89654), .ZN(
        n89637) );
  NAND2_X1 U75209 ( .A1(n89655), .A2(n89656), .ZN(n89654) );
  AOI22_X1 U75210 ( .A1(n105763), .A2(n109186), .B1(n105762), .B2(n109189), 
        .ZN(n89656) );
  AOI22_X1 U75211 ( .A1(n86363), .A2(n109190), .B1(n86364), .B2(n109192), .ZN(
        n89655) );
  NAND2_X1 U75212 ( .A1(n89657), .A2(n89658), .ZN(n89653) );
  AOI22_X1 U75213 ( .A1(n105759), .A2(n109191), .B1(n105758), .B2(n109187), 
        .ZN(n89658) );
  AOI22_X1 U75214 ( .A1(n105757), .A2(n109193), .B1(n105756), .B2(n109188), 
        .ZN(n89657) );
  NAND2_X1 U75215 ( .A1(n89659), .A2(n89660), .ZN(n89652) );
  AOI22_X1 U75216 ( .A1(n105755), .A2(n72043), .B1(n105754), .B2(n72042), .ZN(
        n89660) );
  AOI22_X1 U75217 ( .A1(n105753), .A2(n72045), .B1(n105752), .B2(n109194), 
        .ZN(n89659) );
  NAND2_X1 U75218 ( .A1(n89661), .A2(n89662), .ZN(n89651) );
  AOI22_X1 U75219 ( .A1(n105751), .A2(n109179), .B1(n105750), .B2(n109184), 
        .ZN(n89662) );
  AOI22_X1 U75220 ( .A1(n105749), .A2(n72040), .B1(n86382), .B2(n109182), .ZN(
        n89661) );
  NAND2_X1 U75221 ( .A1(n89663), .A2(n89664), .ZN(n89635) );
  NOR4_X1 U75222 ( .A1(n89665), .A2(n89666), .A3(n89667), .A4(n89668), .ZN(
        n89664) );
  NAND2_X1 U75223 ( .A1(n89669), .A2(n89670), .ZN(n89668) );
  AOI22_X1 U75224 ( .A1(n105747), .A2(n109113), .B1(n105746), .B2(n109115), 
        .ZN(n89670) );
  AOI22_X1 U75225 ( .A1(n105745), .A2(n71958), .B1(n105744), .B2(n109114), 
        .ZN(n89669) );
  NAND2_X1 U75226 ( .A1(n89671), .A2(n89672), .ZN(n89667) );
  AOI22_X1 U75227 ( .A1(n105743), .A2(n71962), .B1(n105742), .B2(n71964), .ZN(
        n89672) );
  AOI22_X1 U75228 ( .A1(n105741), .A2(n109121), .B1(n105740), .B2(n109122), 
        .ZN(n89671) );
  NAND2_X1 U75229 ( .A1(n89673), .A2(n89674), .ZN(n89666) );
  AOI22_X1 U75230 ( .A1(n105739), .A2(n109118), .B1(n105738), .B2(n109120), 
        .ZN(n89674) );
  AOI22_X1 U75231 ( .A1(n105737), .A2(n109123), .B1(n86406), .B2(n109119), 
        .ZN(n89673) );
  NAND2_X1 U75232 ( .A1(n89675), .A2(n89676), .ZN(n89665) );
  AOI22_X1 U75233 ( .A1(n105735), .A2(n109128), .B1(n105734), .B2(n71969), 
        .ZN(n89676) );
  AOI22_X1 U75234 ( .A1(n105733), .A2(n109127), .B1(n105732), .B2(n71967), 
        .ZN(n89675) );
  NOR4_X1 U75235 ( .A1(n89677), .A2(n89678), .A3(n89679), .A4(n89680), .ZN(
        n89663) );
  NAND2_X1 U75236 ( .A1(n89681), .A2(n89682), .ZN(n89680) );
  AOI22_X1 U75237 ( .A1(n105731), .A2(n109108), .B1(n105730), .B2(n109099), 
        .ZN(n89682) );
  AOI22_X1 U75238 ( .A1(n105729), .A2(n109101), .B1(n105728), .B2(n71941), 
        .ZN(n89681) );
  NAND2_X1 U75239 ( .A1(n89683), .A2(n89684), .ZN(n89679) );
  AOI22_X1 U75240 ( .A1(n105727), .A2(n109106), .B1(n105726), .B2(n109110), 
        .ZN(n89684) );
  AOI22_X1 U75241 ( .A1(n86427), .A2(n109112), .B1(n105724), .B2(n109109), 
        .ZN(n89683) );
  NAND2_X1 U75242 ( .A1(n89685), .A2(n89686), .ZN(n89678) );
  AOI22_X1 U75243 ( .A1(n105723), .A2(n71950), .B1(n105722), .B2(n109105), 
        .ZN(n89686) );
  AOI22_X1 U75244 ( .A1(n105721), .A2(n109107), .B1(n105720), .B2(n109111), 
        .ZN(n89685) );
  NAND2_X1 U75245 ( .A1(n89687), .A2(n89688), .ZN(n89677) );
  AOI22_X1 U75246 ( .A1(n105719), .A2(n109117), .B1(n105718), .B2(n71954), 
        .ZN(n89688) );
  AOI22_X1 U75247 ( .A1(n105717), .A2(n71952), .B1(n86440), .B2(n109116), .ZN(
        n89687) );
  NAND2_X1 U75248 ( .A1(n89689), .A2(n89690), .ZN(n89634) );
  NOR4_X1 U75249 ( .A1(n89691), .A2(n89692), .A3(n89693), .A4(n89694), .ZN(
        n89690) );
  NAND2_X1 U75250 ( .A1(n89695), .A2(n89696), .ZN(n89694) );
  AOI22_X1 U75251 ( .A1(n105715), .A2(n71992), .B1(n105714), .B2(n109138), 
        .ZN(n89696) );
  AOI22_X1 U75252 ( .A1(n105713), .A2(n109142), .B1(n105712), .B2(n109141), 
        .ZN(n89695) );
  NAND2_X1 U75253 ( .A1(n89697), .A2(n89698), .ZN(n89693) );
  AOI22_X1 U75254 ( .A1(n86455), .A2(n109147), .B1(n105710), .B2(n109146), 
        .ZN(n89698) );
  AOI22_X1 U75255 ( .A1(n86457), .A2(n109137), .B1(n105708), .B2(n109139), 
        .ZN(n89697) );
  NAND2_X1 U75256 ( .A1(n89699), .A2(n89700), .ZN(n89692) );
  AOI22_X1 U75257 ( .A1(n105707), .A2(n71997), .B1(n105706), .B2(n109144), 
        .ZN(n89700) );
  AOI22_X1 U75258 ( .A1(n105705), .A2(n71996), .B1(n105704), .B2(n71998), .ZN(
        n89699) );
  NAND2_X1 U75259 ( .A1(n89701), .A2(n89702), .ZN(n89691) );
  AOI22_X1 U75260 ( .A1(n105703), .A2(n109150), .B1(n105702), .B2(n72004), 
        .ZN(n89702) );
  AOI22_X1 U75261 ( .A1(n105701), .A2(n109143), .B1(n105700), .B2(n109145), 
        .ZN(n89701) );
  NOR4_X1 U75262 ( .A1(n89703), .A2(n89704), .A3(n89705), .A4(n89706), .ZN(
        n89689) );
  NAND2_X1 U75263 ( .A1(n89707), .A2(n89708), .ZN(n89706) );
  AOI22_X1 U75264 ( .A1(n105699), .A2(n109126), .B1(n105698), .B2(n109131), 
        .ZN(n89708) );
  AOI22_X1 U75265 ( .A1(n86479), .A2(n109125), .B1(n105696), .B2(n71972), .ZN(
        n89707) );
  NAND2_X1 U75266 ( .A1(n89709), .A2(n89710), .ZN(n89705) );
  AOI22_X1 U75267 ( .A1(n105695), .A2(n71981), .B1(n105694), .B2(n109133), 
        .ZN(n89710) );
  AOI22_X1 U75268 ( .A1(n105693), .A2(n109134), .B1(n105692), .B2(n109124), 
        .ZN(n89709) );
  NAND2_X1 U75269 ( .A1(n89711), .A2(n89712), .ZN(n89704) );
  AOI22_X1 U75270 ( .A1(n105691), .A2(n109132), .B1(n105690), .B2(n109136), 
        .ZN(n89712) );
  AOI22_X1 U75271 ( .A1(n105689), .A2(n109130), .B1(n105688), .B2(n109135), 
        .ZN(n89711) );
  NAND2_X1 U75272 ( .A1(n89713), .A2(n89714), .ZN(n89703) );
  AOI22_X1 U75273 ( .A1(n86495), .A2(n71986), .B1(n105686), .B2(n109140), .ZN(
        n89714) );
  AOI22_X1 U75274 ( .A1(n105685), .A2(n71984), .B1(n105684), .B2(n109129), 
        .ZN(n89713) );
  NAND2_X1 U75275 ( .A1(n89715), .A2(n89716), .ZN(n89633) );
  NOR4_X1 U75276 ( .A1(n89717), .A2(n89718), .A3(n89719), .A4(n89720), .ZN(
        n89716) );
  NAND2_X1 U75277 ( .A1(n89721), .A2(n89722), .ZN(n89720) );
  AOI22_X1 U75278 ( .A1(n105683), .A2(n109168), .B1(n105682), .B2(n109167), 
        .ZN(n89722) );
  AOI22_X1 U75279 ( .A1(n105681), .A2(n72020), .B1(n105680), .B2(n109165), 
        .ZN(n89721) );
  NAND2_X1 U75280 ( .A1(n89723), .A2(n89724), .ZN(n89719) );
  AOI22_X1 U75281 ( .A1(n105679), .A2(n109163), .B1(n86514), .B2(n109166), 
        .ZN(n89724) );
  AOI22_X1 U75282 ( .A1(n86515), .A2(n72026), .B1(n105677), .B2(n109164), .ZN(
        n89723) );
  NAND2_X1 U75283 ( .A1(n89725), .A2(n89726), .ZN(n89718) );
  AOI22_X1 U75284 ( .A1(n86519), .A2(n109174), .B1(n86520), .B2(n72032), .ZN(
        n89726) );
  AOI22_X1 U75285 ( .A1(n86521), .A2(n109172), .B1(n86522), .B2(n109173), .ZN(
        n89725) );
  NAND2_X1 U75286 ( .A1(n89727), .A2(n89728), .ZN(n89717) );
  AOI22_X1 U75287 ( .A1(n105676), .A2(n109169), .B1(n86526), .B2(n109171), 
        .ZN(n89728) );
  AOI22_X1 U75288 ( .A1(n86527), .A2(n109175), .B1(n86528), .B2(n109170), .ZN(
        n89727) );
  NOR4_X1 U75289 ( .A1(n89729), .A2(n89730), .A3(n89731), .A4(n89732), .ZN(
        n89715) );
  NAND2_X1 U75290 ( .A1(n89733), .A2(n89734), .ZN(n89732) );
  AOI22_X1 U75291 ( .A1(n86535), .A2(n109149), .B1(n105674), .B2(n109153), 
        .ZN(n89734) );
  AOI22_X1 U75292 ( .A1(n105673), .A2(n109152), .B1(n105672), .B2(n72003), 
        .ZN(n89733) );
  NAND2_X1 U75293 ( .A1(n89735), .A2(n89736), .ZN(n89731) );
  AOI22_X1 U75294 ( .A1(n105671), .A2(n109159), .B1(n105670), .B2(n109148), 
        .ZN(n89736) );
  AOI22_X1 U75295 ( .A1(n105669), .A2(n109151), .B1(n86544), .B2(n109156), 
        .ZN(n89735) );
  NAND2_X1 U75296 ( .A1(n89737), .A2(n89738), .ZN(n89730) );
  AOI22_X1 U75297 ( .A1(n105667), .A2(n109155), .B1(n105666), .B2(n109160), 
        .ZN(n89738) );
  AOI22_X1 U75298 ( .A1(n105665), .A2(n109162), .B1(n105664), .B2(n109158), 
        .ZN(n89737) );
  NAND2_X1 U75299 ( .A1(n89739), .A2(n89740), .ZN(n89729) );
  AOI22_X1 U75300 ( .A1(n105663), .A2(n72021), .B1(n105662), .B2(n109154), 
        .ZN(n89740) );
  AOI22_X1 U75301 ( .A1(n86555), .A2(n109157), .B1(n105660), .B2(n109161), 
        .ZN(n89739) );
  AOI21_X1 U75302 ( .B1(n86302), .B2(n89742), .A(n89743), .ZN(n89741) );
  OAI21_X1 U75303 ( .B1(n89744), .B2(n105787), .A(n89745), .ZN(n89743) );
  OAI21_X1 U75304 ( .B1(n89746), .B2(n89747), .A(n86310), .ZN(n89745) );
  OAI21_X1 U75305 ( .B1(n108734), .B2(n105785), .A(n89748), .ZN(n89747) );
  AOI22_X1 U75306 ( .A1(n86313), .A2(n71462), .B1(n86314), .B2(n108732), .ZN(
        n89748) );
  NAND2_X1 U75307 ( .A1(n89749), .A2(n89750), .ZN(n89746) );
  AOI22_X1 U75308 ( .A1(n105783), .A2(n108730), .B1(n105782), .B2(n108735), 
        .ZN(n89750) );
  AOI22_X1 U75309 ( .A1(n105781), .A2(n108733), .B1(n105780), .B2(n108731), 
        .ZN(n89749) );
  NOR4_X1 U75310 ( .A1(n89751), .A2(n89752), .A3(n89753), .A4(n89754), .ZN(
        n89744) );
  NAND2_X1 U75311 ( .A1(n89755), .A2(n89756), .ZN(n89754) );
  NOR4_X1 U75312 ( .A1(n89757), .A2(n89758), .A3(n89759), .A4(n89760), .ZN(
        n89756) );
  NAND2_X1 U75313 ( .A1(n89761), .A2(n89762), .ZN(n89760) );
  AOI22_X1 U75314 ( .A1(n105779), .A2(n108711), .B1(n105778), .B2(n108712), 
        .ZN(n89762) );
  AOI22_X1 U75315 ( .A1(n105777), .A2(n108720), .B1(n105776), .B2(n108718), 
        .ZN(n89761) );
  NAND2_X1 U75316 ( .A1(n89763), .A2(n89764), .ZN(n89759) );
  AOI22_X1 U75317 ( .A1(n105775), .A2(n71331), .B1(n105774), .B2(n108715), 
        .ZN(n89764) );
  AOI22_X1 U75318 ( .A1(n105773), .A2(n71435), .B1(n105772), .B2(n108633), 
        .ZN(n89763) );
  NAND2_X1 U75319 ( .A1(n89765), .A2(n89766), .ZN(n89758) );
  AOI22_X1 U75320 ( .A1(n105771), .A2(n108637), .B1(n105770), .B2(n71335), 
        .ZN(n89766) );
  AOI22_X1 U75321 ( .A1(n105769), .A2(n108716), .B1(n105768), .B2(n108713), 
        .ZN(n89765) );
  NAND2_X1 U75322 ( .A1(n89767), .A2(n89768), .ZN(n89757) );
  AOI22_X1 U75323 ( .A1(n105767), .A2(n108635), .B1(n105766), .B2(n108639), 
        .ZN(n89768) );
  AOI22_X1 U75324 ( .A1(n105765), .A2(n108638), .B1(n105764), .B2(n71337), 
        .ZN(n89767) );
  NOR4_X1 U75325 ( .A1(n89769), .A2(n89770), .A3(n89771), .A4(n89772), .ZN(
        n89755) );
  NAND2_X1 U75326 ( .A1(n89773), .A2(n89774), .ZN(n89772) );
  AOI22_X1 U75327 ( .A1(n105763), .A2(n108721), .B1(n105762), .B2(n108724), 
        .ZN(n89774) );
  AOI22_X1 U75328 ( .A1(n105761), .A2(n108725), .B1(n86364), .B2(n108727), 
        .ZN(n89773) );
  NAND2_X1 U75329 ( .A1(n89775), .A2(n89776), .ZN(n89771) );
  AOI22_X1 U75330 ( .A1(n105759), .A2(n108726), .B1(n105758), .B2(n108722), 
        .ZN(n89776) );
  AOI22_X1 U75331 ( .A1(n105757), .A2(n108728), .B1(n105756), .B2(n108723), 
        .ZN(n89775) );
  NAND2_X1 U75332 ( .A1(n89777), .A2(n89778), .ZN(n89770) );
  AOI22_X1 U75333 ( .A1(n105755), .A2(n71445), .B1(n105754), .B2(n71444), .ZN(
        n89778) );
  AOI22_X1 U75334 ( .A1(n105753), .A2(n71447), .B1(n105752), .B2(n108729), 
        .ZN(n89777) );
  NAND2_X1 U75335 ( .A1(n89779), .A2(n89780), .ZN(n89769) );
  AOI22_X1 U75336 ( .A1(n105751), .A2(n108714), .B1(n105750), .B2(n108719), 
        .ZN(n89780) );
  AOI22_X1 U75337 ( .A1(n105749), .A2(n71442), .B1(n86382), .B2(n108717), .ZN(
        n89779) );
  NAND2_X1 U75338 ( .A1(n89781), .A2(n89782), .ZN(n89753) );
  NOR4_X1 U75339 ( .A1(n89783), .A2(n89784), .A3(n89785), .A4(n89786), .ZN(
        n89782) );
  NAND2_X1 U75340 ( .A1(n89787), .A2(n89788), .ZN(n89786) );
  AOI22_X1 U75341 ( .A1(n105747), .A2(n108648), .B1(n105746), .B2(n108650), 
        .ZN(n89788) );
  AOI22_X1 U75342 ( .A1(n105745), .A2(n71360), .B1(n105744), .B2(n108649), 
        .ZN(n89787) );
  NAND2_X1 U75343 ( .A1(n89789), .A2(n89790), .ZN(n89785) );
  AOI22_X1 U75344 ( .A1(n105743), .A2(n71364), .B1(n105742), .B2(n71366), .ZN(
        n89790) );
  AOI22_X1 U75345 ( .A1(n105741), .A2(n108656), .B1(n105740), .B2(n108657), 
        .ZN(n89789) );
  NAND2_X1 U75346 ( .A1(n89791), .A2(n89792), .ZN(n89784) );
  AOI22_X1 U75347 ( .A1(n105739), .A2(n108653), .B1(n105738), .B2(n108655), 
        .ZN(n89792) );
  AOI22_X1 U75348 ( .A1(n105737), .A2(n108658), .B1(n86406), .B2(n108654), 
        .ZN(n89791) );
  NAND2_X1 U75349 ( .A1(n89793), .A2(n89794), .ZN(n89783) );
  AOI22_X1 U75350 ( .A1(n105735), .A2(n108663), .B1(n105734), .B2(n71371), 
        .ZN(n89794) );
  AOI22_X1 U75351 ( .A1(n105733), .A2(n108662), .B1(n105732), .B2(n71369), 
        .ZN(n89793) );
  NOR4_X1 U75352 ( .A1(n89795), .A2(n89796), .A3(n89797), .A4(n89798), .ZN(
        n89781) );
  NAND2_X1 U75353 ( .A1(n89799), .A2(n89800), .ZN(n89798) );
  AOI22_X1 U75354 ( .A1(n105731), .A2(n108643), .B1(n105730), .B2(n108634), 
        .ZN(n89800) );
  AOI22_X1 U75355 ( .A1(n105729), .A2(n108636), .B1(n105728), .B2(n71343), 
        .ZN(n89799) );
  NAND2_X1 U75356 ( .A1(n89801), .A2(n89802), .ZN(n89797) );
  AOI22_X1 U75357 ( .A1(n105727), .A2(n108641), .B1(n105726), .B2(n108645), 
        .ZN(n89802) );
  AOI22_X1 U75358 ( .A1(n86427), .A2(n108647), .B1(n105724), .B2(n108644), 
        .ZN(n89801) );
  NAND2_X1 U75359 ( .A1(n89803), .A2(n89804), .ZN(n89796) );
  AOI22_X1 U75360 ( .A1(n105723), .A2(n71352), .B1(n105722), .B2(n108640), 
        .ZN(n89804) );
  AOI22_X1 U75361 ( .A1(n105721), .A2(n108642), .B1(n105720), .B2(n108646), 
        .ZN(n89803) );
  NAND2_X1 U75362 ( .A1(n89805), .A2(n89806), .ZN(n89795) );
  AOI22_X1 U75363 ( .A1(n105719), .A2(n108652), .B1(n105718), .B2(n71356), 
        .ZN(n89806) );
  AOI22_X1 U75364 ( .A1(n105717), .A2(n71354), .B1(n86440), .B2(n108651), .ZN(
        n89805) );
  NAND2_X1 U75365 ( .A1(n89807), .A2(n89808), .ZN(n89752) );
  NOR4_X1 U75366 ( .A1(n89809), .A2(n89810), .A3(n89811), .A4(n89812), .ZN(
        n89808) );
  NAND2_X1 U75367 ( .A1(n89813), .A2(n89814), .ZN(n89812) );
  AOI22_X1 U75368 ( .A1(n105715), .A2(n71394), .B1(n105714), .B2(n108673), 
        .ZN(n89814) );
  AOI22_X1 U75369 ( .A1(n105713), .A2(n108677), .B1(n105712), .B2(n108676), 
        .ZN(n89813) );
  NAND2_X1 U75370 ( .A1(n89815), .A2(n89816), .ZN(n89811) );
  AOI22_X1 U75371 ( .A1(n86455), .A2(n108682), .B1(n105710), .B2(n108681), 
        .ZN(n89816) );
  AOI22_X1 U75372 ( .A1(n86457), .A2(n108672), .B1(n105708), .B2(n108674), 
        .ZN(n89815) );
  NAND2_X1 U75373 ( .A1(n89817), .A2(n89818), .ZN(n89810) );
  AOI22_X1 U75374 ( .A1(n105707), .A2(n108683), .B1(n105706), .B2(n108679), 
        .ZN(n89818) );
  AOI22_X1 U75375 ( .A1(n105705), .A2(n71398), .B1(n105704), .B2(n71400), .ZN(
        n89817) );
  NAND2_X1 U75376 ( .A1(n89819), .A2(n89820), .ZN(n89809) );
  AOI22_X1 U75377 ( .A1(n105703), .A2(n108686), .B1(n105702), .B2(n71406), 
        .ZN(n89820) );
  AOI22_X1 U75378 ( .A1(n105701), .A2(n108678), .B1(n105700), .B2(n108680), 
        .ZN(n89819) );
  NOR4_X1 U75379 ( .A1(n89821), .A2(n89822), .A3(n89823), .A4(n89824), .ZN(
        n89807) );
  NAND2_X1 U75380 ( .A1(n89825), .A2(n89826), .ZN(n89824) );
  AOI22_X1 U75381 ( .A1(n105699), .A2(n108661), .B1(n105698), .B2(n108666), 
        .ZN(n89826) );
  AOI22_X1 U75382 ( .A1(n86479), .A2(n108660), .B1(n105696), .B2(n71374), .ZN(
        n89825) );
  NAND2_X1 U75383 ( .A1(n89827), .A2(n89828), .ZN(n89823) );
  AOI22_X1 U75384 ( .A1(n105695), .A2(n71383), .B1(n86484), .B2(n108668), .ZN(
        n89828) );
  AOI22_X1 U75385 ( .A1(n105693), .A2(n108669), .B1(n105692), .B2(n108659), 
        .ZN(n89827) );
  NAND2_X1 U75386 ( .A1(n89829), .A2(n89830), .ZN(n89822) );
  AOI22_X1 U75387 ( .A1(n105691), .A2(n108667), .B1(n105690), .B2(n108671), 
        .ZN(n89830) );
  AOI22_X1 U75388 ( .A1(n105689), .A2(n108665), .B1(n105688), .B2(n108670), 
        .ZN(n89829) );
  NAND2_X1 U75389 ( .A1(n89831), .A2(n89832), .ZN(n89821) );
  AOI22_X1 U75390 ( .A1(n86495), .A2(n71388), .B1(n105686), .B2(n108675), .ZN(
        n89832) );
  AOI22_X1 U75391 ( .A1(n105685), .A2(n71386), .B1(n105684), .B2(n108664), 
        .ZN(n89831) );
  NAND2_X1 U75392 ( .A1(n89833), .A2(n89834), .ZN(n89751) );
  NOR4_X1 U75393 ( .A1(n89835), .A2(n89836), .A3(n89837), .A4(n89838), .ZN(
        n89834) );
  NAND2_X1 U75394 ( .A1(n89839), .A2(n89840), .ZN(n89838) );
  AOI22_X1 U75395 ( .A1(n105683), .A2(n108704), .B1(n105682), .B2(n108703), 
        .ZN(n89840) );
  AOI22_X1 U75396 ( .A1(n105681), .A2(n71422), .B1(n105680), .B2(n108701), 
        .ZN(n89839) );
  NAND2_X1 U75397 ( .A1(n89841), .A2(n89842), .ZN(n89837) );
  AOI22_X1 U75398 ( .A1(n105679), .A2(n108699), .B1(n86514), .B2(n108702), 
        .ZN(n89842) );
  AOI22_X1 U75399 ( .A1(n86515), .A2(n71428), .B1(n105677), .B2(n108700), .ZN(
        n89841) );
  NAND2_X1 U75400 ( .A1(n89843), .A2(n89844), .ZN(n89836) );
  AOI22_X1 U75401 ( .A1(n86519), .A2(n108709), .B1(n86520), .B2(n71434), .ZN(
        n89844) );
  AOI22_X1 U75402 ( .A1(n86521), .A2(n108707), .B1(n86522), .B2(n108708), .ZN(
        n89843) );
  NAND2_X1 U75403 ( .A1(n89845), .A2(n89846), .ZN(n89835) );
  AOI22_X1 U75404 ( .A1(n105676), .A2(n108705), .B1(n86526), .B2(n71429), .ZN(
        n89846) );
  AOI22_X1 U75405 ( .A1(n86527), .A2(n108710), .B1(n86528), .B2(n108706), .ZN(
        n89845) );
  NOR4_X1 U75406 ( .A1(n89847), .A2(n89848), .A3(n89849), .A4(n89850), .ZN(
        n89833) );
  NAND2_X1 U75407 ( .A1(n89851), .A2(n89852), .ZN(n89850) );
  AOI22_X1 U75408 ( .A1(n86535), .A2(n108685), .B1(n105674), .B2(n108689), 
        .ZN(n89852) );
  AOI22_X1 U75409 ( .A1(n105673), .A2(n108688), .B1(n105672), .B2(n71405), 
        .ZN(n89851) );
  NAND2_X1 U75410 ( .A1(n89853), .A2(n89854), .ZN(n89849) );
  AOI22_X1 U75411 ( .A1(n105671), .A2(n108695), .B1(n105670), .B2(n108684), 
        .ZN(n89854) );
  AOI22_X1 U75412 ( .A1(n105669), .A2(n108687), .B1(n86544), .B2(n108692), 
        .ZN(n89853) );
  NAND2_X1 U75413 ( .A1(n89855), .A2(n89856), .ZN(n89848) );
  AOI22_X1 U75414 ( .A1(n105667), .A2(n108691), .B1(n105666), .B2(n108696), 
        .ZN(n89856) );
  AOI22_X1 U75415 ( .A1(n105665), .A2(n108698), .B1(n105664), .B2(n108694), 
        .ZN(n89855) );
  NAND2_X1 U75416 ( .A1(n89857), .A2(n89858), .ZN(n89847) );
  AOI22_X1 U75417 ( .A1(n105663), .A2(n71423), .B1(n105662), .B2(n108690), 
        .ZN(n89858) );
  AOI22_X1 U75418 ( .A1(n86555), .A2(n108693), .B1(n105660), .B2(n108697), 
        .ZN(n89857) );
  AOI21_X1 U75419 ( .B1(n86302), .B2(n81790), .A(n89860), .ZN(n89859) );
  OAI21_X1 U75420 ( .B1(n89861), .B2(n105787), .A(n89862), .ZN(n89860) );
  OAI21_X1 U75421 ( .B1(n89863), .B2(n89864), .A(n86310), .ZN(n89862) );
  OAI21_X1 U75422 ( .B1(n108962), .B2(n105785), .A(n89865), .ZN(n89864) );
  AOI22_X1 U75423 ( .A1(n86313), .A2(n71757), .B1(n86314), .B2(n108960), .ZN(
        n89865) );
  NAND2_X1 U75424 ( .A1(n89866), .A2(n89867), .ZN(n89863) );
  AOI22_X1 U75425 ( .A1(n105783), .A2(n108958), .B1(n105782), .B2(n108963), 
        .ZN(n89867) );
  AOI22_X1 U75426 ( .A1(n105781), .A2(n108961), .B1(n105780), .B2(n108959), 
        .ZN(n89866) );
  NOR4_X1 U75427 ( .A1(n89868), .A2(n89869), .A3(n89870), .A4(n89871), .ZN(
        n89861) );
  NAND2_X1 U75428 ( .A1(n89872), .A2(n89873), .ZN(n89871) );
  NOR4_X1 U75429 ( .A1(n89874), .A2(n89875), .A3(n89876), .A4(n89877), .ZN(
        n89873) );
  NAND2_X1 U75430 ( .A1(n89878), .A2(n89879), .ZN(n89877) );
  AOI22_X1 U75431 ( .A1(n105779), .A2(n108939), .B1(n105778), .B2(n108940), 
        .ZN(n89879) );
  AOI22_X1 U75432 ( .A1(n105777), .A2(n108948), .B1(n105776), .B2(n108946), 
        .ZN(n89878) );
  NAND2_X1 U75433 ( .A1(n89880), .A2(n89881), .ZN(n89876) );
  AOI22_X1 U75434 ( .A1(n105775), .A2(n71626), .B1(n105774), .B2(n108943), 
        .ZN(n89881) );
  AOI22_X1 U75435 ( .A1(n105773), .A2(n71730), .B1(n105772), .B2(n108860), 
        .ZN(n89880) );
  NAND2_X1 U75436 ( .A1(n89882), .A2(n89883), .ZN(n89875) );
  AOI22_X1 U75437 ( .A1(n105771), .A2(n108864), .B1(n105770), .B2(n71630), 
        .ZN(n89883) );
  AOI22_X1 U75438 ( .A1(n105769), .A2(n108944), .B1(n105768), .B2(n108941), 
        .ZN(n89882) );
  NAND2_X1 U75439 ( .A1(n89884), .A2(n89885), .ZN(n89874) );
  AOI22_X1 U75440 ( .A1(n105767), .A2(n108862), .B1(n105766), .B2(n108866), 
        .ZN(n89885) );
  AOI22_X1 U75441 ( .A1(n105765), .A2(n108865), .B1(n105764), .B2(n71632), 
        .ZN(n89884) );
  NOR4_X1 U75442 ( .A1(n89886), .A2(n89887), .A3(n89888), .A4(n89889), .ZN(
        n89872) );
  NAND2_X1 U75443 ( .A1(n89890), .A2(n89891), .ZN(n89889) );
  AOI22_X1 U75444 ( .A1(n105763), .A2(n108949), .B1(n105762), .B2(n108952), 
        .ZN(n89891) );
  AOI22_X1 U75445 ( .A1(n86363), .A2(n108953), .B1(n86364), .B2(n108955), .ZN(
        n89890) );
  NAND2_X1 U75446 ( .A1(n89892), .A2(n89893), .ZN(n89888) );
  AOI22_X1 U75447 ( .A1(n105759), .A2(n108954), .B1(n105758), .B2(n108950), 
        .ZN(n89893) );
  AOI22_X1 U75448 ( .A1(n105757), .A2(n108956), .B1(n105756), .B2(n108951), 
        .ZN(n89892) );
  NAND2_X1 U75449 ( .A1(n89894), .A2(n89895), .ZN(n89887) );
  AOI22_X1 U75450 ( .A1(n105755), .A2(n71740), .B1(n105754), .B2(n71739), .ZN(
        n89895) );
  AOI22_X1 U75451 ( .A1(n105753), .A2(n71742), .B1(n105752), .B2(n108957), 
        .ZN(n89894) );
  NAND2_X1 U75452 ( .A1(n89896), .A2(n89897), .ZN(n89886) );
  AOI22_X1 U75453 ( .A1(n105751), .A2(n108942), .B1(n105750), .B2(n108947), 
        .ZN(n89897) );
  AOI22_X1 U75454 ( .A1(n105749), .A2(n71737), .B1(n86382), .B2(n108945), .ZN(
        n89896) );
  NAND2_X1 U75455 ( .A1(n89898), .A2(n89899), .ZN(n89870) );
  NOR4_X1 U75456 ( .A1(n89900), .A2(n89901), .A3(n89902), .A4(n89903), .ZN(
        n89899) );
  NAND2_X1 U75457 ( .A1(n89904), .A2(n89905), .ZN(n89903) );
  AOI22_X1 U75458 ( .A1(n105747), .A2(n108875), .B1(n105746), .B2(n108877), 
        .ZN(n89905) );
  AOI22_X1 U75459 ( .A1(n105745), .A2(n71655), .B1(n105744), .B2(n108876), 
        .ZN(n89904) );
  NAND2_X1 U75460 ( .A1(n89906), .A2(n89907), .ZN(n89902) );
  AOI22_X1 U75461 ( .A1(n105743), .A2(n71659), .B1(n105742), .B2(n71661), .ZN(
        n89907) );
  AOI22_X1 U75462 ( .A1(n105741), .A2(n108883), .B1(n105740), .B2(n108884), 
        .ZN(n89906) );
  NAND2_X1 U75463 ( .A1(n89908), .A2(n89909), .ZN(n89901) );
  AOI22_X1 U75464 ( .A1(n105739), .A2(n108880), .B1(n105738), .B2(n108882), 
        .ZN(n89909) );
  AOI22_X1 U75465 ( .A1(n105737), .A2(n108885), .B1(n86406), .B2(n108881), 
        .ZN(n89908) );
  NAND2_X1 U75466 ( .A1(n89910), .A2(n89911), .ZN(n89900) );
  AOI22_X1 U75467 ( .A1(n105735), .A2(n108890), .B1(n105734), .B2(n71666), 
        .ZN(n89911) );
  AOI22_X1 U75468 ( .A1(n105733), .A2(n108889), .B1(n105732), .B2(n71664), 
        .ZN(n89910) );
  NOR4_X1 U75469 ( .A1(n89912), .A2(n89913), .A3(n89914), .A4(n89915), .ZN(
        n89898) );
  NAND2_X1 U75470 ( .A1(n89916), .A2(n89917), .ZN(n89915) );
  AOI22_X1 U75471 ( .A1(n105731), .A2(n108870), .B1(n105730), .B2(n108861), 
        .ZN(n89917) );
  AOI22_X1 U75472 ( .A1(n105729), .A2(n108863), .B1(n105728), .B2(n71638), 
        .ZN(n89916) );
  NAND2_X1 U75473 ( .A1(n89918), .A2(n89919), .ZN(n89914) );
  AOI22_X1 U75474 ( .A1(n105727), .A2(n108868), .B1(n105726), .B2(n108872), 
        .ZN(n89919) );
  AOI22_X1 U75475 ( .A1(n86427), .A2(n108874), .B1(n105724), .B2(n108871), 
        .ZN(n89918) );
  NAND2_X1 U75476 ( .A1(n89920), .A2(n89921), .ZN(n89913) );
  AOI22_X1 U75477 ( .A1(n105723), .A2(n71647), .B1(n105722), .B2(n108867), 
        .ZN(n89921) );
  AOI22_X1 U75478 ( .A1(n105721), .A2(n108869), .B1(n105720), .B2(n108873), 
        .ZN(n89920) );
  NAND2_X1 U75479 ( .A1(n89922), .A2(n89923), .ZN(n89912) );
  AOI22_X1 U75480 ( .A1(n105719), .A2(n108879), .B1(n105718), .B2(n71651), 
        .ZN(n89923) );
  AOI22_X1 U75481 ( .A1(n105717), .A2(n71649), .B1(n86440), .B2(n108878), .ZN(
        n89922) );
  NAND2_X1 U75482 ( .A1(n89924), .A2(n89925), .ZN(n89869) );
  NOR4_X1 U75483 ( .A1(n89926), .A2(n89927), .A3(n89928), .A4(n89929), .ZN(
        n89925) );
  NAND2_X1 U75484 ( .A1(n89930), .A2(n89931), .ZN(n89929) );
  AOI22_X1 U75485 ( .A1(n105715), .A2(n71689), .B1(n105714), .B2(n108900), 
        .ZN(n89931) );
  AOI22_X1 U75486 ( .A1(n105713), .A2(n108904), .B1(n105712), .B2(n108903), 
        .ZN(n89930) );
  NAND2_X1 U75487 ( .A1(n89932), .A2(n89933), .ZN(n89928) );
  AOI22_X1 U75488 ( .A1(n86455), .A2(n108909), .B1(n105710), .B2(n108908), 
        .ZN(n89933) );
  AOI22_X1 U75489 ( .A1(n86457), .A2(n108899), .B1(n105708), .B2(n108901), 
        .ZN(n89932) );
  NAND2_X1 U75490 ( .A1(n89934), .A2(n89935), .ZN(n89927) );
  AOI22_X1 U75491 ( .A1(n105707), .A2(n108910), .B1(n105706), .B2(n108906), 
        .ZN(n89935) );
  AOI22_X1 U75492 ( .A1(n105705), .A2(n71693), .B1(n105704), .B2(n71695), .ZN(
        n89934) );
  NAND2_X1 U75493 ( .A1(n89936), .A2(n89937), .ZN(n89926) );
  AOI22_X1 U75494 ( .A1(n105703), .A2(n108913), .B1(n105702), .B2(n71701), 
        .ZN(n89937) );
  AOI22_X1 U75495 ( .A1(n105701), .A2(n108905), .B1(n105700), .B2(n108907), 
        .ZN(n89936) );
  NOR4_X1 U75496 ( .A1(n89938), .A2(n89939), .A3(n89940), .A4(n89941), .ZN(
        n89924) );
  NAND2_X1 U75497 ( .A1(n89942), .A2(n89943), .ZN(n89941) );
  AOI22_X1 U75498 ( .A1(n105699), .A2(n108888), .B1(n105698), .B2(n108893), 
        .ZN(n89943) );
  AOI22_X1 U75499 ( .A1(n86479), .A2(n108887), .B1(n105696), .B2(n71669), .ZN(
        n89942) );
  NAND2_X1 U75500 ( .A1(n89944), .A2(n89945), .ZN(n89940) );
  AOI22_X1 U75501 ( .A1(n105695), .A2(n71678), .B1(n105694), .B2(n108895), 
        .ZN(n89945) );
  AOI22_X1 U75502 ( .A1(n105693), .A2(n108896), .B1(n105692), .B2(n108886), 
        .ZN(n89944) );
  NAND2_X1 U75503 ( .A1(n89946), .A2(n89947), .ZN(n89939) );
  AOI22_X1 U75504 ( .A1(n105691), .A2(n108894), .B1(n105690), .B2(n108898), 
        .ZN(n89947) );
  AOI22_X1 U75505 ( .A1(n105689), .A2(n108892), .B1(n105688), .B2(n108897), 
        .ZN(n89946) );
  NAND2_X1 U75506 ( .A1(n89948), .A2(n89949), .ZN(n89938) );
  AOI22_X1 U75507 ( .A1(n86495), .A2(n71683), .B1(n105686), .B2(n108902), .ZN(
        n89949) );
  AOI22_X1 U75508 ( .A1(n105685), .A2(n71681), .B1(n105684), .B2(n108891), 
        .ZN(n89948) );
  NAND2_X1 U75509 ( .A1(n89950), .A2(n89951), .ZN(n89868) );
  NOR4_X1 U75510 ( .A1(n89952), .A2(n89953), .A3(n89954), .A4(n89955), .ZN(
        n89951) );
  NAND2_X1 U75511 ( .A1(n89956), .A2(n89957), .ZN(n89955) );
  AOI22_X1 U75512 ( .A1(n105683), .A2(n108931), .B1(n105682), .B2(n108930), 
        .ZN(n89957) );
  AOI22_X1 U75513 ( .A1(n105681), .A2(n71717), .B1(n105680), .B2(n108928), 
        .ZN(n89956) );
  NAND2_X1 U75514 ( .A1(n89958), .A2(n89959), .ZN(n89954) );
  AOI22_X1 U75515 ( .A1(n105679), .A2(n108926), .B1(n86514), .B2(n108929), 
        .ZN(n89959) );
  AOI22_X1 U75516 ( .A1(n86515), .A2(n71723), .B1(n105677), .B2(n108927), .ZN(
        n89958) );
  NAND2_X1 U75517 ( .A1(n89960), .A2(n89961), .ZN(n89953) );
  AOI22_X1 U75518 ( .A1(n86519), .A2(n108937), .B1(n86520), .B2(n71729), .ZN(
        n89961) );
  AOI22_X1 U75519 ( .A1(n86521), .A2(n108935), .B1(n86522), .B2(n108936), .ZN(
        n89960) );
  NAND2_X1 U75520 ( .A1(n89962), .A2(n89963), .ZN(n89952) );
  AOI22_X1 U75521 ( .A1(n105676), .A2(n108932), .B1(n86526), .B2(n108934), 
        .ZN(n89963) );
  AOI22_X1 U75522 ( .A1(n86527), .A2(n108938), .B1(n86528), .B2(n108933), .ZN(
        n89962) );
  NOR4_X1 U75523 ( .A1(n89964), .A2(n89965), .A3(n89966), .A4(n89967), .ZN(
        n89950) );
  NAND2_X1 U75524 ( .A1(n89968), .A2(n89969), .ZN(n89967) );
  AOI22_X1 U75525 ( .A1(n86535), .A2(n108912), .B1(n105674), .B2(n108916), 
        .ZN(n89969) );
  AOI22_X1 U75526 ( .A1(n105673), .A2(n108915), .B1(n105672), .B2(n71700), 
        .ZN(n89968) );
  NAND2_X1 U75527 ( .A1(n89970), .A2(n89971), .ZN(n89966) );
  AOI22_X1 U75528 ( .A1(n105671), .A2(n108922), .B1(n105670), .B2(n108911), 
        .ZN(n89971) );
  AOI22_X1 U75529 ( .A1(n105669), .A2(n108914), .B1(n86544), .B2(n108919), 
        .ZN(n89970) );
  NAND2_X1 U75530 ( .A1(n89972), .A2(n89973), .ZN(n89965) );
  AOI22_X1 U75531 ( .A1(n105667), .A2(n108918), .B1(n105666), .B2(n108923), 
        .ZN(n89973) );
  AOI22_X1 U75532 ( .A1(n105665), .A2(n108925), .B1(n105664), .B2(n108921), 
        .ZN(n89972) );
  NAND2_X1 U75533 ( .A1(n89974), .A2(n89975), .ZN(n89964) );
  AOI22_X1 U75534 ( .A1(n105663), .A2(n71718), .B1(n105662), .B2(n108917), 
        .ZN(n89975) );
  AOI22_X1 U75535 ( .A1(n86555), .A2(n108920), .B1(n105660), .B2(n108924), 
        .ZN(n89974) );
  AOI21_X1 U75536 ( .B1(n86302), .B2(n89977), .A(n89978), .ZN(n89976) );
  OAI21_X1 U75537 ( .B1(n89979), .B2(n105787), .A(n89980), .ZN(n89978) );
  OAI21_X1 U75538 ( .B1(n89981), .B2(n89982), .A(n86310), .ZN(n89980) );
  OAI21_X1 U75539 ( .B1(n108850), .B2(n105785), .A(n89983), .ZN(n89982) );
  AOI22_X1 U75540 ( .A1(n86313), .A2(n71613), .B1(n86314), .B2(n108848), .ZN(
        n89983) );
  NAND2_X1 U75541 ( .A1(n89984), .A2(n89985), .ZN(n89981) );
  AOI22_X1 U75542 ( .A1(n105783), .A2(n108846), .B1(n105782), .B2(n108851), 
        .ZN(n89985) );
  AOI22_X1 U75543 ( .A1(n105781), .A2(n108849), .B1(n105780), .B2(n108847), 
        .ZN(n89984) );
  NOR4_X1 U75544 ( .A1(n89986), .A2(n89987), .A3(n89988), .A4(n89989), .ZN(
        n89979) );
  NAND2_X1 U75545 ( .A1(n89990), .A2(n89991), .ZN(n89989) );
  NOR4_X1 U75546 ( .A1(n89992), .A2(n89993), .A3(n89994), .A4(n89995), .ZN(
        n89991) );
  NAND2_X1 U75547 ( .A1(n89996), .A2(n89997), .ZN(n89995) );
  AOI22_X1 U75548 ( .A1(n105779), .A2(n108827), .B1(n105778), .B2(n108828), 
        .ZN(n89997) );
  AOI22_X1 U75549 ( .A1(n105777), .A2(n108836), .B1(n105776), .B2(n108834), 
        .ZN(n89996) );
  NAND2_X1 U75550 ( .A1(n89998), .A2(n89999), .ZN(n89994) );
  AOI22_X1 U75551 ( .A1(n105775), .A2(n71482), .B1(n105774), .B2(n108831), 
        .ZN(n89999) );
  AOI22_X1 U75552 ( .A1(n105773), .A2(n71586), .B1(n105772), .B2(n108748), 
        .ZN(n89998) );
  NAND2_X1 U75553 ( .A1(n90000), .A2(n90001), .ZN(n89993) );
  AOI22_X1 U75554 ( .A1(n105771), .A2(n108752), .B1(n105770), .B2(n71486), 
        .ZN(n90001) );
  AOI22_X1 U75555 ( .A1(n105769), .A2(n108832), .B1(n105768), .B2(n108829), 
        .ZN(n90000) );
  NAND2_X1 U75556 ( .A1(n90002), .A2(n90003), .ZN(n89992) );
  AOI22_X1 U75557 ( .A1(n105767), .A2(n108750), .B1(n105766), .B2(n108754), 
        .ZN(n90003) );
  AOI22_X1 U75558 ( .A1(n105765), .A2(n108753), .B1(n105764), .B2(n71488), 
        .ZN(n90002) );
  NOR4_X1 U75559 ( .A1(n90004), .A2(n90005), .A3(n90006), .A4(n90007), .ZN(
        n89990) );
  NAND2_X1 U75560 ( .A1(n90008), .A2(n90009), .ZN(n90007) );
  AOI22_X1 U75561 ( .A1(n105763), .A2(n108837), .B1(n105762), .B2(n108840), 
        .ZN(n90009) );
  AOI22_X1 U75562 ( .A1(n105761), .A2(n108841), .B1(n86364), .B2(n108843), 
        .ZN(n90008) );
  NAND2_X1 U75563 ( .A1(n90010), .A2(n90011), .ZN(n90006) );
  AOI22_X1 U75564 ( .A1(n105759), .A2(n108842), .B1(n105758), .B2(n108838), 
        .ZN(n90011) );
  AOI22_X1 U75565 ( .A1(n105757), .A2(n108844), .B1(n105756), .B2(n108839), 
        .ZN(n90010) );
  NAND2_X1 U75566 ( .A1(n90012), .A2(n90013), .ZN(n90005) );
  AOI22_X1 U75567 ( .A1(n105755), .A2(n71596), .B1(n105754), .B2(n71595), .ZN(
        n90013) );
  AOI22_X1 U75568 ( .A1(n105753), .A2(n71598), .B1(n105752), .B2(n108845), 
        .ZN(n90012) );
  NAND2_X1 U75569 ( .A1(n90014), .A2(n90015), .ZN(n90004) );
  AOI22_X1 U75570 ( .A1(n105751), .A2(n108830), .B1(n105750), .B2(n108835), 
        .ZN(n90015) );
  AOI22_X1 U75571 ( .A1(n105749), .A2(n71593), .B1(n86382), .B2(n108833), .ZN(
        n90014) );
  NAND2_X1 U75572 ( .A1(n90016), .A2(n90017), .ZN(n89988) );
  NOR4_X1 U75573 ( .A1(n90018), .A2(n90019), .A3(n90020), .A4(n90021), .ZN(
        n90017) );
  NAND2_X1 U75574 ( .A1(n90022), .A2(n90023), .ZN(n90021) );
  AOI22_X1 U75575 ( .A1(n105747), .A2(n108763), .B1(n105746), .B2(n108765), 
        .ZN(n90023) );
  AOI22_X1 U75576 ( .A1(n105745), .A2(n71511), .B1(n105744), .B2(n108764), 
        .ZN(n90022) );
  NAND2_X1 U75577 ( .A1(n90024), .A2(n90025), .ZN(n90020) );
  AOI22_X1 U75578 ( .A1(n105743), .A2(n71515), .B1(n105742), .B2(n71517), .ZN(
        n90025) );
  AOI22_X1 U75579 ( .A1(n105741), .A2(n108771), .B1(n105740), .B2(n108772), 
        .ZN(n90024) );
  NAND2_X1 U75580 ( .A1(n90026), .A2(n90027), .ZN(n90019) );
  AOI22_X1 U75581 ( .A1(n105739), .A2(n108768), .B1(n105738), .B2(n108770), 
        .ZN(n90027) );
  AOI22_X1 U75582 ( .A1(n105737), .A2(n108773), .B1(n86406), .B2(n108769), 
        .ZN(n90026) );
  NAND2_X1 U75583 ( .A1(n90028), .A2(n90029), .ZN(n90018) );
  AOI22_X1 U75584 ( .A1(n105735), .A2(n108778), .B1(n105734), .B2(n71522), 
        .ZN(n90029) );
  AOI22_X1 U75585 ( .A1(n105733), .A2(n108777), .B1(n105732), .B2(n71520), 
        .ZN(n90028) );
  NOR4_X1 U75586 ( .A1(n90030), .A2(n90031), .A3(n90032), .A4(n90033), .ZN(
        n90016) );
  NAND2_X1 U75587 ( .A1(n90034), .A2(n90035), .ZN(n90033) );
  AOI22_X1 U75588 ( .A1(n105731), .A2(n108758), .B1(n105730), .B2(n108749), 
        .ZN(n90035) );
  AOI22_X1 U75589 ( .A1(n105729), .A2(n108751), .B1(n105728), .B2(n71494), 
        .ZN(n90034) );
  NAND2_X1 U75590 ( .A1(n90036), .A2(n90037), .ZN(n90032) );
  AOI22_X1 U75591 ( .A1(n105727), .A2(n108756), .B1(n105726), .B2(n108760), 
        .ZN(n90037) );
  AOI22_X1 U75592 ( .A1(n86427), .A2(n108762), .B1(n105724), .B2(n108759), 
        .ZN(n90036) );
  NAND2_X1 U75593 ( .A1(n90038), .A2(n90039), .ZN(n90031) );
  AOI22_X1 U75594 ( .A1(n105723), .A2(n71503), .B1(n105722), .B2(n108755), 
        .ZN(n90039) );
  AOI22_X1 U75595 ( .A1(n105721), .A2(n108757), .B1(n105720), .B2(n108761), 
        .ZN(n90038) );
  NAND2_X1 U75596 ( .A1(n90040), .A2(n90041), .ZN(n90030) );
  AOI22_X1 U75597 ( .A1(n105719), .A2(n108767), .B1(n105718), .B2(n71507), 
        .ZN(n90041) );
  AOI22_X1 U75598 ( .A1(n105717), .A2(n71505), .B1(n86440), .B2(n108766), .ZN(
        n90040) );
  NAND2_X1 U75599 ( .A1(n90042), .A2(n90043), .ZN(n89987) );
  NOR4_X1 U75600 ( .A1(n90044), .A2(n90045), .A3(n90046), .A4(n90047), .ZN(
        n90043) );
  NAND2_X1 U75601 ( .A1(n90048), .A2(n90049), .ZN(n90047) );
  AOI22_X1 U75602 ( .A1(n105715), .A2(n71545), .B1(n105714), .B2(n108788), 
        .ZN(n90049) );
  AOI22_X1 U75603 ( .A1(n105713), .A2(n108792), .B1(n105712), .B2(n108791), 
        .ZN(n90048) );
  NAND2_X1 U75604 ( .A1(n90050), .A2(n90051), .ZN(n90046) );
  AOI22_X1 U75605 ( .A1(n86455), .A2(n108797), .B1(n105710), .B2(n108796), 
        .ZN(n90051) );
  AOI22_X1 U75606 ( .A1(n86457), .A2(n108787), .B1(n105708), .B2(n108789), 
        .ZN(n90050) );
  NAND2_X1 U75607 ( .A1(n90052), .A2(n90053), .ZN(n90045) );
  AOI22_X1 U75608 ( .A1(n105707), .A2(n108798), .B1(n105706), .B2(n108794), 
        .ZN(n90053) );
  AOI22_X1 U75609 ( .A1(n105705), .A2(n71549), .B1(n105704), .B2(n71551), .ZN(
        n90052) );
  NAND2_X1 U75610 ( .A1(n90054), .A2(n90055), .ZN(n90044) );
  AOI22_X1 U75611 ( .A1(n105703), .A2(n108801), .B1(n105702), .B2(n71557), 
        .ZN(n90055) );
  AOI22_X1 U75612 ( .A1(n105701), .A2(n108793), .B1(n105700), .B2(n108795), 
        .ZN(n90054) );
  NOR4_X1 U75613 ( .A1(n90056), .A2(n90057), .A3(n90058), .A4(n90059), .ZN(
        n90042) );
  NAND2_X1 U75614 ( .A1(n90060), .A2(n90061), .ZN(n90059) );
  AOI22_X1 U75615 ( .A1(n105699), .A2(n108776), .B1(n105698), .B2(n108781), 
        .ZN(n90061) );
  AOI22_X1 U75616 ( .A1(n86479), .A2(n108775), .B1(n105696), .B2(n71525), .ZN(
        n90060) );
  NAND2_X1 U75617 ( .A1(n90062), .A2(n90063), .ZN(n90058) );
  AOI22_X1 U75618 ( .A1(n105695), .A2(n71534), .B1(n86484), .B2(n108783), .ZN(
        n90063) );
  AOI22_X1 U75619 ( .A1(n105693), .A2(n108784), .B1(n105692), .B2(n108774), 
        .ZN(n90062) );
  NAND2_X1 U75620 ( .A1(n90064), .A2(n90065), .ZN(n90057) );
  AOI22_X1 U75621 ( .A1(n105691), .A2(n108782), .B1(n105690), .B2(n108786), 
        .ZN(n90065) );
  AOI22_X1 U75622 ( .A1(n105689), .A2(n108780), .B1(n105688), .B2(n108785), 
        .ZN(n90064) );
  NAND2_X1 U75623 ( .A1(n90066), .A2(n90067), .ZN(n90056) );
  AOI22_X1 U75624 ( .A1(n86495), .A2(n71539), .B1(n105686), .B2(n108790), .ZN(
        n90067) );
  AOI22_X1 U75625 ( .A1(n105685), .A2(n71537), .B1(n105684), .B2(n108779), 
        .ZN(n90066) );
  NAND2_X1 U75626 ( .A1(n90068), .A2(n90069), .ZN(n89986) );
  NOR4_X1 U75627 ( .A1(n90070), .A2(n90071), .A3(n90072), .A4(n90073), .ZN(
        n90069) );
  NAND2_X1 U75628 ( .A1(n90074), .A2(n90075), .ZN(n90073) );
  AOI22_X1 U75629 ( .A1(n105683), .A2(n108819), .B1(n105682), .B2(n108818), 
        .ZN(n90075) );
  AOI22_X1 U75630 ( .A1(n105681), .A2(n71573), .B1(n105680), .B2(n108816), 
        .ZN(n90074) );
  NAND2_X1 U75631 ( .A1(n90076), .A2(n90077), .ZN(n90072) );
  AOI22_X1 U75632 ( .A1(n105679), .A2(n108814), .B1(n86514), .B2(n108817), 
        .ZN(n90077) );
  AOI22_X1 U75633 ( .A1(n86515), .A2(n71579), .B1(n105677), .B2(n108815), .ZN(
        n90076) );
  NAND2_X1 U75634 ( .A1(n90078), .A2(n90079), .ZN(n90071) );
  AOI22_X1 U75635 ( .A1(n86519), .A2(n108825), .B1(n86520), .B2(n71585), .ZN(
        n90079) );
  AOI22_X1 U75636 ( .A1(n86521), .A2(n108823), .B1(n86522), .B2(n108824), .ZN(
        n90078) );
  NAND2_X1 U75637 ( .A1(n90080), .A2(n90081), .ZN(n90070) );
  AOI22_X1 U75638 ( .A1(n105676), .A2(n108820), .B1(n86526), .B2(n108822), 
        .ZN(n90081) );
  AOI22_X1 U75639 ( .A1(n86527), .A2(n108826), .B1(n86528), .B2(n108821), .ZN(
        n90080) );
  NOR4_X1 U75640 ( .A1(n90082), .A2(n90083), .A3(n90084), .A4(n90085), .ZN(
        n90068) );
  NAND2_X1 U75641 ( .A1(n90086), .A2(n90087), .ZN(n90085) );
  AOI22_X1 U75642 ( .A1(n86535), .A2(n108800), .B1(n105674), .B2(n108804), 
        .ZN(n90087) );
  AOI22_X1 U75643 ( .A1(n105673), .A2(n108803), .B1(n105672), .B2(n71556), 
        .ZN(n90086) );
  NAND2_X1 U75644 ( .A1(n90088), .A2(n90089), .ZN(n90084) );
  AOI22_X1 U75645 ( .A1(n105671), .A2(n108810), .B1(n105670), .B2(n108799), 
        .ZN(n90089) );
  AOI22_X1 U75646 ( .A1(n105669), .A2(n108802), .B1(n86544), .B2(n108807), 
        .ZN(n90088) );
  NAND2_X1 U75647 ( .A1(n90090), .A2(n90091), .ZN(n90083) );
  AOI22_X1 U75648 ( .A1(n105667), .A2(n108806), .B1(n105666), .B2(n108811), 
        .ZN(n90091) );
  AOI22_X1 U75649 ( .A1(n105665), .A2(n108813), .B1(n105664), .B2(n108809), 
        .ZN(n90090) );
  NAND2_X1 U75650 ( .A1(n90092), .A2(n90093), .ZN(n90082) );
  AOI22_X1 U75651 ( .A1(n105663), .A2(n71574), .B1(n105662), .B2(n108805), 
        .ZN(n90093) );
  AOI22_X1 U75652 ( .A1(n86555), .A2(n108808), .B1(n105660), .B2(n108812), 
        .ZN(n90092) );
  OAI21_X1 U75653 ( .B1(n90094), .B2(n105787), .A(n90095), .ZN(
        \DLX_Datapath/RegisterFile/N46866 ) );
  AOI22_X1 U75654 ( .A1(n86302), .A2(n90096), .B1(n86310), .B2(n90097), .ZN(
        n90095) );
  OR2_X1 U75655 ( .A1(n90098), .A2(n90099), .ZN(n90097) );
  OAI21_X1 U75656 ( .B1(n107167), .B2(n105785), .A(n90100), .ZN(n90099) );
  AOI22_X1 U75657 ( .A1(n86313), .A2(n69430), .B1(n86314), .B2(n107171), .ZN(
        n90100) );
  NOR2_X1 U75658 ( .A1(n90101), .A2(n59442), .ZN(n86314) );
  AND2_X2 U75659 ( .A1(n90102), .A2(n107137), .ZN(n86313) );
  OR2_X1 U75660 ( .A1(n90103), .A2(n107136), .ZN(n86311) );
  NAND2_X1 U75661 ( .A1(n90104), .A2(n90105), .ZN(n90098) );
  AOI22_X1 U75662 ( .A1(n105783), .A2(n107175), .B1(n105782), .B2(n106767), 
        .ZN(n90105) );
  NOR2_X1 U75663 ( .A1(n107136), .A2(n90101), .ZN(n86318) );
  OR2_X1 U75664 ( .A1(n90106), .A2(n107134), .ZN(n90101) );
  NOR2_X1 U75665 ( .A1(n90107), .A2(n59442), .ZN(n86317) );
  AOI22_X1 U75666 ( .A1(n105781), .A2(n107169), .B1(n105780), .B2(n107173), 
        .ZN(n90104) );
  NOR2_X1 U75667 ( .A1(n90103), .A2(n59442), .ZN(n86320) );
  NAND2_X1 U75668 ( .A1(n59435), .A2(n107134), .ZN(n90103) );
  NOR2_X1 U75669 ( .A1(n107136), .A2(n90107), .ZN(n86319) );
  OR2_X1 U75670 ( .A1(n90106), .A2(n59441), .ZN(n90107) );
  AOI21_X1 U75671 ( .B1(n69424), .B2(n90109), .A(n90110), .ZN(n86310) );
  AND2_X2 U75672 ( .A1(n90111), .A2(n90112), .ZN(n86302) );
  AOI22_X1 U75673 ( .A1(n90102), .A2(n90108), .B1(n107140), .B2(n107120), .ZN(
        n90112) );
  NOR4_X1 U75674 ( .A1(n90113), .A2(n90114), .A3(n107121), .A4(n107124), .ZN(
        n90109) );
  NOR3_X1 U75675 ( .A1(n90116), .A2(n107131), .A3(n107125), .ZN(n90115) );
  AOI22_X1 U75676 ( .A1(n90119), .A2(n107134), .B1(n90120), .B2(n107132), .ZN(
        n90118) );
  NOR2_X1 U75677 ( .A1(n107142), .A2(n107137), .ZN(n90108) );
  NOR2_X1 U75678 ( .A1(n90121), .A2(n107134), .ZN(n90102) );
  AOI21_X1 U75679 ( .B1(n90122), .B2(n90110), .A(n111056), .ZN(n90111) );
  OAI21_X1 U75680 ( .B1(n111056), .B2(n90122), .A(n90110), .ZN(n86306) );
  NAND2_X1 U75681 ( .A1(n90123), .A2(n90124), .ZN(n90122) );
  NOR4_X1 U75682 ( .A1(n90125), .A2(n90126), .A3(n90114), .A4(n90113), .ZN(
        n90124) );
  NOR2_X1 U75683 ( .A1(n90120), .A2(n107132), .ZN(n90113) );
  NOR2_X1 U75684 ( .A1(n90119), .A2(n107134), .ZN(n90114) );
  NOR2_X1 U75685 ( .A1(n59441), .A2(n107122), .ZN(n90126) );
  OAI21_X1 U75686 ( .B1(n59435), .B2(n107114), .A(n90117), .ZN(n90125) );
  XNOR2_X1 U75687 ( .A(n90127), .B(n59442), .ZN(n90117) );
  NOR4_X1 U75688 ( .A1(n90128), .A2(n90129), .A3(n90130), .A4(n90131), .ZN(
        n90123) );
  XNOR2_X1 U75689 ( .A(\DLX_Datapath/RegisterFile/N46177 ), .B(n90132), .ZN(
        n90131) );
  XNOR2_X1 U75690 ( .A(n90133), .B(n90134), .ZN(n90130) );
  XOR2_X1 U75691 ( .A(\DLX_Datapath/RegisterFile/N46178 ), .B(n90135), .Z(
        n90129) );
  OR2_X1 U75692 ( .A1(n90136), .A2(n90116), .ZN(n90128) );
  XOR2_X1 U75693 ( .A(n104762), .B(n107139), .Z(n90116) );
  NOR4_X1 U75694 ( .A1(n90138), .A2(n90139), .A3(n90140), .A4(n90141), .ZN(
        n90094) );
  NAND2_X1 U75695 ( .A1(n90142), .A2(n90143), .ZN(n90141) );
  NOR4_X1 U75696 ( .A1(n90144), .A2(n90145), .A3(n90146), .A4(n90147), .ZN(
        n90143) );
  NAND2_X1 U75697 ( .A1(n90148), .A2(n90149), .ZN(n90147) );
  AOI22_X1 U75698 ( .A1(n105779), .A2(n107213), .B1(n105778), .B2(n107211), 
        .ZN(n90149) );
  NOR2_X1 U75699 ( .A1(n90150), .A2(n90151), .ZN(n86334) );
  NOR2_X1 U75700 ( .A1(n90152), .A2(n90153), .ZN(n86333) );
  AOI22_X1 U75701 ( .A1(n105777), .A2(n107195), .B1(n105776), .B2(n107199), 
        .ZN(n90148) );
  NOR2_X1 U75702 ( .A1(n90150), .A2(n90154), .ZN(n86336) );
  NOR2_X1 U75703 ( .A1(n90155), .A2(n90156), .ZN(n86335) );
  NAND2_X1 U75704 ( .A1(n90157), .A2(n90158), .ZN(n90146) );
  AOI22_X1 U75705 ( .A1(n105775), .A2(n69591), .B1(n105774), .B2(n107205), 
        .ZN(n90158) );
  NOR2_X1 U75706 ( .A1(n90159), .A2(n90153), .ZN(n86340) );
  NOR2_X1 U75707 ( .A1(n90160), .A2(n90161), .ZN(n86339) );
  AOI22_X1 U75708 ( .A1(n105773), .A2(n69484), .B1(n105772), .B2(n107288), 
        .ZN(n90157) );
  NOR2_X1 U75709 ( .A1(n90160), .A2(n90162), .ZN(n86342) );
  NOR2_X1 U75710 ( .A1(n90152), .A2(n90151), .ZN(n86341) );
  NAND2_X1 U75711 ( .A1(n90163), .A2(n90164), .ZN(n90145) );
  AOI22_X1 U75712 ( .A1(n105771), .A2(n107292), .B1(n105770), .B2(n69595), 
        .ZN(n90164) );
  NOR2_X1 U75713 ( .A1(n90165), .A2(n90161), .ZN(n86346) );
  NOR2_X1 U75714 ( .A1(n90166), .A2(n90162), .ZN(n86345) );
  AOI22_X1 U75715 ( .A1(n105769), .A2(n107203), .B1(n105768), .B2(n107209), 
        .ZN(n90163) );
  NOR2_X1 U75716 ( .A1(n90150), .A2(n90153), .ZN(n86348) );
  NOR2_X1 U75717 ( .A1(n90155), .A2(n90151), .ZN(n86347) );
  NAND2_X1 U75718 ( .A1(n90167), .A2(n90168), .ZN(n90144) );
  AOI22_X1 U75719 ( .A1(n105767), .A2(n107290), .B1(n105766), .B2(n107294), 
        .ZN(n90168) );
  NOR2_X1 U75720 ( .A1(n90160), .A2(n90169), .ZN(n86352) );
  NOR2_X1 U75721 ( .A1(n90170), .A2(n90162), .ZN(n86351) );
  AOI22_X1 U75722 ( .A1(n105765), .A2(n107293), .B1(n105764), .B2(n69597), 
        .ZN(n90167) );
  NOR2_X1 U75723 ( .A1(n90166), .A2(n90161), .ZN(n86354) );
  NOR2_X1 U75724 ( .A1(n90160), .A2(n90171), .ZN(n86353) );
  NOR4_X1 U75725 ( .A1(n90172), .A2(n90173), .A3(n90174), .A4(n90175), .ZN(
        n90142) );
  NAND2_X1 U75726 ( .A1(n90176), .A2(n90177), .ZN(n90175) );
  AOI22_X1 U75727 ( .A1(n105763), .A2(n107193), .B1(n105762), .B2(n107187), 
        .ZN(n90177) );
  NOR2_X1 U75728 ( .A1(n90150), .A2(n90169), .ZN(n86362) );
  NOR2_X1 U75729 ( .A1(n90155), .A2(n90154), .ZN(n86361) );
  AOI22_X1 U75730 ( .A1(n105761), .A2(n107185), .B1(n86364), .B2(n107181), 
        .ZN(n90176) );
  NOR2_X1 U75731 ( .A1(n90159), .A2(n90171), .ZN(n86364) );
  NOR2_X1 U75732 ( .A1(n90150), .A2(n90171), .ZN(n86363) );
  NAND2_X1 U75733 ( .A1(n90178), .A2(n90179), .ZN(n90174) );
  AOI22_X1 U75734 ( .A1(n105759), .A2(n107183), .B1(n105758), .B2(n107191), 
        .ZN(n90179) );
  NOR2_X1 U75735 ( .A1(n90152), .A2(n90169), .ZN(n86368) );
  NOR2_X1 U75736 ( .A1(n90159), .A2(n90169), .ZN(n86367) );
  AOI22_X1 U75737 ( .A1(n105757), .A2(n107179), .B1(n105756), .B2(n107189), 
        .ZN(n90178) );
  NOR2_X1 U75738 ( .A1(n90152), .A2(n90171), .ZN(n86370) );
  NOR2_X1 U75739 ( .A1(n90155), .A2(n90169), .ZN(n86369) );
  NAND2_X1 U75740 ( .A1(n90180), .A2(n90181), .ZN(n90173) );
  AOI22_X1 U75741 ( .A1(n105755), .A2(n69464), .B1(n105754), .B2(n69466), .ZN(
        n90181) );
  NOR2_X1 U75742 ( .A1(n90152), .A2(n90154), .ZN(n86374) );
  NOR2_X1 U75743 ( .A1(n90150), .A2(n90156), .ZN(n86373) );
  NAND2_X1 U75744 ( .A1(n90182), .A2(n90183), .ZN(n90150) );
  AOI22_X1 U75745 ( .A1(n105753), .A2(n69460), .B1(n105752), .B2(n107177), 
        .ZN(n90180) );
  NOR2_X1 U75746 ( .A1(n90155), .A2(n90171), .ZN(n86376) );
  NOR2_X1 U75747 ( .A1(n90159), .A2(n90156), .ZN(n86375) );
  NAND2_X1 U75748 ( .A1(n90184), .A2(n90185), .ZN(n90172) );
  AOI22_X1 U75749 ( .A1(n105751), .A2(n107207), .B1(n105750), .B2(n107197), 
        .ZN(n90185) );
  NOR2_X1 U75750 ( .A1(n90159), .A2(n90154), .ZN(n86380) );
  NOR2_X1 U75751 ( .A1(n90159), .A2(n90151), .ZN(n86379) );
  NAND2_X1 U75752 ( .A1(n90182), .A2(n90186), .ZN(n90159) );
  AOI22_X1 U75753 ( .A1(n105749), .A2(n69470), .B1(n86382), .B2(n107201), .ZN(
        n90184) );
  NOR2_X1 U75754 ( .A1(n90152), .A2(n90156), .ZN(n86382) );
  NAND2_X1 U75755 ( .A1(n90182), .A2(n90187), .ZN(n90152) );
  NOR2_X1 U75756 ( .A1(n90155), .A2(n90153), .ZN(n86381) );
  NAND2_X1 U75757 ( .A1(n90182), .A2(n90188), .ZN(n90155) );
  NOR2_X1 U75758 ( .A1(n90189), .A2(n90190), .ZN(n90182) );
  NAND2_X1 U75759 ( .A1(n90191), .A2(n90192), .ZN(n90140) );
  NOR4_X1 U75760 ( .A1(n90193), .A2(n90194), .A3(n90195), .A4(n90196), .ZN(
        n90192) );
  NAND2_X1 U75761 ( .A1(n90197), .A2(n90198), .ZN(n90196) );
  AOI22_X1 U75762 ( .A1(n105747), .A2(n107303), .B1(n105746), .B2(n107305), 
        .ZN(n90198) );
  NOR2_X1 U75763 ( .A1(n90166), .A2(n90154), .ZN(n86392) );
  NOR2_X1 U75764 ( .A1(n90170), .A2(n90156), .ZN(n86391) );
  AOI22_X1 U75765 ( .A1(n105745), .A2(n69620), .B1(n105744), .B2(n107304), 
        .ZN(n90197) );
  NOR2_X1 U75766 ( .A1(n90165), .A2(n90154), .ZN(n86394) );
  NOR2_X1 U75767 ( .A1(n90165), .A2(n90151), .ZN(n86393) );
  NAND2_X1 U75768 ( .A1(n90199), .A2(n90200), .ZN(n90195) );
  AOI22_X1 U75769 ( .A1(n105743), .A2(n69624), .B1(n105742), .B2(n69626), .ZN(
        n90200) );
  NOR2_X1 U75770 ( .A1(n90201), .A2(n90162), .ZN(n86398) );
  NOR2_X1 U75771 ( .A1(n90202), .A2(n90162), .ZN(n86397) );
  AOI22_X1 U75772 ( .A1(n105741), .A2(n107311), .B1(n105740), .B2(n107312), 
        .ZN(n90199) );
  NOR2_X1 U75773 ( .A1(n90202), .A2(n90161), .ZN(n86400) );
  NOR2_X1 U75774 ( .A1(n90166), .A2(n90151), .ZN(n86399) );
  NAND2_X1 U75775 ( .A1(n90203), .A2(n90204), .ZN(n90194) );
  AOI22_X1 U75776 ( .A1(n105739), .A2(n107308), .B1(n105738), .B2(n107310), 
        .ZN(n90204) );
  NOR2_X1 U75777 ( .A1(n90166), .A2(n90153), .ZN(n86404) );
  NOR2_X1 U75778 ( .A1(n90170), .A2(n90151), .ZN(n86403) );
  AOI22_X1 U75779 ( .A1(n105737), .A2(n107313), .B1(n86406), .B2(n107309), 
        .ZN(n90203) );
  NOR2_X1 U75780 ( .A1(n90165), .A2(n90153), .ZN(n86406) );
  NOR2_X1 U75781 ( .A1(n90201), .A2(n90161), .ZN(n86405) );
  NAND2_X1 U75782 ( .A1(n90205), .A2(n90206), .ZN(n90193) );
  AOI22_X1 U75783 ( .A1(n105735), .A2(n107318), .B1(n105734), .B2(n69631), 
        .ZN(n90206) );
  NOR2_X1 U75784 ( .A1(n90202), .A2(n90171), .ZN(n86410) );
  NOR2_X1 U75785 ( .A1(n90201), .A2(n90171), .ZN(n86409) );
  AOI22_X1 U75786 ( .A1(n105733), .A2(n107317), .B1(n105732), .B2(n69629), 
        .ZN(n90205) );
  NOR2_X1 U75787 ( .A1(n90207), .A2(n90161), .ZN(n86412) );
  NOR2_X1 U75788 ( .A1(n90202), .A2(n90169), .ZN(n86411) );
  NOR4_X1 U75789 ( .A1(n90208), .A2(n90209), .A3(n90210), .A4(n90211), .ZN(
        n90191) );
  NAND2_X1 U75790 ( .A1(n90212), .A2(n90213), .ZN(n90211) );
  AOI22_X1 U75791 ( .A1(n105731), .A2(n107298), .B1(n105730), .B2(n107289), 
        .ZN(n90213) );
  NOR2_X1 U75792 ( .A1(n90170), .A2(n90161), .ZN(n86420) );
  NOR2_X1 U75793 ( .A1(n90166), .A2(n90171), .ZN(n86419) );
  AOI22_X1 U75794 ( .A1(n105729), .A2(n107291), .B1(n105728), .B2(n69603), 
        .ZN(n90212) );
  NOR2_X1 U75795 ( .A1(n90165), .A2(n90171), .ZN(n86422) );
  NOR2_X1 U75796 ( .A1(n90165), .A2(n90162), .ZN(n86421) );
  NAND2_X1 U75797 ( .A1(n90214), .A2(n90215), .ZN(n90210) );
  AOI22_X1 U75798 ( .A1(n105727), .A2(n107296), .B1(n105726), .B2(n107300), 
        .ZN(n90215) );
  NOR2_X1 U75799 ( .A1(n90160), .A2(n90154), .ZN(n86426) );
  NOR2_X1 U75800 ( .A1(n90170), .A2(n90169), .ZN(n86425) );
  AOI22_X1 U75801 ( .A1(n105725), .A2(n107302), .B1(n105724), .B2(n107299), 
        .ZN(n90214) );
  NOR2_X1 U75802 ( .A1(n90166), .A2(n90169), .ZN(n86428) );
  NOR2_X1 U75803 ( .A1(n90170), .A2(n90154), .ZN(n86427) );
  NAND2_X1 U75804 ( .A1(n90216), .A2(n90217), .ZN(n90209) );
  AOI22_X1 U75805 ( .A1(n105723), .A2(n69612), .B1(n105722), .B2(n107295), 
        .ZN(n90217) );
  NOR2_X1 U75806 ( .A1(n90170), .A2(n90171), .ZN(n86432) );
  NOR2_X1 U75807 ( .A1(n90165), .A2(n90156), .ZN(n86431) );
  AOI22_X1 U75808 ( .A1(n105721), .A2(n107297), .B1(n105720), .B2(n107301), 
        .ZN(n90216) );
  NOR2_X1 U75809 ( .A1(n90160), .A2(n90156), .ZN(n86434) );
  NOR2_X1 U75810 ( .A1(n90165), .A2(n90169), .ZN(n86433) );
  NAND2_X1 U75811 ( .A1(n90218), .A2(n90183), .ZN(n90165) );
  NAND2_X1 U75812 ( .A1(n90219), .A2(n90220), .ZN(n90208) );
  AOI22_X1 U75813 ( .A1(n105719), .A2(n107307), .B1(n105718), .B2(n69616), 
        .ZN(n90220) );
  NOR2_X1 U75814 ( .A1(n90160), .A2(n90151), .ZN(n86438) );
  NOR2_X1 U75815 ( .A1(n90170), .A2(n90153), .ZN(n86437) );
  NAND2_X1 U75816 ( .A1(n90218), .A2(n90186), .ZN(n90170) );
  AOI22_X1 U75817 ( .A1(n105717), .A2(n69614), .B1(n86440), .B2(n107306), .ZN(
        n90219) );
  NOR2_X1 U75818 ( .A1(n90160), .A2(n90153), .ZN(n86440) );
  NAND2_X1 U75819 ( .A1(n90218), .A2(n90188), .ZN(n90160) );
  NOR2_X1 U75820 ( .A1(n90166), .A2(n90156), .ZN(n86439) );
  NAND2_X1 U75821 ( .A1(n90218), .A2(n90187), .ZN(n90166) );
  NOR2_X1 U75822 ( .A1(n90189), .A2(n107093), .ZN(n90218) );
  NAND2_X1 U75823 ( .A1(n90221), .A2(n90222), .ZN(n90139) );
  NOR4_X1 U75824 ( .A1(n90223), .A2(n90224), .A3(n90225), .A4(n90226), .ZN(
        n90222) );
  NAND2_X1 U75825 ( .A1(n90227), .A2(n90228), .ZN(n90226) );
  AOI22_X1 U75826 ( .A1(n105715), .A2(n69654), .B1(n105714), .B2(n107328), 
        .ZN(n90228) );
  NOR2_X1 U75827 ( .A1(n90207), .A2(n90154), .ZN(n86450) );
  NOR2_X1 U75828 ( .A1(n90207), .A2(n90151), .ZN(n86449) );
  AOI22_X1 U75829 ( .A1(n105713), .A2(n107332), .B1(n105712), .B2(n107331), 
        .ZN(n90227) );
  NOR2_X1 U75830 ( .A1(n90201), .A2(n90151), .ZN(n86452) );
  NOR2_X1 U75831 ( .A1(n90229), .A2(n90153), .ZN(n86451) );
  NAND2_X1 U75832 ( .A1(n90230), .A2(n90231), .ZN(n90225) );
  AOI22_X1 U75833 ( .A1(n105711), .A2(n107337), .B1(n105710), .B2(n107336), 
        .ZN(n90231) );
  NOR2_X1 U75834 ( .A1(n90162), .A2(n90232), .ZN(n86456) );
  NOR2_X1 U75835 ( .A1(n90161), .A2(n90233), .ZN(n86455) );
  AOI22_X1 U75836 ( .A1(n105709), .A2(n107327), .B1(n105708), .B2(n107329), 
        .ZN(n90230) );
  NOR2_X1 U75837 ( .A1(n90202), .A2(n90153), .ZN(n86458) );
  NOR2_X1 U75838 ( .A1(n90229), .A2(n90156), .ZN(n86457) );
  NAND2_X1 U75839 ( .A1(n90234), .A2(n90235), .ZN(n90224) );
  AOI22_X1 U75840 ( .A1(n105707), .A2(n107338), .B1(n105706), .B2(n107334), 
        .ZN(n90235) );
  NOR2_X1 U75841 ( .A1(n90207), .A2(n90153), .ZN(n86462) );
  NOR2_X1 U75842 ( .A1(n90161), .A2(n90236), .ZN(n86461) );
  AOI22_X1 U75843 ( .A1(n105705), .A2(n69658), .B1(n105704), .B2(n69660), .ZN(
        n90234) );
  NOR2_X1 U75844 ( .A1(n90162), .A2(n90236), .ZN(n86464) );
  NOR2_X1 U75845 ( .A1(n90162), .A2(n90233), .ZN(n86463) );
  NAND2_X1 U75846 ( .A1(n90237), .A2(n90238), .ZN(n90223) );
  AOI22_X1 U75847 ( .A1(n105703), .A2(n107341), .B1(n105702), .B2(n69666), 
        .ZN(n90238) );
  NOR2_X1 U75848 ( .A1(n90169), .A2(n90233), .ZN(n86468) );
  NOR2_X1 U75849 ( .A1(n90171), .A2(n90232), .ZN(n86467) );
  AOI22_X1 U75850 ( .A1(n105701), .A2(n107333), .B1(n105700), .B2(n107335), 
        .ZN(n90237) );
  NOR2_X1 U75851 ( .A1(n90161), .A2(n90232), .ZN(n86470) );
  NOR2_X1 U75852 ( .A1(n90229), .A2(n90151), .ZN(n86469) );
  NOR4_X1 U75853 ( .A1(n90239), .A2(n90240), .A3(n90241), .A4(n90242), .ZN(
        n90221) );
  NAND2_X1 U75854 ( .A1(n90243), .A2(n90244), .ZN(n90242) );
  AOI22_X1 U75855 ( .A1(n105699), .A2(n107316), .B1(n105698), .B2(n107321), 
        .ZN(n90244) );
  NOR2_X1 U75856 ( .A1(n90207), .A2(n90171), .ZN(n86478) );
  NOR2_X1 U75857 ( .A1(n90207), .A2(n90162), .ZN(n86477) );
  AOI22_X1 U75858 ( .A1(n105697), .A2(n107315), .B1(n105696), .B2(n69634), 
        .ZN(n90243) );
  NOR2_X1 U75859 ( .A1(n90201), .A2(n90169), .ZN(n86480) );
  NOR2_X1 U75860 ( .A1(n90229), .A2(n90162), .ZN(n86479) );
  NAND2_X1 U75861 ( .A1(n90245), .A2(n90246), .ZN(n90241) );
  AOI22_X1 U75862 ( .A1(n105695), .A2(n69643), .B1(n105694), .B2(n107323), 
        .ZN(n90246) );
  NOR2_X1 U75863 ( .A1(n90202), .A2(n90154), .ZN(n86484) );
  NOR2_X1 U75864 ( .A1(n90229), .A2(n90154), .ZN(n86483) );
  AOI22_X1 U75865 ( .A1(n105693), .A2(n107324), .B1(n105692), .B2(n107314), 
        .ZN(n90245) );
  NOR2_X1 U75866 ( .A1(n90229), .A2(n90161), .ZN(n86486) );
  NOR2_X1 U75867 ( .A1(n90202), .A2(n90156), .ZN(n86485) );
  NAND2_X1 U75868 ( .A1(n90247), .A2(n90248), .ZN(n90240) );
  AOI22_X1 U75869 ( .A1(n105691), .A2(n107322), .B1(n105690), .B2(n107326), 
        .ZN(n90248) );
  NOR2_X1 U75870 ( .A1(n90201), .A2(n90156), .ZN(n86490) );
  NOR2_X1 U75871 ( .A1(n90207), .A2(n90169), .ZN(n86489) );
  AOI22_X1 U75872 ( .A1(n105689), .A2(n107320), .B1(n105688), .B2(n107325), 
        .ZN(n90247) );
  NOR2_X1 U75873 ( .A1(n90201), .A2(n90154), .ZN(n86492) );
  NOR2_X1 U75874 ( .A1(n90229), .A2(n90169), .ZN(n86491) );
  NAND2_X1 U75875 ( .A1(n90249), .A2(n90250), .ZN(n90239) );
  AOI22_X1 U75876 ( .A1(n105687), .A2(n69648), .B1(n105686), .B2(n107330), 
        .ZN(n90250) );
  NOR2_X1 U75877 ( .A1(n90201), .A2(n90153), .ZN(n86496) );
  NAND2_X1 U75878 ( .A1(n90251), .A2(n90186), .ZN(n90201) );
  NOR2_X1 U75879 ( .A1(n90202), .A2(n90151), .ZN(n86495) );
  NAND2_X1 U75880 ( .A1(n90251), .A2(n90188), .ZN(n90202) );
  AOI22_X1 U75881 ( .A1(n105685), .A2(n69646), .B1(n105684), .B2(n107319), 
        .ZN(n90249) );
  NOR2_X1 U75882 ( .A1(n90229), .A2(n90171), .ZN(n86498) );
  NAND2_X1 U75883 ( .A1(n90251), .A2(n90183), .ZN(n90229) );
  NOR2_X1 U75884 ( .A1(n90207), .A2(n90156), .ZN(n86497) );
  NAND2_X1 U75885 ( .A1(n90251), .A2(n90187), .ZN(n90207) );
  NOR2_X1 U75886 ( .A1(n90190), .A2(n107059), .ZN(n90251) );
  NAND2_X1 U75887 ( .A1(n90252), .A2(n90253), .ZN(n90138) );
  NOR4_X1 U75888 ( .A1(n90254), .A2(n90255), .A3(n90256), .A4(n90257), .ZN(
        n90253) );
  NAND2_X1 U75889 ( .A1(n90258), .A2(n90259), .ZN(n90257) );
  AOI22_X1 U75890 ( .A1(n105683), .A2(n107359), .B1(n105682), .B2(n107358), 
        .ZN(n90259) );
  NOR2_X1 U75891 ( .A1(n90236), .A2(n90151), .ZN(n86508) );
  NOR2_X1 U75892 ( .A1(n90153), .A2(n90260), .ZN(n86507) );
  AOI22_X1 U75893 ( .A1(n105681), .A2(n69682), .B1(n105680), .B2(n107356), 
        .ZN(n90258) );
  NOR2_X1 U75894 ( .A1(n90232), .A2(n90151), .ZN(n86510) );
  NOR2_X1 U75895 ( .A1(n90233), .A2(n90151), .ZN(n86509) );
  NAND2_X1 U75896 ( .A1(n90261), .A2(n90262), .ZN(n90256) );
  AOI22_X1 U75897 ( .A1(n105679), .A2(n107354), .B1(n86514), .B2(n107357), 
        .ZN(n90262) );
  NOR2_X1 U75898 ( .A1(n90233), .A2(n90153), .ZN(n86514) );
  NOR2_X1 U75899 ( .A1(n90156), .A2(n90260), .ZN(n86513) );
  AOI22_X1 U75900 ( .A1(n86515), .A2(n69688), .B1(n105677), .B2(n107355), .ZN(
        n90261) );
  NOR2_X1 U75901 ( .A1(n90232), .A2(n90153), .ZN(n86516) );
  AND2_X2 U75902 ( .A1(n90263), .A2(n90188), .ZN(n86515) );
  NAND2_X1 U75903 ( .A1(n90264), .A2(n90265), .ZN(n90255) );
  AOI22_X1 U75904 ( .A1(n86519), .A2(n107364), .B1(n86520), .B2(n69694), .ZN(
        n90265) );
  AND2_X2 U75905 ( .A1(n90263), .A2(n90187), .ZN(n86520) );
  AND2_X2 U75906 ( .A1(n90183), .A2(n90263), .ZN(n86519) );
  AOI22_X1 U75907 ( .A1(n86521), .A2(n107362), .B1(n86522), .B2(n107363), .ZN(
        n90264) );
  AND2_X2 U75908 ( .A1(n90183), .A2(n90266), .ZN(n86522) );
  AND2_X2 U75909 ( .A1(n90263), .A2(n90186), .ZN(n86521) );
  NOR2_X1 U75910 ( .A1(n90267), .A2(n59435), .ZN(n90263) );
  NAND2_X1 U75911 ( .A1(n90268), .A2(n90269), .ZN(n90254) );
  AOI22_X1 U75912 ( .A1(n105676), .A2(n107360), .B1(n86526), .B2(n69689), .ZN(
        n90269) );
  AND2_X2 U75913 ( .A1(n90186), .A2(n90266), .ZN(n86526) );
  NOR2_X1 U75914 ( .A1(n90151), .A2(n90260), .ZN(n86525) );
  OR2_X1 U75915 ( .A1(n90270), .A2(n90271), .ZN(n90151) );
  AOI22_X1 U75916 ( .A1(n86527), .A2(n107365), .B1(n86528), .B2(n107361), .ZN(
        n90268) );
  AND2_X2 U75917 ( .A1(n90188), .A2(n90266), .ZN(n86528) );
  AND2_X2 U75918 ( .A1(n90266), .A2(n90187), .ZN(n86527) );
  NOR2_X1 U75919 ( .A1(n90267), .A2(n107132), .ZN(n90266) );
  NAND2_X1 U75920 ( .A1(n90272), .A2(n90135), .ZN(n90267) );
  NOR4_X1 U75921 ( .A1(n90273), .A2(n90274), .A3(n90275), .A4(n90276), .ZN(
        n90252) );
  NAND2_X1 U75922 ( .A1(n90277), .A2(n90278), .ZN(n90276) );
  AOI22_X1 U75923 ( .A1(n105675), .A2(n107340), .B1(n105674), .B2(n107344), 
        .ZN(n90278) );
  NOR2_X1 U75924 ( .A1(n90169), .A2(n90236), .ZN(n86536) );
  NOR2_X1 U75925 ( .A1(n90162), .A2(n90260), .ZN(n86535) );
  OR2_X1 U75926 ( .A1(n90106), .A2(n107100), .ZN(n90162) );
  AOI22_X1 U75927 ( .A1(n105673), .A2(n107343), .B1(n105672), .B2(n69665), 
        .ZN(n90277) );
  NOR2_X1 U75928 ( .A1(n90171), .A2(n90233), .ZN(n86538) );
  NOR2_X1 U75929 ( .A1(n90171), .A2(n90236), .ZN(n86537) );
  NAND2_X1 U75930 ( .A1(n90279), .A2(n90280), .ZN(n90275) );
  AOI22_X1 U75931 ( .A1(n105671), .A2(n107350), .B1(n105670), .B2(n107339), 
        .ZN(n90280) );
  NOR2_X1 U75932 ( .A1(n90161), .A2(n90260), .ZN(n86542) );
  NOR2_X1 U75935 ( .A1(n90233), .A2(n90156), .ZN(n86541) );
  AOI22_X1 U75936 ( .A1(n105669), .A2(n107342), .B1(n86544), .B2(n107347), 
        .ZN(n90279) );
  NOR2_X1 U75937 ( .A1(n90154), .A2(n90232), .ZN(n86544) );
  NOR2_X1 U75938 ( .A1(n90169), .A2(n90232), .ZN(n86543) );
  NAND2_X1 U75939 ( .A1(n90282), .A2(n90283), .ZN(n90274) );
  AOI22_X1 U75940 ( .A1(n105667), .A2(n107346), .B1(n105666), .B2(n107351), 
        .ZN(n90283) );
  NOR2_X1 U75941 ( .A1(n90154), .A2(n90236), .ZN(n86548) );
  NOR2_X1 U75942 ( .A1(n90169), .A2(n90260), .ZN(n86547) );
  OR2_X1 U75943 ( .A1(n90270), .A2(n107100), .ZN(n90169) );
  NAND2_X1 U75944 ( .A1(n107132), .A2(n107139), .ZN(n90270) );
  AOI22_X1 U75945 ( .A1(n105665), .A2(n107353), .B1(n105664), .B2(n107349), 
        .ZN(n90282) );
  NOR2_X1 U75946 ( .A1(n90154), .A2(n90233), .ZN(n86550) );
  NAND2_X1 U75947 ( .A1(n90186), .A2(n90284), .ZN(n90233) );
  NOR2_X1 U75948 ( .A1(n107137), .A2(n59441), .ZN(n90186) );
  NOR2_X1 U75949 ( .A1(n90154), .A2(n90260), .ZN(n86549) );
  OR2_X1 U75950 ( .A1(n90121), .A2(n90271), .ZN(n90154) );
  NAND2_X1 U75951 ( .A1(n59443), .A2(n59435), .ZN(n90121) );
  NAND2_X1 U75952 ( .A1(n90285), .A2(n90286), .ZN(n90273) );
  AOI22_X1 U75953 ( .A1(n105663), .A2(n69683), .B1(n105662), .B2(n107345), 
        .ZN(n90286) );
  NOR2_X1 U75954 ( .A1(n90171), .A2(n90260), .ZN(n86554) );
  NAND2_X1 U75955 ( .A1(n90187), .A2(n90284), .ZN(n90260) );
  NOR2_X1 U75956 ( .A1(n59442), .A2(n59441), .ZN(n90187) );
  NOR2_X1 U75959 ( .A1(n90236), .A2(n90153), .ZN(n86553) );
  AOI22_X1 U75962 ( .A1(n86555), .A2(n107348), .B1(n105660), .B2(n107352), 
        .ZN(n90285) );
  NOR2_X1 U75963 ( .A1(n90236), .A2(n90156), .ZN(n86556) );
  NAND2_X1 U75964 ( .A1(n90183), .A2(n90284), .ZN(n90236) );
  NOR2_X1 U75965 ( .A1(n107134), .A2(n59442), .ZN(n90183) );
  NOR2_X1 U75966 ( .A1(n90232), .A2(n90156), .ZN(n86555) );
  OR2_X1 U75967 ( .A1(n90271), .A2(n90106), .ZN(n90156) );
  NAND2_X1 U75968 ( .A1(n59443), .A2(n107132), .ZN(n90106) );
  XOR2_X1 U75969 ( .A(n107139), .B(n90134), .Z(n90271) );
  NAND2_X1 U75970 ( .A1(n90188), .A2(n90284), .ZN(n90232) );
  NOR2_X1 U75971 ( .A1(n107093), .A2(n107059), .ZN(n90284) );
  XOR2_X1 U75972 ( .A(n90272), .B(n90135), .Z(n90189) );
  NOR2_X1 U75975 ( .A1(n90292), .A2(n90132), .ZN(n90272) );
  XOR2_X1 U75976 ( .A(n90132), .B(n90292), .Z(n90190) );
  NAND2_X1 U75977 ( .A1(n59443), .A2(n90134), .ZN(n90292) );
  OAI21_X1 U75978 ( .B1(n59443), .B2(n90293), .A(n90290), .ZN(n90134) );
  XOR2_X1 U75979 ( .A(n90291), .B(n90290), .Z(n90132) );
  NAND2_X1 U75980 ( .A1(n90293), .A2(n59443), .ZN(n90290) );
  NOR2_X1 U75981 ( .A1(n107134), .A2(n107137), .ZN(n90188) );
  AOI21_X1 U75982 ( .B1(n90295), .B2(n86303), .A(n90296), .ZN(n90294) );
  OAI21_X1 U75983 ( .B1(n90297), .B2(n105659), .A(n90299), .ZN(n90296) );
  OAI21_X1 U75984 ( .B1(n90300), .B2(n90301), .A(n90302), .ZN(n90299) );
  OAI21_X1 U75985 ( .B1(n102179), .B2(n90303), .A(n90304), .ZN(n90301) );
  AOI22_X1 U75986 ( .A1(n90305), .A2(n107941), .B1(n90306), .B2(n70424), .ZN(
        n90304) );
  NAND2_X1 U75987 ( .A1(n90307), .A2(n90308), .ZN(n90300) );
  AOI22_X1 U75988 ( .A1(n90309), .A2(n107946), .B1(n105653), .B2(n107943), 
        .ZN(n90308) );
  AOI22_X1 U75989 ( .A1(n90311), .A2(n70422), .B1(n90312), .B2(n107942), .ZN(
        n90307) );
  NOR4_X1 U75990 ( .A1(n90313), .A2(n90314), .A3(n90315), .A4(n90316), .ZN(
        n90297) );
  NAND2_X1 U75991 ( .A1(n90317), .A2(n90318), .ZN(n90316) );
  NOR4_X1 U75992 ( .A1(n90319), .A2(n90320), .A3(n90321), .A4(n90322), .ZN(
        n90318) );
  NAND2_X1 U75993 ( .A1(n90323), .A2(n90324), .ZN(n90322) );
  AOI22_X1 U75994 ( .A1(n90325), .A2(n107922), .B1(n90326), .B2(n107923), .ZN(
        n90324) );
  AOI22_X1 U75995 ( .A1(n90327), .A2(n107931), .B1(n90328), .B2(n107929), .ZN(
        n90323) );
  NAND2_X1 U75996 ( .A1(n90329), .A2(n90330), .ZN(n90321) );
  AOI22_X1 U75997 ( .A1(n90331), .A2(n70291), .B1(n90332), .B2(n107926), .ZN(
        n90330) );
  AOI22_X1 U75998 ( .A1(n90333), .A2(n70395), .B1(n90334), .B2(n107855), .ZN(
        n90329) );
  NAND2_X1 U75999 ( .A1(n90335), .A2(n90336), .ZN(n90320) );
  AOI22_X1 U76000 ( .A1(n90337), .A2(n107859), .B1(n90338), .B2(n70295), .ZN(
        n90336) );
  AOI22_X1 U76001 ( .A1(n90339), .A2(n107927), .B1(n90340), .B2(n107924), .ZN(
        n90335) );
  NAND2_X1 U76002 ( .A1(n90341), .A2(n90342), .ZN(n90319) );
  AOI22_X1 U76003 ( .A1(n90343), .A2(n107857), .B1(n90344), .B2(n107861), .ZN(
        n90342) );
  AOI22_X1 U76004 ( .A1(n90345), .A2(n107860), .B1(n90346), .B2(n70297), .ZN(
        n90341) );
  NOR4_X1 U76005 ( .A1(n90347), .A2(n90348), .A3(n90349), .A4(n90350), .ZN(
        n90317) );
  NAND2_X1 U76006 ( .A1(n90351), .A2(n90352), .ZN(n90350) );
  AOI22_X1 U76007 ( .A1(n90353), .A2(n107932), .B1(n90354), .B2(n107935), .ZN(
        n90352) );
  AOI22_X1 U76008 ( .A1(n90355), .A2(n107936), .B1(n90356), .B2(n107938), .ZN(
        n90351) );
  NAND2_X1 U76009 ( .A1(n90357), .A2(n90358), .ZN(n90349) );
  AOI22_X1 U76010 ( .A1(n90359), .A2(n107937), .B1(n90360), .B2(n107933), .ZN(
        n90358) );
  AOI22_X1 U76011 ( .A1(n90361), .A2(n107939), .B1(n90362), .B2(n107934), .ZN(
        n90357) );
  NAND2_X1 U76012 ( .A1(n90363), .A2(n90364), .ZN(n90348) );
  AOI22_X1 U76013 ( .A1(n90365), .A2(n70405), .B1(n90366), .B2(n70404), .ZN(
        n90364) );
  AOI22_X1 U76014 ( .A1(n90367), .A2(n70407), .B1(n90368), .B2(n107940), .ZN(
        n90363) );
  NAND2_X1 U76015 ( .A1(n90369), .A2(n90370), .ZN(n90347) );
  AOI22_X1 U76016 ( .A1(n90371), .A2(n107925), .B1(n90372), .B2(n107930), .ZN(
        n90370) );
  AOI22_X1 U76017 ( .A1(n90373), .A2(n70402), .B1(n90374), .B2(n107928), .ZN(
        n90369) );
  NAND2_X1 U76018 ( .A1(n90375), .A2(n90376), .ZN(n90315) );
  NOR4_X1 U76019 ( .A1(n90377), .A2(n90378), .A3(n90379), .A4(n90380), .ZN(
        n90376) );
  NAND2_X1 U76020 ( .A1(n90381), .A2(n90382), .ZN(n90380) );
  AOI22_X1 U76021 ( .A1(n90383), .A2(n107869), .B1(n90384), .B2(n107871), .ZN(
        n90382) );
  AOI22_X1 U76022 ( .A1(n90385), .A2(n70320), .B1(n90386), .B2(n107870), .ZN(
        n90381) );
  NAND2_X1 U76023 ( .A1(n90387), .A2(n90388), .ZN(n90379) );
  AOI22_X1 U76024 ( .A1(n90389), .A2(n70324), .B1(n90390), .B2(n70326), .ZN(
        n90388) );
  AOI22_X1 U76025 ( .A1(n90391), .A2(n107875), .B1(n90392), .B2(n107876), .ZN(
        n90387) );
  NAND2_X1 U76026 ( .A1(n90393), .A2(n90394), .ZN(n90378) );
  AOI22_X1 U76027 ( .A1(n90395), .A2(n107873), .B1(n90396), .B2(n70321), .ZN(
        n90394) );
  AOI22_X1 U76028 ( .A1(n90397), .A2(n107877), .B1(n90398), .B2(n107874), .ZN(
        n90393) );
  NAND2_X1 U76029 ( .A1(n90399), .A2(n90400), .ZN(n90377) );
  AOI22_X1 U76030 ( .A1(n90401), .A2(n107881), .B1(n90402), .B2(n70331), .ZN(
        n90400) );
  AOI22_X1 U76031 ( .A1(n90403), .A2(n107880), .B1(n90404), .B2(n70329), .ZN(
        n90399) );
  NOR4_X1 U76032 ( .A1(n90405), .A2(n90406), .A3(n90407), .A4(n90408), .ZN(
        n90375) );
  NAND2_X1 U76033 ( .A1(n90409), .A2(n90410), .ZN(n90408) );
  AOI22_X1 U76034 ( .A1(n90411), .A2(n107864), .B1(n90412), .B2(n107856), .ZN(
        n90410) );
  AOI22_X1 U76035 ( .A1(n90413), .A2(n107858), .B1(n90414), .B2(n70303), .ZN(
        n90409) );
  NAND2_X1 U76036 ( .A1(n90415), .A2(n90416), .ZN(n90407) );
  AOI22_X1 U76037 ( .A1(n90417), .A2(n107863), .B1(n90418), .B2(n107866), .ZN(
        n90416) );
  AOI22_X1 U76038 ( .A1(n90419), .A2(n107868), .B1(n90420), .B2(n107865), .ZN(
        n90415) );
  NAND2_X1 U76039 ( .A1(n90421), .A2(n90422), .ZN(n90406) );
  AOI22_X1 U76040 ( .A1(n90423), .A2(n70312), .B1(n90424), .B2(n107862), .ZN(
        n90422) );
  AOI22_X1 U76041 ( .A1(n90425), .A2(n70304), .B1(n90426), .B2(n70308), .ZN(
        n90421) );
  NAND2_X1 U76042 ( .A1(n90427), .A2(n90428), .ZN(n90405) );
  AOI22_X1 U76043 ( .A1(n90429), .A2(n70317), .B1(n90430), .B2(n70316), .ZN(
        n90428) );
  AOI22_X1 U76044 ( .A1(n90431), .A2(n70314), .B1(n90432), .B2(n107872), .ZN(
        n90427) );
  NAND2_X1 U76045 ( .A1(n90433), .A2(n90434), .ZN(n90314) );
  NOR4_X1 U76046 ( .A1(n90435), .A2(n90436), .A3(n90437), .A4(n90438), .ZN(
        n90434) );
  NAND2_X1 U76047 ( .A1(n90439), .A2(n90440), .ZN(n90438) );
  AOI22_X1 U76048 ( .A1(n90441), .A2(n70354), .B1(n90442), .B2(n107890), .ZN(
        n90440) );
  AOI22_X1 U76049 ( .A1(n90443), .A2(n107893), .B1(n90444), .B2(n70350), .ZN(
        n90439) );
  NAND2_X1 U76050 ( .A1(n90445), .A2(n90446), .ZN(n90437) );
  AOI22_X1 U76051 ( .A1(n90447), .A2(n107897), .B1(n90448), .B2(n107896), .ZN(
        n90446) );
  AOI22_X1 U76052 ( .A1(n90449), .A2(n107889), .B1(n90450), .B2(n107891), .ZN(
        n90445) );
  NAND2_X1 U76053 ( .A1(n90451), .A2(n90452), .ZN(n90436) );
  AOI22_X1 U76054 ( .A1(n90453), .A2(n107898), .B1(n90454), .B2(n107895), .ZN(
        n90452) );
  AOI22_X1 U76055 ( .A1(n90455), .A2(n70358), .B1(n90456), .B2(n70360), .ZN(
        n90451) );
  NAND2_X1 U76056 ( .A1(n90457), .A2(n90458), .ZN(n90435) );
  AOI22_X1 U76057 ( .A1(n90459), .A2(n70363), .B1(n90460), .B2(n70366), .ZN(
        n90458) );
  AOI22_X1 U76058 ( .A1(n90461), .A2(n107894), .B1(n90462), .B2(n70355), .ZN(
        n90457) );
  NOR4_X1 U76059 ( .A1(n90463), .A2(n90464), .A3(n90465), .A4(n90466), .ZN(
        n90433) );
  NAND2_X1 U76060 ( .A1(n90467), .A2(n90468), .ZN(n90466) );
  AOI22_X1 U76061 ( .A1(n90469), .A2(n70330), .B1(n90470), .B2(n107884), .ZN(
        n90468) );
  AOI22_X1 U76062 ( .A1(n90471), .A2(n107879), .B1(n90472), .B2(n70334), .ZN(
        n90467) );
  NAND2_X1 U76063 ( .A1(n90473), .A2(n90474), .ZN(n90465) );
  AOI22_X1 U76064 ( .A1(n90475), .A2(n70343), .B1(n90476), .B2(n107886), .ZN(
        n90474) );
  AOI22_X1 U76065 ( .A1(n90477), .A2(n107887), .B1(n90478), .B2(n107878), .ZN(
        n90473) );
  NAND2_X1 U76066 ( .A1(n90479), .A2(n90480), .ZN(n90464) );
  AOI22_X1 U76067 ( .A1(n90481), .A2(n107885), .B1(n90482), .B2(n70342), .ZN(
        n90480) );
  AOI22_X1 U76068 ( .A1(n90483), .A2(n107883), .B1(n90484), .B2(n107888), .ZN(
        n90479) );
  NAND2_X1 U76069 ( .A1(n90485), .A2(n90486), .ZN(n90463) );
  AOI22_X1 U76070 ( .A1(n90487), .A2(n70348), .B1(n90488), .B2(n107892), .ZN(
        n90486) );
  AOI22_X1 U76071 ( .A1(n90489), .A2(n70346), .B1(n90490), .B2(n107882), .ZN(
        n90485) );
  NAND2_X1 U76072 ( .A1(n90491), .A2(n90492), .ZN(n90313) );
  NOR4_X1 U76073 ( .A1(n90493), .A2(n90494), .A3(n90495), .A4(n90496), .ZN(
        n90492) );
  NAND2_X1 U76074 ( .A1(n90497), .A2(n90498), .ZN(n90496) );
  AOI22_X1 U76075 ( .A1(n90499), .A2(n107914), .B1(n90500), .B2(n107913), .ZN(
        n90498) );
  AOI22_X1 U76076 ( .A1(n90501), .A2(n70382), .B1(n90502), .B2(n107911), .ZN(
        n90497) );
  NAND2_X1 U76077 ( .A1(n90503), .A2(n90504), .ZN(n90495) );
  AOI22_X1 U76078 ( .A1(n90505), .A2(n107909), .B1(n90506), .B2(n107912), .ZN(
        n90504) );
  AOI22_X1 U76079 ( .A1(n90507), .A2(n70388), .B1(n90508), .B2(n107910), .ZN(
        n90503) );
  NAND2_X1 U76080 ( .A1(n90509), .A2(n90510), .ZN(n90494) );
  AOI22_X1 U76081 ( .A1(n105650), .A2(n107919), .B1(n90512), .B2(n70394), .ZN(
        n90510) );
  AOI22_X1 U76082 ( .A1(n90513), .A2(n107917), .B1(n90514), .B2(n107918), .ZN(
        n90509) );
  NAND2_X1 U76083 ( .A1(n90515), .A2(n90516), .ZN(n90493) );
  AOI22_X1 U76084 ( .A1(n90517), .A2(n70386), .B1(n90518), .B2(n107916), .ZN(
        n90516) );
  AOI22_X1 U76085 ( .A1(n90519), .A2(n107920), .B1(n105644), .B2(n107915), 
        .ZN(n90515) );
  NOR4_X1 U76086 ( .A1(n90521), .A2(n90522), .A3(n90523), .A4(n90524), .ZN(
        n90491) );
  NAND2_X1 U76087 ( .A1(n90525), .A2(n90526), .ZN(n90524) );
  AOI22_X1 U76088 ( .A1(n90527), .A2(n107900), .B1(n90528), .B2(n107901), .ZN(
        n90526) );
  AOI22_X1 U76089 ( .A1(n90529), .A2(n70367), .B1(n90530), .B2(n70365), .ZN(
        n90525) );
  NAND2_X1 U76090 ( .A1(n90531), .A2(n90532), .ZN(n90523) );
  AOI22_X1 U76091 ( .A1(n90533), .A2(n107906), .B1(n90534), .B2(n107899), .ZN(
        n90532) );
  AOI22_X1 U76092 ( .A1(n90535), .A2(n70364), .B1(n90536), .B2(n107903), .ZN(
        n90531) );
  NAND2_X1 U76093 ( .A1(n90537), .A2(n90538), .ZN(n90522) );
  AOI22_X1 U76094 ( .A1(n90539), .A2(n107902), .B1(n90540), .B2(n107907), .ZN(
        n90538) );
  AOI22_X1 U76095 ( .A1(n90541), .A2(n107908), .B1(n90542), .B2(n107905), .ZN(
        n90537) );
  NAND2_X1 U76096 ( .A1(n90543), .A2(n90544), .ZN(n90521) );
  AOI22_X1 U76097 ( .A1(n90545), .A2(n70383), .B1(n90546), .B2(n70369), .ZN(
        n90544) );
  AOI22_X1 U76098 ( .A1(n90547), .A2(n70372), .B1(n90548), .B2(n70376), .ZN(
        n90543) );
  AOI21_X1 U76099 ( .B1(n90295), .B2(n86558), .A(n90550), .ZN(n90549) );
  OAI21_X1 U76100 ( .B1(n90551), .B2(n105659), .A(n90552), .ZN(n90550) );
  OAI21_X1 U76101 ( .B1(n90553), .B2(n90554), .A(n90302), .ZN(n90552) );
  OAI21_X1 U76102 ( .B1(n102165), .B2(n90303), .A(n90555), .ZN(n90554) );
  AOI22_X1 U76103 ( .A1(n90305), .A2(n108037), .B1(n90306), .B2(n70566), .ZN(
        n90555) );
  NAND2_X1 U76104 ( .A1(n90556), .A2(n90557), .ZN(n90553) );
  AOI22_X1 U76105 ( .A1(n90309), .A2(n108042), .B1(n105653), .B2(n108039), 
        .ZN(n90557) );
  AOI22_X1 U76106 ( .A1(n90311), .A2(n70564), .B1(n90312), .B2(n108038), .ZN(
        n90556) );
  NOR4_X1 U76107 ( .A1(n90558), .A2(n90559), .A3(n90560), .A4(n90561), .ZN(
        n90551) );
  NAND2_X1 U76108 ( .A1(n90562), .A2(n90563), .ZN(n90561) );
  NOR4_X1 U76109 ( .A1(n90564), .A2(n90565), .A3(n90566), .A4(n90567), .ZN(
        n90563) );
  NAND2_X1 U76110 ( .A1(n90568), .A2(n90569), .ZN(n90567) );
  AOI22_X1 U76111 ( .A1(n90325), .A2(n108018), .B1(n90326), .B2(n108019), .ZN(
        n90569) );
  AOI22_X1 U76112 ( .A1(n90327), .A2(n108027), .B1(n90328), .B2(n108025), .ZN(
        n90568) );
  NAND2_X1 U76113 ( .A1(n90570), .A2(n90571), .ZN(n90566) );
  AOI22_X1 U76114 ( .A1(n90331), .A2(n70433), .B1(n90332), .B2(n108022), .ZN(
        n90571) );
  AOI22_X1 U76115 ( .A1(n90333), .A2(n70537), .B1(n90334), .B2(n107952), .ZN(
        n90570) );
  NAND2_X1 U76116 ( .A1(n90572), .A2(n90573), .ZN(n90565) );
  AOI22_X1 U76117 ( .A1(n90337), .A2(n107956), .B1(n90338), .B2(n70437), .ZN(
        n90573) );
  AOI22_X1 U76118 ( .A1(n90339), .A2(n108023), .B1(n90340), .B2(n108020), .ZN(
        n90572) );
  NAND2_X1 U76119 ( .A1(n90574), .A2(n90575), .ZN(n90564) );
  AOI22_X1 U76120 ( .A1(n90343), .A2(n107954), .B1(n90344), .B2(n107958), .ZN(
        n90575) );
  AOI22_X1 U76121 ( .A1(n90345), .A2(n107957), .B1(n90346), .B2(n70439), .ZN(
        n90574) );
  NOR4_X1 U76122 ( .A1(n90576), .A2(n90577), .A3(n90578), .A4(n90579), .ZN(
        n90562) );
  NAND2_X1 U76123 ( .A1(n90580), .A2(n90581), .ZN(n90579) );
  AOI22_X1 U76124 ( .A1(n90353), .A2(n108028), .B1(n90354), .B2(n108031), .ZN(
        n90581) );
  AOI22_X1 U76125 ( .A1(n90355), .A2(n108032), .B1(n90356), .B2(n108034), .ZN(
        n90580) );
  NAND2_X1 U76126 ( .A1(n90582), .A2(n90583), .ZN(n90578) );
  AOI22_X1 U76127 ( .A1(n90359), .A2(n108033), .B1(n90360), .B2(n108029), .ZN(
        n90583) );
  AOI22_X1 U76128 ( .A1(n90361), .A2(n108035), .B1(n90362), .B2(n108030), .ZN(
        n90582) );
  NAND2_X1 U76129 ( .A1(n90584), .A2(n90585), .ZN(n90577) );
  AOI22_X1 U76130 ( .A1(n90365), .A2(n70547), .B1(n90366), .B2(n70546), .ZN(
        n90585) );
  AOI22_X1 U76131 ( .A1(n90367), .A2(n70549), .B1(n90368), .B2(n108036), .ZN(
        n90584) );
  NAND2_X1 U76132 ( .A1(n90586), .A2(n90587), .ZN(n90576) );
  AOI22_X1 U76133 ( .A1(n90371), .A2(n108021), .B1(n90372), .B2(n108026), .ZN(
        n90587) );
  AOI22_X1 U76134 ( .A1(n90373), .A2(n70544), .B1(n90374), .B2(n108024), .ZN(
        n90586) );
  NAND2_X1 U76135 ( .A1(n90588), .A2(n90589), .ZN(n90560) );
  NOR4_X1 U76136 ( .A1(n90590), .A2(n90591), .A3(n90592), .A4(n90593), .ZN(
        n90589) );
  NAND2_X1 U76137 ( .A1(n90594), .A2(n90595), .ZN(n90593) );
  AOI22_X1 U76138 ( .A1(n90383), .A2(n107966), .B1(n90384), .B2(n107968), .ZN(
        n90595) );
  AOI22_X1 U76139 ( .A1(n90385), .A2(n70462), .B1(n90386), .B2(n107967), .ZN(
        n90594) );
  NAND2_X1 U76140 ( .A1(n90596), .A2(n90597), .ZN(n90592) );
  AOI22_X1 U76141 ( .A1(n90389), .A2(n70466), .B1(n90390), .B2(n70468), .ZN(
        n90597) );
  AOI22_X1 U76142 ( .A1(n90391), .A2(n107972), .B1(n90392), .B2(n107973), .ZN(
        n90596) );
  NAND2_X1 U76143 ( .A1(n90598), .A2(n90599), .ZN(n90591) );
  AOI22_X1 U76144 ( .A1(n90395), .A2(n107971), .B1(n90396), .B2(n70463), .ZN(
        n90599) );
  AOI22_X1 U76145 ( .A1(n90397), .A2(n107974), .B1(n90398), .B2(n70461), .ZN(
        n90598) );
  NAND2_X1 U76146 ( .A1(n90600), .A2(n90601), .ZN(n90590) );
  AOI22_X1 U76147 ( .A1(n90401), .A2(n107976), .B1(n90402), .B2(n70473), .ZN(
        n90601) );
  AOI22_X1 U76148 ( .A1(n90403), .A2(n70474), .B1(n90404), .B2(n70471), .ZN(
        n90600) );
  NOR4_X1 U76149 ( .A1(n90602), .A2(n90603), .A3(n90604), .A4(n90605), .ZN(
        n90588) );
  NAND2_X1 U76150 ( .A1(n90606), .A2(n90607), .ZN(n90605) );
  AOI22_X1 U76151 ( .A1(n90411), .A2(n107961), .B1(n90412), .B2(n107953), .ZN(
        n90607) );
  AOI22_X1 U76152 ( .A1(n90413), .A2(n107955), .B1(n90414), .B2(n70445), .ZN(
        n90606) );
  NAND2_X1 U76153 ( .A1(n90608), .A2(n90609), .ZN(n90604) );
  AOI22_X1 U76154 ( .A1(n90417), .A2(n107960), .B1(n90418), .B2(n107963), .ZN(
        n90609) );
  AOI22_X1 U76155 ( .A1(n90419), .A2(n107965), .B1(n90420), .B2(n107962), .ZN(
        n90608) );
  NAND2_X1 U76156 ( .A1(n90610), .A2(n90611), .ZN(n90603) );
  AOI22_X1 U76157 ( .A1(n90423), .A2(n70454), .B1(n90424), .B2(n107959), .ZN(
        n90611) );
  AOI22_X1 U76158 ( .A1(n90425), .A2(n70446), .B1(n90426), .B2(n70450), .ZN(
        n90610) );
  NAND2_X1 U76159 ( .A1(n90612), .A2(n90613), .ZN(n90602) );
  AOI22_X1 U76160 ( .A1(n90429), .A2(n107970), .B1(n90430), .B2(n70458), .ZN(
        n90613) );
  AOI22_X1 U76161 ( .A1(n90431), .A2(n70456), .B1(n90432), .B2(n107969), .ZN(
        n90612) );
  NAND2_X1 U76162 ( .A1(n90614), .A2(n90615), .ZN(n90559) );
  NOR4_X1 U76163 ( .A1(n90616), .A2(n90617), .A3(n90618), .A4(n90619), .ZN(
        n90615) );
  NAND2_X1 U76164 ( .A1(n90620), .A2(n90621), .ZN(n90619) );
  AOI22_X1 U76165 ( .A1(n90441), .A2(n70496), .B1(n90442), .B2(n107985), .ZN(
        n90621) );
  AOI22_X1 U76166 ( .A1(n90443), .A2(n107988), .B1(n90444), .B2(n70492), .ZN(
        n90620) );
  NAND2_X1 U76167 ( .A1(n90622), .A2(n90623), .ZN(n90618) );
  AOI22_X1 U76168 ( .A1(n90447), .A2(n107991), .B1(n90448), .B2(n107990), .ZN(
        n90623) );
  AOI22_X1 U76169 ( .A1(n90449), .A2(n107984), .B1(n90450), .B2(n107986), .ZN(
        n90622) );
  NAND2_X1 U76170 ( .A1(n90624), .A2(n90625), .ZN(n90617) );
  AOI22_X1 U76171 ( .A1(n90453), .A2(n107992), .B1(n90454), .B2(n107989), .ZN(
        n90625) );
  AOI22_X1 U76172 ( .A1(n90455), .A2(n70500), .B1(n90456), .B2(n70502), .ZN(
        n90624) );
  NAND2_X1 U76173 ( .A1(n90626), .A2(n90627), .ZN(n90616) );
  AOI22_X1 U76174 ( .A1(n90459), .A2(n107995), .B1(n90460), .B2(n70508), .ZN(
        n90627) );
  AOI22_X1 U76175 ( .A1(n90461), .A2(n70494), .B1(n90462), .B2(n70497), .ZN(
        n90626) );
  NOR4_X1 U76176 ( .A1(n90628), .A2(n90629), .A3(n90630), .A4(n90631), .ZN(
        n90614) );
  NAND2_X1 U76177 ( .A1(n90632), .A2(n90633), .ZN(n90631) );
  AOI22_X1 U76178 ( .A1(n90469), .A2(n70472), .B1(n90470), .B2(n107979), .ZN(
        n90633) );
  AOI22_X1 U76179 ( .A1(n90471), .A2(n70470), .B1(n90472), .B2(n70476), .ZN(
        n90632) );
  NAND2_X1 U76180 ( .A1(n90634), .A2(n90635), .ZN(n90630) );
  AOI22_X1 U76181 ( .A1(n90475), .A2(n70485), .B1(n90476), .B2(n107981), .ZN(
        n90635) );
  AOI22_X1 U76182 ( .A1(n90477), .A2(n107982), .B1(n90478), .B2(n107975), .ZN(
        n90634) );
  NAND2_X1 U76183 ( .A1(n90636), .A2(n90637), .ZN(n90629) );
  AOI22_X1 U76184 ( .A1(n90481), .A2(n107980), .B1(n90482), .B2(n70484), .ZN(
        n90637) );
  AOI22_X1 U76185 ( .A1(n90483), .A2(n107978), .B1(n90484), .B2(n107983), .ZN(
        n90636) );
  NAND2_X1 U76186 ( .A1(n90638), .A2(n90639), .ZN(n90628) );
  AOI22_X1 U76187 ( .A1(n90487), .A2(n70490), .B1(n90488), .B2(n107987), .ZN(
        n90639) );
  AOI22_X1 U76188 ( .A1(n90489), .A2(n70488), .B1(n90490), .B2(n107977), .ZN(
        n90638) );
  NAND2_X1 U76189 ( .A1(n90640), .A2(n90641), .ZN(n90558) );
  NOR4_X1 U76190 ( .A1(n90642), .A2(n90643), .A3(n90644), .A4(n90645), .ZN(
        n90641) );
  NAND2_X1 U76191 ( .A1(n90646), .A2(n90647), .ZN(n90645) );
  AOI22_X1 U76192 ( .A1(n90499), .A2(n108010), .B1(n90500), .B2(n108009), .ZN(
        n90647) );
  AOI22_X1 U76193 ( .A1(n90501), .A2(n70524), .B1(n90502), .B2(n108007), .ZN(
        n90646) );
  NAND2_X1 U76194 ( .A1(n90648), .A2(n90649), .ZN(n90644) );
  AOI22_X1 U76195 ( .A1(n90505), .A2(n108005), .B1(n90506), .B2(n108008), .ZN(
        n90649) );
  AOI22_X1 U76196 ( .A1(n90507), .A2(n70530), .B1(n90508), .B2(n108006), .ZN(
        n90648) );
  NAND2_X1 U76197 ( .A1(n90650), .A2(n90651), .ZN(n90643) );
  AOI22_X1 U76198 ( .A1(n105650), .A2(n108016), .B1(n90512), .B2(n70536), .ZN(
        n90651) );
  AOI22_X1 U76199 ( .A1(n90513), .A2(n108014), .B1(n90514), .B2(n108015), .ZN(
        n90650) );
  NAND2_X1 U76200 ( .A1(n90652), .A2(n90653), .ZN(n90642) );
  AOI22_X1 U76201 ( .A1(n90517), .A2(n108011), .B1(n90518), .B2(n108013), .ZN(
        n90653) );
  AOI22_X1 U76202 ( .A1(n90519), .A2(n70535), .B1(n105644), .B2(n108012), .ZN(
        n90652) );
  NOR4_X1 U76203 ( .A1(n90654), .A2(n90655), .A3(n90656), .A4(n90657), .ZN(
        n90640) );
  NAND2_X1 U76204 ( .A1(n90658), .A2(n90659), .ZN(n90657) );
  AOI22_X1 U76205 ( .A1(n90527), .A2(n107994), .B1(n90528), .B2(n107997), .ZN(
        n90659) );
  AOI22_X1 U76206 ( .A1(n90529), .A2(n107996), .B1(n90530), .B2(n70507), .ZN(
        n90658) );
  NAND2_X1 U76207 ( .A1(n90660), .A2(n90661), .ZN(n90656) );
  AOI22_X1 U76208 ( .A1(n90533), .A2(n108002), .B1(n90534), .B2(n107993), .ZN(
        n90661) );
  AOI22_X1 U76209 ( .A1(n90535), .A2(n70506), .B1(n90536), .B2(n107999), .ZN(
        n90660) );
  NAND2_X1 U76210 ( .A1(n90662), .A2(n90663), .ZN(n90655) );
  AOI22_X1 U76211 ( .A1(n90539), .A2(n107998), .B1(n90540), .B2(n108003), .ZN(
        n90663) );
  AOI22_X1 U76212 ( .A1(n90541), .A2(n108004), .B1(n90542), .B2(n108001), .ZN(
        n90662) );
  NAND2_X1 U76213 ( .A1(n90664), .A2(n90665), .ZN(n90654) );
  AOI22_X1 U76214 ( .A1(n90545), .A2(n70525), .B1(n90546), .B2(n70511), .ZN(
        n90665) );
  AOI22_X1 U76215 ( .A1(n90547), .A2(n70514), .B1(n90548), .B2(n70518), .ZN(
        n90664) );
  AOI21_X1 U76216 ( .B1(n90295), .B2(n86676), .A(n90667), .ZN(n90666) );
  OAI21_X1 U76217 ( .B1(n90668), .B2(n105659), .A(n90669), .ZN(n90667) );
  OAI21_X1 U76218 ( .B1(n90670), .B2(n90671), .A(n90302), .ZN(n90669) );
  OAI21_X1 U76219 ( .B1(n102150), .B2(n90303), .A(n90672), .ZN(n90671) );
  AOI22_X1 U76220 ( .A1(n90305), .A2(n107174), .B1(n90306), .B2(n69425), .ZN(
        n90672) );
  NAND2_X1 U76221 ( .A1(n90673), .A2(n90674), .ZN(n90670) );
  AOI22_X1 U76222 ( .A1(n90309), .A2(n106838), .B1(n105653), .B2(n107170), 
        .ZN(n90674) );
  AOI22_X1 U76223 ( .A1(n90311), .A2(n69429), .B1(n90312), .B2(n107172), .ZN(
        n90673) );
  NOR4_X1 U76224 ( .A1(n90675), .A2(n90676), .A3(n90677), .A4(n90678), .ZN(
        n90668) );
  NAND2_X1 U76225 ( .A1(n90679), .A2(n90680), .ZN(n90678) );
  NOR4_X1 U76226 ( .A1(n90681), .A2(n90682), .A3(n90683), .A4(n90684), .ZN(
        n90680) );
  NAND2_X1 U76227 ( .A1(n90685), .A2(n90686), .ZN(n90684) );
  AOI22_X1 U76228 ( .A1(n90325), .A2(n107212), .B1(n90326), .B2(n107210), .ZN(
        n90686) );
  AOI22_X1 U76229 ( .A1(n90327), .A2(n107194), .B1(n90328), .B2(n107198), .ZN(
        n90685) );
  NAND2_X1 U76230 ( .A1(n90687), .A2(n90688), .ZN(n90683) );
  AOI22_X1 U76231 ( .A1(n90331), .A2(n69486), .B1(n90332), .B2(n107204), .ZN(
        n90688) );
  AOI22_X1 U76232 ( .A1(n90333), .A2(n69483), .B1(n90334), .B2(n107214), .ZN(
        n90687) );
  NAND2_X1 U76233 ( .A1(n90689), .A2(n90690), .ZN(n90682) );
  AOI22_X1 U76234 ( .A1(n90337), .A2(n107218), .B1(n90338), .B2(n69490), .ZN(
        n90690) );
  AOI22_X1 U76235 ( .A1(n90339), .A2(n107202), .B1(n90340), .B2(n107208), .ZN(
        n90689) );
  NAND2_X1 U76236 ( .A1(n90691), .A2(n90692), .ZN(n90681) );
  AOI22_X1 U76237 ( .A1(n90343), .A2(n107216), .B1(n90344), .B2(n107220), .ZN(
        n90692) );
  AOI22_X1 U76238 ( .A1(n90345), .A2(n107219), .B1(n90346), .B2(n69492), .ZN(
        n90691) );
  NOR4_X1 U76239 ( .A1(n90693), .A2(n90694), .A3(n90695), .A4(n90696), .ZN(
        n90679) );
  NAND2_X1 U76240 ( .A1(n90697), .A2(n90698), .ZN(n90696) );
  AOI22_X1 U76241 ( .A1(n90353), .A2(n107192), .B1(n90354), .B2(n107186), .ZN(
        n90698) );
  AOI22_X1 U76242 ( .A1(n90355), .A2(n107184), .B1(n90356), .B2(n107180), .ZN(
        n90697) );
  NAND2_X1 U76243 ( .A1(n90699), .A2(n90700), .ZN(n90695) );
  AOI22_X1 U76244 ( .A1(n90359), .A2(n107182), .B1(n90360), .B2(n107190), .ZN(
        n90700) );
  AOI22_X1 U76245 ( .A1(n90361), .A2(n107178), .B1(n90362), .B2(n107188), .ZN(
        n90699) );
  NAND2_X1 U76246 ( .A1(n90701), .A2(n90702), .ZN(n90694) );
  AOI22_X1 U76247 ( .A1(n90365), .A2(n69463), .B1(n90366), .B2(n69465), .ZN(
        n90702) );
  AOI22_X1 U76248 ( .A1(n90367), .A2(n69459), .B1(n90368), .B2(n107176), .ZN(
        n90701) );
  NAND2_X1 U76249 ( .A1(n90703), .A2(n90704), .ZN(n90693) );
  AOI22_X1 U76250 ( .A1(n90371), .A2(n107206), .B1(n90372), .B2(n107196), .ZN(
        n90704) );
  AOI22_X1 U76251 ( .A1(n90373), .A2(n69469), .B1(n90374), .B2(n107200), .ZN(
        n90703) );
  NAND2_X1 U76252 ( .A1(n90705), .A2(n90706), .ZN(n90677) );
  NOR4_X1 U76253 ( .A1(n90707), .A2(n90708), .A3(n90709), .A4(n90710), .ZN(
        n90706) );
  NAND2_X1 U76254 ( .A1(n90711), .A2(n90712), .ZN(n90710) );
  AOI22_X1 U76255 ( .A1(n90383), .A2(n107229), .B1(n90384), .B2(n107231), .ZN(
        n90712) );
  AOI22_X1 U76256 ( .A1(n90385), .A2(n69515), .B1(n90386), .B2(n107230), .ZN(
        n90711) );
  NAND2_X1 U76257 ( .A1(n90713), .A2(n90714), .ZN(n90709) );
  AOI22_X1 U76258 ( .A1(n90389), .A2(n69519), .B1(n90390), .B2(n69521), .ZN(
        n90714) );
  AOI22_X1 U76259 ( .A1(n90391), .A2(n107236), .B1(n90392), .B2(n107237), .ZN(
        n90713) );
  NAND2_X1 U76260 ( .A1(n90715), .A2(n90716), .ZN(n90708) );
  AOI22_X1 U76261 ( .A1(n90395), .A2(n107234), .B1(n90396), .B2(n107235), .ZN(
        n90716) );
  AOI22_X1 U76262 ( .A1(n90397), .A2(n107238), .B1(n90398), .B2(n69514), .ZN(
        n90715) );
  NAND2_X1 U76263 ( .A1(n90717), .A2(n90718), .ZN(n90707) );
  AOI22_X1 U76264 ( .A1(n90401), .A2(n107243), .B1(n90402), .B2(n69526), .ZN(
        n90718) );
  AOI22_X1 U76265 ( .A1(n90403), .A2(n107242), .B1(n90404), .B2(n69524), .ZN(
        n90717) );
  NOR4_X1 U76266 ( .A1(n90719), .A2(n90720), .A3(n90721), .A4(n90722), .ZN(
        n90705) );
  NAND2_X1 U76267 ( .A1(n90723), .A2(n90724), .ZN(n90722) );
  AOI22_X1 U76268 ( .A1(n90411), .A2(n107224), .B1(n90412), .B2(n107215), .ZN(
        n90724) );
  AOI22_X1 U76269 ( .A1(n90413), .A2(n107217), .B1(n90414), .B2(n69498), .ZN(
        n90723) );
  NAND2_X1 U76270 ( .A1(n90725), .A2(n90726), .ZN(n90721) );
  AOI22_X1 U76271 ( .A1(n90417), .A2(n107222), .B1(n90418), .B2(n107226), .ZN(
        n90726) );
  AOI22_X1 U76272 ( .A1(n90419), .A2(n107228), .B1(n90420), .B2(n107225), .ZN(
        n90725) );
  NAND2_X1 U76273 ( .A1(n90727), .A2(n90728), .ZN(n90720) );
  AOI22_X1 U76274 ( .A1(n90423), .A2(n69507), .B1(n90424), .B2(n107221), .ZN(
        n90728) );
  AOI22_X1 U76275 ( .A1(n90425), .A2(n107223), .B1(n90426), .B2(n69503), .ZN(
        n90727) );
  NAND2_X1 U76276 ( .A1(n90729), .A2(n90730), .ZN(n90719) );
  AOI22_X1 U76277 ( .A1(n90429), .A2(n107233), .B1(n90430), .B2(n69511), .ZN(
        n90730) );
  AOI22_X1 U76278 ( .A1(n90431), .A2(n69509), .B1(n90432), .B2(n107232), .ZN(
        n90729) );
  NAND2_X1 U76279 ( .A1(n90731), .A2(n90732), .ZN(n90676) );
  NOR4_X1 U76280 ( .A1(n90733), .A2(n90734), .A3(n90735), .A4(n90736), .ZN(
        n90732) );
  NAND2_X1 U76281 ( .A1(n90737), .A2(n90738), .ZN(n90736) );
  AOI22_X1 U76282 ( .A1(n90441), .A2(n69549), .B1(n90442), .B2(n107253), .ZN(
        n90738) );
  AOI22_X1 U76283 ( .A1(n90443), .A2(n107256), .B1(n90444), .B2(n69545), .ZN(
        n90737) );
  NAND2_X1 U76284 ( .A1(n90739), .A2(n90740), .ZN(n90735) );
  AOI22_X1 U76285 ( .A1(n90447), .A2(n107261), .B1(n90448), .B2(n107260), .ZN(
        n90740) );
  AOI22_X1 U76286 ( .A1(n90449), .A2(n107252), .B1(n90450), .B2(n107254), .ZN(
        n90739) );
  NAND2_X1 U76287 ( .A1(n90741), .A2(n90742), .ZN(n90734) );
  AOI22_X1 U76288 ( .A1(n90453), .A2(n107262), .B1(n90454), .B2(n107258), .ZN(
        n90742) );
  AOI22_X1 U76289 ( .A1(n90455), .A2(n69553), .B1(n90456), .B2(n69555), .ZN(
        n90741) );
  NAND2_X1 U76290 ( .A1(n90743), .A2(n90744), .ZN(n90733) );
  AOI22_X1 U76291 ( .A1(n90459), .A2(n107265), .B1(n90460), .B2(n69561), .ZN(
        n90744) );
  AOI22_X1 U76292 ( .A1(n90461), .A2(n107257), .B1(n90462), .B2(n107259), .ZN(
        n90743) );
  NOR4_X1 U76293 ( .A1(n90745), .A2(n90746), .A3(n90747), .A4(n90748), .ZN(
        n90731) );
  NAND2_X1 U76294 ( .A1(n90749), .A2(n90750), .ZN(n90748) );
  AOI22_X1 U76295 ( .A1(n90469), .A2(n107241), .B1(n90470), .B2(n107246), .ZN(
        n90750) );
  AOI22_X1 U76296 ( .A1(n90471), .A2(n107240), .B1(n90472), .B2(n69529), .ZN(
        n90749) );
  NAND2_X1 U76297 ( .A1(n90751), .A2(n90752), .ZN(n90747) );
  AOI22_X1 U76298 ( .A1(n90475), .A2(n69538), .B1(n90476), .B2(n107248), .ZN(
        n90752) );
  AOI22_X1 U76299 ( .A1(n90477), .A2(n107249), .B1(n90478), .B2(n107239), .ZN(
        n90751) );
  NAND2_X1 U76300 ( .A1(n90753), .A2(n90754), .ZN(n90746) );
  AOI22_X1 U76301 ( .A1(n90481), .A2(n107247), .B1(n90482), .B2(n107251), .ZN(
        n90754) );
  AOI22_X1 U76302 ( .A1(n90483), .A2(n107245), .B1(n90484), .B2(n107250), .ZN(
        n90753) );
  NAND2_X1 U76303 ( .A1(n90755), .A2(n90756), .ZN(n90745) );
  AOI22_X1 U76304 ( .A1(n90487), .A2(n69543), .B1(n90488), .B2(n107255), .ZN(
        n90756) );
  AOI22_X1 U76305 ( .A1(n90489), .A2(n69541), .B1(n90490), .B2(n107244), .ZN(
        n90755) );
  NAND2_X1 U76306 ( .A1(n90757), .A2(n90758), .ZN(n90675) );
  NOR4_X1 U76307 ( .A1(n90759), .A2(n90760), .A3(n90761), .A4(n90762), .ZN(
        n90758) );
  NAND2_X1 U76308 ( .A1(n90763), .A2(n90764), .ZN(n90762) );
  AOI22_X1 U76309 ( .A1(n90499), .A2(n107281), .B1(n90500), .B2(n107280), .ZN(
        n90764) );
  AOI22_X1 U76310 ( .A1(n90501), .A2(n69577), .B1(n90502), .B2(n107278), .ZN(
        n90763) );
  NAND2_X1 U76311 ( .A1(n90765), .A2(n90766), .ZN(n90761) );
  AOI22_X1 U76312 ( .A1(n90505), .A2(n107276), .B1(n90506), .B2(n107279), .ZN(
        n90766) );
  AOI22_X1 U76313 ( .A1(n90507), .A2(n69583), .B1(n90508), .B2(n107277), .ZN(
        n90765) );
  NAND2_X1 U76314 ( .A1(n90767), .A2(n90768), .ZN(n90760) );
  AOI22_X1 U76315 ( .A1(n105650), .A2(n107286), .B1(n90512), .B2(n69589), .ZN(
        n90768) );
  AOI22_X1 U76316 ( .A1(n90513), .A2(n107284), .B1(n90514), .B2(n107285), .ZN(
        n90767) );
  NAND2_X1 U76317 ( .A1(n90769), .A2(n90770), .ZN(n90759) );
  AOI22_X1 U76318 ( .A1(n90517), .A2(n69581), .B1(n90518), .B2(n107283), .ZN(
        n90770) );
  AOI22_X1 U76319 ( .A1(n90519), .A2(n69588), .B1(n105644), .B2(n107282), .ZN(
        n90769) );
  NOR4_X1 U76320 ( .A1(n90771), .A2(n90772), .A3(n90773), .A4(n90774), .ZN(
        n90757) );
  NAND2_X1 U76321 ( .A1(n90775), .A2(n90776), .ZN(n90774) );
  AOI22_X1 U76322 ( .A1(n90527), .A2(n107264), .B1(n90528), .B2(n107268), .ZN(
        n90776) );
  AOI22_X1 U76323 ( .A1(n90529), .A2(n107267), .B1(n90530), .B2(n69560), .ZN(
        n90775) );
  NAND2_X1 U76324 ( .A1(n90777), .A2(n90778), .ZN(n90773) );
  AOI22_X1 U76325 ( .A1(n90533), .A2(n107273), .B1(n90534), .B2(n107263), .ZN(
        n90778) );
  AOI22_X1 U76326 ( .A1(n90535), .A2(n107266), .B1(n90536), .B2(n107270), .ZN(
        n90777) );
  NAND2_X1 U76327 ( .A1(n90779), .A2(n90780), .ZN(n90772) );
  AOI22_X1 U76328 ( .A1(n90539), .A2(n107269), .B1(n90540), .B2(n107274), .ZN(
        n90780) );
  AOI22_X1 U76329 ( .A1(n90541), .A2(n107275), .B1(n90542), .B2(n107272), .ZN(
        n90779) );
  NAND2_X1 U76330 ( .A1(n90781), .A2(n90782), .ZN(n90771) );
  AOI22_X1 U76331 ( .A1(n90545), .A2(n69578), .B1(n90546), .B2(n69564), .ZN(
        n90782) );
  AOI22_X1 U76332 ( .A1(n90547), .A2(n69567), .B1(n90548), .B2(n69571), .ZN(
        n90781) );
  AOI21_X1 U76333 ( .B1(n90295), .B2(n86794), .A(n90784), .ZN(n90783) );
  OAI21_X1 U76334 ( .B1(n90785), .B2(n105659), .A(n90786), .ZN(n90784) );
  OAI21_X1 U76335 ( .B1(n90787), .B2(n90788), .A(n90302), .ZN(n90786) );
  OAI21_X1 U76336 ( .B1(n102134), .B2(n90303), .A(n90789), .ZN(n90788) );
  AOI22_X1 U76337 ( .A1(n90305), .A2(n107846), .B1(n90306), .B2(n70280), .ZN(
        n90789) );
  NAND2_X1 U76338 ( .A1(n90790), .A2(n90791), .ZN(n90787) );
  AOI22_X1 U76339 ( .A1(n90309), .A2(n107851), .B1(n105653), .B2(n107848), 
        .ZN(n90791) );
  AOI22_X1 U76340 ( .A1(n90311), .A2(n70278), .B1(n90312), .B2(n107847), .ZN(
        n90790) );
  NOR4_X1 U76341 ( .A1(n90792), .A2(n90793), .A3(n90794), .A4(n90795), .ZN(
        n90785) );
  NAND2_X1 U76342 ( .A1(n90796), .A2(n90797), .ZN(n90795) );
  NOR4_X1 U76343 ( .A1(n90798), .A2(n90799), .A3(n90800), .A4(n90801), .ZN(
        n90797) );
  NAND2_X1 U76344 ( .A1(n90802), .A2(n90803), .ZN(n90801) );
  AOI22_X1 U76345 ( .A1(n90325), .A2(n107826), .B1(n90326), .B2(n107827), .ZN(
        n90803) );
  AOI22_X1 U76346 ( .A1(n90327), .A2(n107836), .B1(n90328), .B2(n107834), .ZN(
        n90802) );
  NAND2_X1 U76347 ( .A1(n90804), .A2(n90805), .ZN(n90800) );
  AOI22_X1 U76348 ( .A1(n90331), .A2(n70147), .B1(n90332), .B2(n107830), .ZN(
        n90805) );
  AOI22_X1 U76349 ( .A1(n90333), .A2(n70251), .B1(n90334), .B2(n107752), .ZN(
        n90804) );
  NAND2_X1 U76350 ( .A1(n90806), .A2(n90807), .ZN(n90799) );
  AOI22_X1 U76351 ( .A1(n90337), .A2(n107756), .B1(n90338), .B2(n70151), .ZN(
        n90807) );
  AOI22_X1 U76352 ( .A1(n90339), .A2(n107831), .B1(n90340), .B2(n107828), .ZN(
        n90806) );
  NAND2_X1 U76353 ( .A1(n90808), .A2(n90809), .ZN(n90798) );
  AOI22_X1 U76354 ( .A1(n90343), .A2(n107754), .B1(n90344), .B2(n107758), .ZN(
        n90809) );
  AOI22_X1 U76355 ( .A1(n90345), .A2(n107757), .B1(n90346), .B2(n70153), .ZN(
        n90808) );
  NOR4_X1 U76356 ( .A1(n90810), .A2(n90811), .A3(n90812), .A4(n90813), .ZN(
        n90796) );
  NAND2_X1 U76357 ( .A1(n90814), .A2(n90815), .ZN(n90813) );
  AOI22_X1 U76358 ( .A1(n90353), .A2(n107837), .B1(n90354), .B2(n107840), .ZN(
        n90815) );
  AOI22_X1 U76359 ( .A1(n90355), .A2(n107841), .B1(n90356), .B2(n107843), .ZN(
        n90814) );
  NAND2_X1 U76360 ( .A1(n90816), .A2(n90817), .ZN(n90812) );
  AOI22_X1 U76361 ( .A1(n90359), .A2(n107842), .B1(n90360), .B2(n107838), .ZN(
        n90817) );
  AOI22_X1 U76362 ( .A1(n90361), .A2(n107844), .B1(n90362), .B2(n107839), .ZN(
        n90816) );
  NAND2_X1 U76363 ( .A1(n90818), .A2(n90819), .ZN(n90811) );
  AOI22_X1 U76364 ( .A1(n90365), .A2(n70261), .B1(n90366), .B2(n70260), .ZN(
        n90819) );
  AOI22_X1 U76365 ( .A1(n90367), .A2(n70263), .B1(n90368), .B2(n107845), .ZN(
        n90818) );
  NAND2_X1 U76366 ( .A1(n90820), .A2(n90821), .ZN(n90810) );
  AOI22_X1 U76367 ( .A1(n90371), .A2(n107829), .B1(n90372), .B2(n107835), .ZN(
        n90821) );
  AOI22_X1 U76368 ( .A1(n90373), .A2(n70258), .B1(n90374), .B2(n107833), .ZN(
        n90820) );
  NAND2_X1 U76369 ( .A1(n90822), .A2(n90823), .ZN(n90794) );
  NOR4_X1 U76370 ( .A1(n90824), .A2(n90825), .A3(n90826), .A4(n90827), .ZN(
        n90823) );
  NAND2_X1 U76371 ( .A1(n90828), .A2(n90829), .ZN(n90827) );
  AOI22_X1 U76372 ( .A1(n90383), .A2(n107767), .B1(n90384), .B2(n107769), .ZN(
        n90829) );
  AOI22_X1 U76373 ( .A1(n90385), .A2(n70176), .B1(n90386), .B2(n107768), .ZN(
        n90828) );
  NAND2_X1 U76374 ( .A1(n90830), .A2(n90831), .ZN(n90826) );
  AOI22_X1 U76375 ( .A1(n90389), .A2(n70180), .B1(n90390), .B2(n70182), .ZN(
        n90831) );
  AOI22_X1 U76376 ( .A1(n90391), .A2(n107775), .B1(n90392), .B2(n107776), .ZN(
        n90830) );
  NAND2_X1 U76377 ( .A1(n90832), .A2(n90833), .ZN(n90825) );
  AOI22_X1 U76378 ( .A1(n90395), .A2(n107772), .B1(n90396), .B2(n107774), .ZN(
        n90833) );
  AOI22_X1 U76379 ( .A1(n90397), .A2(n107777), .B1(n90398), .B2(n107773), .ZN(
        n90832) );
  NAND2_X1 U76380 ( .A1(n90834), .A2(n90835), .ZN(n90824) );
  AOI22_X1 U76381 ( .A1(n90401), .A2(n107782), .B1(n90402), .B2(n70187), .ZN(
        n90835) );
  AOI22_X1 U76382 ( .A1(n90403), .A2(n107781), .B1(n90404), .B2(n70185), .ZN(
        n90834) );
  NOR4_X1 U76383 ( .A1(n90836), .A2(n90837), .A3(n90838), .A4(n90839), .ZN(
        n90822) );
  NAND2_X1 U76384 ( .A1(n90840), .A2(n90841), .ZN(n90839) );
  AOI22_X1 U76385 ( .A1(n90411), .A2(n107762), .B1(n90412), .B2(n107753), .ZN(
        n90841) );
  AOI22_X1 U76386 ( .A1(n90413), .A2(n107755), .B1(n90414), .B2(n70159), .ZN(
        n90840) );
  NAND2_X1 U76387 ( .A1(n90842), .A2(n90843), .ZN(n90838) );
  AOI22_X1 U76388 ( .A1(n90417), .A2(n107760), .B1(n90418), .B2(n107764), .ZN(
        n90843) );
  AOI22_X1 U76389 ( .A1(n90419), .A2(n107766), .B1(n90420), .B2(n107763), .ZN(
        n90842) );
  NAND2_X1 U76390 ( .A1(n90844), .A2(n90845), .ZN(n90837) );
  AOI22_X1 U76391 ( .A1(n90423), .A2(n70168), .B1(n90424), .B2(n107759), .ZN(
        n90845) );
  AOI22_X1 U76392 ( .A1(n90425), .A2(n107761), .B1(n90426), .B2(n107765), .ZN(
        n90844) );
  NAND2_X1 U76393 ( .A1(n90846), .A2(n90847), .ZN(n90836) );
  AOI22_X1 U76394 ( .A1(n90429), .A2(n107771), .B1(n90430), .B2(n70172), .ZN(
        n90847) );
  AOI22_X1 U76395 ( .A1(n90431), .A2(n70170), .B1(n90432), .B2(n107770), .ZN(
        n90846) );
  NAND2_X1 U76396 ( .A1(n90848), .A2(n90849), .ZN(n90793) );
  NOR4_X1 U76397 ( .A1(n90850), .A2(n90851), .A3(n90852), .A4(n90853), .ZN(
        n90849) );
  NAND2_X1 U76398 ( .A1(n90854), .A2(n90855), .ZN(n90853) );
  AOI22_X1 U76399 ( .A1(n90441), .A2(n70210), .B1(n90442), .B2(n107792), .ZN(
        n90855) );
  AOI22_X1 U76400 ( .A1(n90443), .A2(n107795), .B1(n90444), .B2(n70206), .ZN(
        n90854) );
  NAND2_X1 U76401 ( .A1(n90856), .A2(n90857), .ZN(n90852) );
  AOI22_X1 U76402 ( .A1(n90447), .A2(n107798), .B1(n90448), .B2(n107797), .ZN(
        n90857) );
  AOI22_X1 U76403 ( .A1(n90449), .A2(n107791), .B1(n90450), .B2(n107793), .ZN(
        n90856) );
  NAND2_X1 U76404 ( .A1(n90858), .A2(n90859), .ZN(n90851) );
  AOI22_X1 U76405 ( .A1(n90453), .A2(n107799), .B1(n90454), .B2(n70209), .ZN(
        n90859) );
  AOI22_X1 U76406 ( .A1(n90455), .A2(n70214), .B1(n90456), .B2(n70216), .ZN(
        n90858) );
  NAND2_X1 U76407 ( .A1(n90860), .A2(n90861), .ZN(n90850) );
  AOI22_X1 U76408 ( .A1(n90459), .A2(n107802), .B1(n90460), .B2(n70222), .ZN(
        n90861) );
  AOI22_X1 U76409 ( .A1(n90461), .A2(n70208), .B1(n90462), .B2(n107796), .ZN(
        n90860) );
  NOR4_X1 U76410 ( .A1(n90862), .A2(n90863), .A3(n90864), .A4(n90865), .ZN(
        n90848) );
  NAND2_X1 U76411 ( .A1(n90866), .A2(n90867), .ZN(n90865) );
  AOI22_X1 U76412 ( .A1(n90469), .A2(n107780), .B1(n90470), .B2(n107785), .ZN(
        n90867) );
  AOI22_X1 U76413 ( .A1(n90471), .A2(n107779), .B1(n90472), .B2(n70190), .ZN(
        n90866) );
  NAND2_X1 U76414 ( .A1(n90868), .A2(n90869), .ZN(n90864) );
  AOI22_X1 U76415 ( .A1(n90475), .A2(n70199), .B1(n90476), .B2(n107787), .ZN(
        n90869) );
  AOI22_X1 U76416 ( .A1(n90477), .A2(n107788), .B1(n90478), .B2(n107778), .ZN(
        n90868) );
  NAND2_X1 U76417 ( .A1(n90870), .A2(n90871), .ZN(n90863) );
  AOI22_X1 U76418 ( .A1(n90481), .A2(n107786), .B1(n90482), .B2(n107790), .ZN(
        n90871) );
  AOI22_X1 U76419 ( .A1(n90483), .A2(n107784), .B1(n90484), .B2(n107789), .ZN(
        n90870) );
  NAND2_X1 U76420 ( .A1(n90872), .A2(n90873), .ZN(n90862) );
  AOI22_X1 U76421 ( .A1(n90487), .A2(n70204), .B1(n90488), .B2(n107794), .ZN(
        n90873) );
  AOI22_X1 U76422 ( .A1(n90489), .A2(n70202), .B1(n90490), .B2(n107783), .ZN(
        n90872) );
  NAND2_X1 U76423 ( .A1(n90874), .A2(n90875), .ZN(n90792) );
  NOR4_X1 U76424 ( .A1(n90876), .A2(n90877), .A3(n90878), .A4(n90879), .ZN(
        n90875) );
  NAND2_X1 U76425 ( .A1(n90880), .A2(n90881), .ZN(n90879) );
  AOI22_X1 U76426 ( .A1(n90499), .A2(n107819), .B1(n90500), .B2(n107818), .ZN(
        n90881) );
  AOI22_X1 U76427 ( .A1(n90501), .A2(n70238), .B1(n90502), .B2(n107816), .ZN(
        n90880) );
  NAND2_X1 U76428 ( .A1(n90882), .A2(n90883), .ZN(n90878) );
  AOI22_X1 U76429 ( .A1(n90505), .A2(n107814), .B1(n90506), .B2(n107817), .ZN(
        n90883) );
  AOI22_X1 U76430 ( .A1(n90507), .A2(n70244), .B1(n90508), .B2(n107815), .ZN(
        n90882) );
  NAND2_X1 U76431 ( .A1(n90884), .A2(n90885), .ZN(n90877) );
  AOI22_X1 U76432 ( .A1(n105650), .A2(n107824), .B1(n90512), .B2(n70250), .ZN(
        n90885) );
  AOI22_X1 U76433 ( .A1(n90513), .A2(n107822), .B1(n90514), .B2(n107823), .ZN(
        n90884) );
  NAND2_X1 U76434 ( .A1(n90886), .A2(n90887), .ZN(n90876) );
  AOI22_X1 U76435 ( .A1(n90517), .A2(n70242), .B1(n90518), .B2(n107821), .ZN(
        n90887) );
  AOI22_X1 U76436 ( .A1(n90519), .A2(n70249), .B1(n105644), .B2(n107820), .ZN(
        n90886) );
  NOR4_X1 U76437 ( .A1(n90888), .A2(n90889), .A3(n90890), .A4(n90891), .ZN(
        n90874) );
  NAND2_X1 U76438 ( .A1(n90892), .A2(n90893), .ZN(n90891) );
  AOI22_X1 U76439 ( .A1(n90527), .A2(n107801), .B1(n90528), .B2(n107805), .ZN(
        n90893) );
  AOI22_X1 U76440 ( .A1(n90529), .A2(n107804), .B1(n90530), .B2(n70221), .ZN(
        n90892) );
  NAND2_X1 U76441 ( .A1(n90894), .A2(n90895), .ZN(n90890) );
  AOI22_X1 U76442 ( .A1(n90533), .A2(n107810), .B1(n90534), .B2(n107800), .ZN(
        n90895) );
  AOI22_X1 U76443 ( .A1(n90535), .A2(n107803), .B1(n90536), .B2(n107807), .ZN(
        n90894) );
  NAND2_X1 U76444 ( .A1(n90896), .A2(n90897), .ZN(n90889) );
  AOI22_X1 U76445 ( .A1(n90539), .A2(n107806), .B1(n90540), .B2(n107811), .ZN(
        n90897) );
  AOI22_X1 U76446 ( .A1(n90541), .A2(n107813), .B1(n90542), .B2(n107809), .ZN(
        n90896) );
  NAND2_X1 U76447 ( .A1(n90898), .A2(n90899), .ZN(n90888) );
  AOI22_X1 U76448 ( .A1(n90545), .A2(n70239), .B1(n90546), .B2(n70225), .ZN(
        n90899) );
  AOI22_X1 U76449 ( .A1(n90547), .A2(n70228), .B1(n90548), .B2(n107812), .ZN(
        n90898) );
  AOI21_X1 U76450 ( .B1(n90295), .B2(n86912), .A(n90901), .ZN(n90900) );
  OAI21_X1 U76451 ( .B1(n90902), .B2(n105659), .A(n90903), .ZN(n90901) );
  OAI21_X1 U76452 ( .B1(n90904), .B2(n90905), .A(n90302), .ZN(n90903) );
  OAI21_X1 U76453 ( .B1(n102120), .B2(n90303), .A(n90906), .ZN(n90905) );
  AOI22_X1 U76454 ( .A1(n90305), .A2(n110741), .B1(n90306), .B2(n74126), .ZN(
        n90906) );
  NAND2_X1 U76455 ( .A1(n90907), .A2(n90908), .ZN(n90904) );
  AOI22_X1 U76456 ( .A1(n90309), .A2(n110746), .B1(n105653), .B2(n110743), 
        .ZN(n90908) );
  AOI22_X1 U76457 ( .A1(n90311), .A2(n74124), .B1(n90312), .B2(n110742), .ZN(
        n90907) );
  NOR4_X1 U76458 ( .A1(n90909), .A2(n90910), .A3(n90911), .A4(n90912), .ZN(
        n90902) );
  NAND2_X1 U76459 ( .A1(n90913), .A2(n90914), .ZN(n90912) );
  NOR4_X1 U76460 ( .A1(n90915), .A2(n90916), .A3(n90917), .A4(n90918), .ZN(
        n90914) );
  NAND2_X1 U76461 ( .A1(n90919), .A2(n90920), .ZN(n90918) );
  AOI22_X1 U76462 ( .A1(n90325), .A2(n110722), .B1(n90326), .B2(n110723), .ZN(
        n90920) );
  AOI22_X1 U76463 ( .A1(n90327), .A2(n110731), .B1(n90328), .B2(n110729), .ZN(
        n90919) );
  NAND2_X1 U76464 ( .A1(n90921), .A2(n90922), .ZN(n90917) );
  AOI22_X1 U76465 ( .A1(n90331), .A2(n73993), .B1(n90332), .B2(n110726), .ZN(
        n90922) );
  AOI22_X1 U76466 ( .A1(n90333), .A2(n74097), .B1(n90334), .B2(n110655), .ZN(
        n90921) );
  NAND2_X1 U76467 ( .A1(n90923), .A2(n90924), .ZN(n90916) );
  AOI22_X1 U76468 ( .A1(n90337), .A2(n110659), .B1(n90338), .B2(n73997), .ZN(
        n90924) );
  AOI22_X1 U76469 ( .A1(n90339), .A2(n110727), .B1(n90340), .B2(n110724), .ZN(
        n90923) );
  NAND2_X1 U76470 ( .A1(n90925), .A2(n90926), .ZN(n90915) );
  AOI22_X1 U76471 ( .A1(n90343), .A2(n110657), .B1(n90344), .B2(n110661), .ZN(
        n90926) );
  AOI22_X1 U76472 ( .A1(n90345), .A2(n110660), .B1(n90346), .B2(n73999), .ZN(
        n90925) );
  NOR4_X1 U76473 ( .A1(n90927), .A2(n90928), .A3(n90929), .A4(n90930), .ZN(
        n90913) );
  NAND2_X1 U76474 ( .A1(n90931), .A2(n90932), .ZN(n90930) );
  AOI22_X1 U76475 ( .A1(n90353), .A2(n110732), .B1(n90354), .B2(n110735), .ZN(
        n90932) );
  AOI22_X1 U76476 ( .A1(n90355), .A2(n110736), .B1(n90356), .B2(n110738), .ZN(
        n90931) );
  NAND2_X1 U76477 ( .A1(n90933), .A2(n90934), .ZN(n90929) );
  AOI22_X1 U76478 ( .A1(n90359), .A2(n110737), .B1(n90360), .B2(n110733), .ZN(
        n90934) );
  AOI22_X1 U76479 ( .A1(n90361), .A2(n110739), .B1(n90362), .B2(n110734), .ZN(
        n90933) );
  NAND2_X1 U76480 ( .A1(n90935), .A2(n90936), .ZN(n90928) );
  AOI22_X1 U76481 ( .A1(n90365), .A2(n74107), .B1(n90366), .B2(n74106), .ZN(
        n90936) );
  AOI22_X1 U76482 ( .A1(n90367), .A2(n74109), .B1(n90368), .B2(n110740), .ZN(
        n90935) );
  NAND2_X1 U76483 ( .A1(n90937), .A2(n90938), .ZN(n90927) );
  AOI22_X1 U76484 ( .A1(n90371), .A2(n110725), .B1(n90372), .B2(n110730), .ZN(
        n90938) );
  AOI22_X1 U76485 ( .A1(n90373), .A2(n74104), .B1(n90374), .B2(n110728), .ZN(
        n90937) );
  NAND2_X1 U76486 ( .A1(n90939), .A2(n90940), .ZN(n90911) );
  NOR4_X1 U76487 ( .A1(n90941), .A2(n90942), .A3(n90943), .A4(n90944), .ZN(
        n90940) );
  NAND2_X1 U76488 ( .A1(n90945), .A2(n90946), .ZN(n90944) );
  AOI22_X1 U76489 ( .A1(n90383), .A2(n110670), .B1(n90384), .B2(n110672), .ZN(
        n90946) );
  AOI22_X1 U76490 ( .A1(n90385), .A2(n74022), .B1(n90386), .B2(n110671), .ZN(
        n90945) );
  NAND2_X1 U76491 ( .A1(n90947), .A2(n90948), .ZN(n90943) );
  AOI22_X1 U76492 ( .A1(n90389), .A2(n74026), .B1(n90390), .B2(n74028), .ZN(
        n90948) );
  AOI22_X1 U76493 ( .A1(n90391), .A2(n110677), .B1(n90392), .B2(n110678), .ZN(
        n90947) );
  NAND2_X1 U76494 ( .A1(n90949), .A2(n90950), .ZN(n90942) );
  AOI22_X1 U76495 ( .A1(n90395), .A2(n110675), .B1(n90396), .B2(n110676), .ZN(
        n90950) );
  AOI22_X1 U76496 ( .A1(n90397), .A2(n110679), .B1(n90398), .B2(n74021), .ZN(
        n90949) );
  NAND2_X1 U76497 ( .A1(n90951), .A2(n90952), .ZN(n90941) );
  AOI22_X1 U76498 ( .A1(n90401), .A2(n110683), .B1(n90402), .B2(n74033), .ZN(
        n90952) );
  AOI22_X1 U76499 ( .A1(n90403), .A2(n110682), .B1(n90404), .B2(n74031), .ZN(
        n90951) );
  NOR4_X1 U76500 ( .A1(n90953), .A2(n90954), .A3(n90955), .A4(n90956), .ZN(
        n90939) );
  NAND2_X1 U76501 ( .A1(n90957), .A2(n90958), .ZN(n90956) );
  AOI22_X1 U76502 ( .A1(n90411), .A2(n110665), .B1(n90412), .B2(n110656), .ZN(
        n90958) );
  AOI22_X1 U76503 ( .A1(n90413), .A2(n110658), .B1(n90414), .B2(n74005), .ZN(
        n90957) );
  NAND2_X1 U76504 ( .A1(n90959), .A2(n90960), .ZN(n90955) );
  AOI22_X1 U76505 ( .A1(n90417), .A2(n110663), .B1(n90418), .B2(n110667), .ZN(
        n90960) );
  AOI22_X1 U76506 ( .A1(n90419), .A2(n110669), .B1(n90420), .B2(n110666), .ZN(
        n90959) );
  NAND2_X1 U76507 ( .A1(n90961), .A2(n90962), .ZN(n90954) );
  AOI22_X1 U76508 ( .A1(n90423), .A2(n74014), .B1(n90424), .B2(n110662), .ZN(
        n90962) );
  AOI22_X1 U76509 ( .A1(n90425), .A2(n110664), .B1(n90426), .B2(n110668), .ZN(
        n90961) );
  NAND2_X1 U76510 ( .A1(n90963), .A2(n90964), .ZN(n90953) );
  AOI22_X1 U76511 ( .A1(n90429), .A2(n110674), .B1(n90430), .B2(n74018), .ZN(
        n90964) );
  AOI22_X1 U76512 ( .A1(n90431), .A2(n74016), .B1(n90432), .B2(n110673), .ZN(
        n90963) );
  NAND2_X1 U76513 ( .A1(n90965), .A2(n90966), .ZN(n90910) );
  NOR4_X1 U76514 ( .A1(n90967), .A2(n90968), .A3(n90969), .A4(n90970), .ZN(
        n90966) );
  NAND2_X1 U76515 ( .A1(n90971), .A2(n90972), .ZN(n90970) );
  AOI22_X1 U76516 ( .A1(n90441), .A2(n74056), .B1(n90442), .B2(n110692), .ZN(
        n90972) );
  AOI22_X1 U76517 ( .A1(n90443), .A2(n110695), .B1(n90444), .B2(n74052), .ZN(
        n90971) );
  NAND2_X1 U76518 ( .A1(n90973), .A2(n90974), .ZN(n90969) );
  AOI22_X1 U76519 ( .A1(n90447), .A2(n110698), .B1(n90448), .B2(n110697), .ZN(
        n90974) );
  AOI22_X1 U76520 ( .A1(n90449), .A2(n110691), .B1(n90450), .B2(n110693), .ZN(
        n90973) );
  NAND2_X1 U76521 ( .A1(n90975), .A2(n90976), .ZN(n90968) );
  AOI22_X1 U76522 ( .A1(n90453), .A2(n74061), .B1(n90454), .B2(n74055), .ZN(
        n90976) );
  AOI22_X1 U76523 ( .A1(n90455), .A2(n74060), .B1(n90456), .B2(n74062), .ZN(
        n90975) );
  NAND2_X1 U76524 ( .A1(n90977), .A2(n90978), .ZN(n90967) );
  AOI22_X1 U76525 ( .A1(n90459), .A2(n74065), .B1(n90460), .B2(n74068), .ZN(
        n90978) );
  AOI22_X1 U76526 ( .A1(n90461), .A2(n110696), .B1(n90462), .B2(n74057), .ZN(
        n90977) );
  NOR4_X1 U76527 ( .A1(n90979), .A2(n90980), .A3(n90981), .A4(n90982), .ZN(
        n90965) );
  NAND2_X1 U76528 ( .A1(n90983), .A2(n90984), .ZN(n90982) );
  AOI22_X1 U76529 ( .A1(n90469), .A2(n74032), .B1(n90470), .B2(n110686), .ZN(
        n90984) );
  AOI22_X1 U76530 ( .A1(n90471), .A2(n110681), .B1(n90472), .B2(n74036), .ZN(
        n90983) );
  NAND2_X1 U76531 ( .A1(n90985), .A2(n90986), .ZN(n90981) );
  AOI22_X1 U76532 ( .A1(n90475), .A2(n74045), .B1(n90476), .B2(n110688), .ZN(
        n90986) );
  AOI22_X1 U76533 ( .A1(n90477), .A2(n110689), .B1(n90478), .B2(n110680), .ZN(
        n90985) );
  NAND2_X1 U76534 ( .A1(n90987), .A2(n90988), .ZN(n90980) );
  AOI22_X1 U76535 ( .A1(n90481), .A2(n110687), .B1(n90482), .B2(n74044), .ZN(
        n90988) );
  AOI22_X1 U76536 ( .A1(n90483), .A2(n110685), .B1(n90484), .B2(n110690), .ZN(
        n90987) );
  NAND2_X1 U76537 ( .A1(n90989), .A2(n90990), .ZN(n90979) );
  AOI22_X1 U76538 ( .A1(n90487), .A2(n74050), .B1(n90488), .B2(n110694), .ZN(
        n90990) );
  AOI22_X1 U76539 ( .A1(n90489), .A2(n74048), .B1(n90490), .B2(n110684), .ZN(
        n90989) );
  NAND2_X1 U76540 ( .A1(n90991), .A2(n90992), .ZN(n90909) );
  NOR4_X1 U76541 ( .A1(n90993), .A2(n90994), .A3(n90995), .A4(n90996), .ZN(
        n90992) );
  NAND2_X1 U76542 ( .A1(n90997), .A2(n90998), .ZN(n90996) );
  AOI22_X1 U76543 ( .A1(n90499), .A2(n110715), .B1(n90500), .B2(n110714), .ZN(
        n90998) );
  AOI22_X1 U76544 ( .A1(n90501), .A2(n74084), .B1(n90502), .B2(n110712), .ZN(
        n90997) );
  NAND2_X1 U76545 ( .A1(n90999), .A2(n91000), .ZN(n90995) );
  AOI22_X1 U76546 ( .A1(n90505), .A2(n110710), .B1(n90506), .B2(n110713), .ZN(
        n91000) );
  AOI22_X1 U76547 ( .A1(n90507), .A2(n74090), .B1(n90508), .B2(n110711), .ZN(
        n90999) );
  NAND2_X1 U76548 ( .A1(n91001), .A2(n91002), .ZN(n90994) );
  AOI22_X1 U76549 ( .A1(n105650), .A2(n110720), .B1(n90512), .B2(n74096), .ZN(
        n91002) );
  AOI22_X1 U76550 ( .A1(n90513), .A2(n110718), .B1(n90514), .B2(n110719), .ZN(
        n91001) );
  NAND2_X1 U76551 ( .A1(n91003), .A2(n91004), .ZN(n90993) );
  AOI22_X1 U76552 ( .A1(n90517), .A2(n74088), .B1(n90518), .B2(n110717), .ZN(
        n91004) );
  AOI22_X1 U76553 ( .A1(n90519), .A2(n74095), .B1(n105644), .B2(n110716), .ZN(
        n91003) );
  NOR4_X1 U76554 ( .A1(n91005), .A2(n91006), .A3(n91007), .A4(n91008), .ZN(
        n90991) );
  NAND2_X1 U76555 ( .A1(n91009), .A2(n91010), .ZN(n91008) );
  AOI22_X1 U76556 ( .A1(n90527), .A2(n110700), .B1(n90528), .B2(n110702), .ZN(
        n91010) );
  AOI22_X1 U76557 ( .A1(n90529), .A2(n74069), .B1(n90530), .B2(n74067), .ZN(
        n91009) );
  NAND2_X1 U76558 ( .A1(n91011), .A2(n91012), .ZN(n91007) );
  AOI22_X1 U76559 ( .A1(n90533), .A2(n110707), .B1(n90534), .B2(n110699), .ZN(
        n91012) );
  AOI22_X1 U76560 ( .A1(n90535), .A2(n110701), .B1(n90536), .B2(n110704), .ZN(
        n91011) );
  NAND2_X1 U76561 ( .A1(n91013), .A2(n91014), .ZN(n91006) );
  AOI22_X1 U76562 ( .A1(n90539), .A2(n110703), .B1(n90540), .B2(n74077), .ZN(
        n91014) );
  AOI22_X1 U76563 ( .A1(n90541), .A2(n110709), .B1(n90542), .B2(n110706), .ZN(
        n91013) );
  NAND2_X1 U76564 ( .A1(n91015), .A2(n91016), .ZN(n91005) );
  AOI22_X1 U76565 ( .A1(n90545), .A2(n74085), .B1(n90546), .B2(n74071), .ZN(
        n91016) );
  AOI22_X1 U76566 ( .A1(n90547), .A2(n110705), .B1(n90548), .B2(n110708), .ZN(
        n91015) );
  AOI21_X1 U76567 ( .B1(n90295), .B2(n87030), .A(n91018), .ZN(n91017) );
  OAI21_X1 U76568 ( .B1(n91019), .B2(n105659), .A(n91020), .ZN(n91018) );
  OAI21_X1 U76569 ( .B1(n91021), .B2(n91022), .A(n90302), .ZN(n91020) );
  OAI21_X1 U76570 ( .B1(n102106), .B2(n90303), .A(n91023), .ZN(n91022) );
  AOI22_X1 U76571 ( .A1(n90305), .A2(n108146), .B1(n90306), .B2(n70713), .ZN(
        n91023) );
  NAND2_X1 U76572 ( .A1(n91024), .A2(n91025), .ZN(n91021) );
  AOI22_X1 U76573 ( .A1(n90309), .A2(n108151), .B1(n105653), .B2(n108148), 
        .ZN(n91025) );
  AOI22_X1 U76574 ( .A1(n90311), .A2(n70711), .B1(n90312), .B2(n108147), .ZN(
        n91024) );
  NOR4_X1 U76575 ( .A1(n91026), .A2(n91027), .A3(n91028), .A4(n91029), .ZN(
        n91019) );
  NAND2_X1 U76576 ( .A1(n91030), .A2(n91031), .ZN(n91029) );
  NOR4_X1 U76577 ( .A1(n91032), .A2(n91033), .A3(n91034), .A4(n91035), .ZN(
        n91031) );
  NAND2_X1 U76578 ( .A1(n91036), .A2(n91037), .ZN(n91035) );
  AOI22_X1 U76579 ( .A1(n90325), .A2(n108126), .B1(n90326), .B2(n108127), .ZN(
        n91037) );
  AOI22_X1 U76580 ( .A1(n90327), .A2(n108136), .B1(n90328), .B2(n108134), .ZN(
        n91036) );
  NAND2_X1 U76581 ( .A1(n91038), .A2(n91039), .ZN(n91034) );
  AOI22_X1 U76582 ( .A1(n90331), .A2(n70580), .B1(n90332), .B2(n108130), .ZN(
        n91039) );
  AOI22_X1 U76583 ( .A1(n90333), .A2(n70684), .B1(n90334), .B2(n108054), .ZN(
        n91038) );
  NAND2_X1 U76584 ( .A1(n91040), .A2(n91041), .ZN(n91033) );
  AOI22_X1 U76585 ( .A1(n90337), .A2(n108058), .B1(n90338), .B2(n70584), .ZN(
        n91041) );
  AOI22_X1 U76586 ( .A1(n90339), .A2(n108131), .B1(n90340), .B2(n108128), .ZN(
        n91040) );
  NAND2_X1 U76587 ( .A1(n91042), .A2(n91043), .ZN(n91032) );
  AOI22_X1 U76588 ( .A1(n90343), .A2(n108056), .B1(n90344), .B2(n108060), .ZN(
        n91043) );
  AOI22_X1 U76589 ( .A1(n90345), .A2(n108059), .B1(n90346), .B2(n70586), .ZN(
        n91042) );
  NOR4_X1 U76590 ( .A1(n91044), .A2(n91045), .A3(n91046), .A4(n91047), .ZN(
        n91030) );
  NAND2_X1 U76591 ( .A1(n91048), .A2(n91049), .ZN(n91047) );
  AOI22_X1 U76592 ( .A1(n90353), .A2(n108137), .B1(n90354), .B2(n108140), .ZN(
        n91049) );
  AOI22_X1 U76593 ( .A1(n90355), .A2(n108141), .B1(n90356), .B2(n108143), .ZN(
        n91048) );
  NAND2_X1 U76594 ( .A1(n91050), .A2(n91051), .ZN(n91046) );
  AOI22_X1 U76595 ( .A1(n90359), .A2(n108142), .B1(n90360), .B2(n108138), .ZN(
        n91051) );
  AOI22_X1 U76596 ( .A1(n90361), .A2(n108144), .B1(n90362), .B2(n108139), .ZN(
        n91050) );
  NAND2_X1 U76597 ( .A1(n91052), .A2(n91053), .ZN(n91045) );
  AOI22_X1 U76598 ( .A1(n90365), .A2(n70694), .B1(n90366), .B2(n70693), .ZN(
        n91053) );
  AOI22_X1 U76599 ( .A1(n90367), .A2(n70696), .B1(n90368), .B2(n108145), .ZN(
        n91052) );
  NAND2_X1 U76600 ( .A1(n91054), .A2(n91055), .ZN(n91044) );
  AOI22_X1 U76601 ( .A1(n90371), .A2(n108129), .B1(n90372), .B2(n108135), .ZN(
        n91055) );
  AOI22_X1 U76602 ( .A1(n90373), .A2(n70691), .B1(n90374), .B2(n108133), .ZN(
        n91054) );
  NAND2_X1 U76603 ( .A1(n91056), .A2(n91057), .ZN(n91028) );
  NOR4_X1 U76604 ( .A1(n91058), .A2(n91059), .A3(n91060), .A4(n91061), .ZN(
        n91057) );
  NAND2_X1 U76605 ( .A1(n91062), .A2(n91063), .ZN(n91061) );
  AOI22_X1 U76606 ( .A1(n90383), .A2(n108069), .B1(n90384), .B2(n108071), .ZN(
        n91063) );
  AOI22_X1 U76607 ( .A1(n90385), .A2(n70609), .B1(n90386), .B2(n108070), .ZN(
        n91062) );
  NAND2_X1 U76608 ( .A1(n91064), .A2(n91065), .ZN(n91060) );
  AOI22_X1 U76609 ( .A1(n90389), .A2(n70613), .B1(n90390), .B2(n70615), .ZN(
        n91065) );
  AOI22_X1 U76610 ( .A1(n90391), .A2(n108077), .B1(n90392), .B2(n108078), .ZN(
        n91064) );
  NAND2_X1 U76611 ( .A1(n91066), .A2(n91067), .ZN(n91059) );
  AOI22_X1 U76612 ( .A1(n90395), .A2(n108074), .B1(n90396), .B2(n108076), .ZN(
        n91067) );
  AOI22_X1 U76613 ( .A1(n90397), .A2(n108079), .B1(n90398), .B2(n108075), .ZN(
        n91066) );
  NAND2_X1 U76614 ( .A1(n91068), .A2(n91069), .ZN(n91058) );
  AOI22_X1 U76615 ( .A1(n90401), .A2(n108083), .B1(n90402), .B2(n70620), .ZN(
        n91069) );
  AOI22_X1 U76616 ( .A1(n90403), .A2(n108082), .B1(n90404), .B2(n70618), .ZN(
        n91068) );
  NOR4_X1 U76617 ( .A1(n91070), .A2(n91071), .A3(n91072), .A4(n91073), .ZN(
        n91056) );
  NAND2_X1 U76618 ( .A1(n91074), .A2(n91075), .ZN(n91073) );
  AOI22_X1 U76619 ( .A1(n90411), .A2(n108064), .B1(n90412), .B2(n108055), .ZN(
        n91075) );
  AOI22_X1 U76620 ( .A1(n90413), .A2(n108057), .B1(n90414), .B2(n70592), .ZN(
        n91074) );
  NAND2_X1 U76621 ( .A1(n91076), .A2(n91077), .ZN(n91072) );
  AOI22_X1 U76622 ( .A1(n90417), .A2(n108062), .B1(n90418), .B2(n108066), .ZN(
        n91077) );
  AOI22_X1 U76623 ( .A1(n90419), .A2(n108068), .B1(n90420), .B2(n108065), .ZN(
        n91076) );
  NAND2_X1 U76624 ( .A1(n91078), .A2(n91079), .ZN(n91071) );
  AOI22_X1 U76625 ( .A1(n90423), .A2(n70601), .B1(n90424), .B2(n108061), .ZN(
        n91079) );
  AOI22_X1 U76626 ( .A1(n90425), .A2(n108063), .B1(n90426), .B2(n108067), .ZN(
        n91078) );
  NAND2_X1 U76627 ( .A1(n91080), .A2(n91081), .ZN(n91070) );
  AOI22_X1 U76628 ( .A1(n90429), .A2(n108073), .B1(n90430), .B2(n70605), .ZN(
        n91081) );
  AOI22_X1 U76629 ( .A1(n90431), .A2(n70603), .B1(n90432), .B2(n108072), .ZN(
        n91080) );
  NAND2_X1 U76630 ( .A1(n91082), .A2(n91083), .ZN(n91027) );
  NOR4_X1 U76631 ( .A1(n91084), .A2(n91085), .A3(n91086), .A4(n91087), .ZN(
        n91083) );
  NAND2_X1 U76632 ( .A1(n91088), .A2(n91089), .ZN(n91087) );
  AOI22_X1 U76633 ( .A1(n90441), .A2(n70643), .B1(n90442), .B2(n108092), .ZN(
        n91089) );
  AOI22_X1 U76634 ( .A1(n90443), .A2(n108095), .B1(n90444), .B2(n70639), .ZN(
        n91088) );
  NAND2_X1 U76635 ( .A1(n91090), .A2(n91091), .ZN(n91086) );
  AOI22_X1 U76636 ( .A1(n90447), .A2(n108100), .B1(n90448), .B2(n108099), .ZN(
        n91091) );
  AOI22_X1 U76637 ( .A1(n90449), .A2(n108091), .B1(n90450), .B2(n108093), .ZN(
        n91090) );
  NAND2_X1 U76638 ( .A1(n91092), .A2(n91093), .ZN(n91085) );
  AOI22_X1 U76639 ( .A1(n90453), .A2(n108101), .B1(n90454), .B2(n108097), .ZN(
        n91093) );
  AOI22_X1 U76640 ( .A1(n90455), .A2(n70647), .B1(n90456), .B2(n70649), .ZN(
        n91092) );
  NAND2_X1 U76641 ( .A1(n91094), .A2(n91095), .ZN(n91084) );
  AOI22_X1 U76642 ( .A1(n90459), .A2(n70652), .B1(n90460), .B2(n70655), .ZN(
        n91095) );
  AOI22_X1 U76643 ( .A1(n90461), .A2(n108096), .B1(n90462), .B2(n108098), .ZN(
        n91094) );
  NOR4_X1 U76644 ( .A1(n91096), .A2(n91097), .A3(n91098), .A4(n91099), .ZN(
        n91082) );
  NAND2_X1 U76645 ( .A1(n91100), .A2(n91101), .ZN(n91099) );
  AOI22_X1 U76646 ( .A1(n90469), .A2(n70619), .B1(n90470), .B2(n108086), .ZN(
        n91101) );
  AOI22_X1 U76647 ( .A1(n90471), .A2(n108081), .B1(n90472), .B2(n70623), .ZN(
        n91100) );
  NAND2_X1 U76648 ( .A1(n91102), .A2(n91103), .ZN(n91098) );
  AOI22_X1 U76649 ( .A1(n90475), .A2(n70632), .B1(n90476), .B2(n108088), .ZN(
        n91103) );
  AOI22_X1 U76650 ( .A1(n90477), .A2(n108089), .B1(n90478), .B2(n108080), .ZN(
        n91102) );
  NAND2_X1 U76651 ( .A1(n91104), .A2(n91105), .ZN(n91097) );
  AOI22_X1 U76652 ( .A1(n90481), .A2(n108087), .B1(n90482), .B2(n70631), .ZN(
        n91105) );
  AOI22_X1 U76653 ( .A1(n90483), .A2(n108085), .B1(n90484), .B2(n108090), .ZN(
        n91104) );
  NAND2_X1 U76654 ( .A1(n91106), .A2(n91107), .ZN(n91096) );
  AOI22_X1 U76655 ( .A1(n90487), .A2(n70637), .B1(n90488), .B2(n108094), .ZN(
        n91107) );
  AOI22_X1 U76656 ( .A1(n90489), .A2(n70635), .B1(n90490), .B2(n108084), .ZN(
        n91106) );
  NAND2_X1 U76657 ( .A1(n91108), .A2(n91109), .ZN(n91026) );
  NOR4_X1 U76658 ( .A1(n91110), .A2(n91111), .A3(n91112), .A4(n91113), .ZN(
        n91109) );
  NAND2_X1 U76659 ( .A1(n91114), .A2(n91115), .ZN(n91113) );
  AOI22_X1 U76660 ( .A1(n90499), .A2(n108118), .B1(n90500), .B2(n108117), .ZN(
        n91115) );
  AOI22_X1 U76661 ( .A1(n90501), .A2(n70671), .B1(n90502), .B2(n108115), .ZN(
        n91114) );
  NAND2_X1 U76662 ( .A1(n91116), .A2(n91117), .ZN(n91112) );
  AOI22_X1 U76663 ( .A1(n90505), .A2(n108113), .B1(n90506), .B2(n108116), .ZN(
        n91117) );
  AOI22_X1 U76664 ( .A1(n90507), .A2(n70677), .B1(n90508), .B2(n108114), .ZN(
        n91116) );
  NAND2_X1 U76665 ( .A1(n91118), .A2(n91119), .ZN(n91111) );
  AOI22_X1 U76666 ( .A1(n105650), .A2(n108123), .B1(n90512), .B2(n70683), .ZN(
        n91119) );
  AOI22_X1 U76667 ( .A1(n90513), .A2(n108121), .B1(n90514), .B2(n108122), .ZN(
        n91118) );
  NAND2_X1 U76668 ( .A1(n91120), .A2(n91121), .ZN(n91110) );
  AOI22_X1 U76669 ( .A1(n90517), .A2(n70675), .B1(n90518), .B2(n108120), .ZN(
        n91121) );
  AOI22_X1 U76670 ( .A1(n90519), .A2(n108124), .B1(n105644), .B2(n108119), 
        .ZN(n91120) );
  NOR4_X1 U76671 ( .A1(n91122), .A2(n91123), .A3(n91124), .A4(n91125), .ZN(
        n91108) );
  NAND2_X1 U76672 ( .A1(n91126), .A2(n91127), .ZN(n91125) );
  AOI22_X1 U76673 ( .A1(n90527), .A2(n108103), .B1(n90528), .B2(n108105), .ZN(
        n91127) );
  AOI22_X1 U76674 ( .A1(n90529), .A2(n70656), .B1(n90530), .B2(n70654), .ZN(
        n91126) );
  NAND2_X1 U76675 ( .A1(n91128), .A2(n91129), .ZN(n91124) );
  AOI22_X1 U76676 ( .A1(n90533), .A2(n108110), .B1(n90534), .B2(n108102), .ZN(
        n91129) );
  AOI22_X1 U76677 ( .A1(n90535), .A2(n108104), .B1(n90536), .B2(n108107), .ZN(
        n91128) );
  NAND2_X1 U76678 ( .A1(n91130), .A2(n91131), .ZN(n91123) );
  AOI22_X1 U76679 ( .A1(n90539), .A2(n108106), .B1(n90540), .B2(n70664), .ZN(
        n91131) );
  AOI22_X1 U76680 ( .A1(n90541), .A2(n108112), .B1(n90542), .B2(n108109), .ZN(
        n91130) );
  NAND2_X1 U76681 ( .A1(n91132), .A2(n91133), .ZN(n91122) );
  AOI22_X1 U76682 ( .A1(n90545), .A2(n70672), .B1(n90546), .B2(n70658), .ZN(
        n91133) );
  AOI22_X1 U76683 ( .A1(n90547), .A2(n108108), .B1(n90548), .B2(n108111), .ZN(
        n91132) );
  AOI21_X1 U76684 ( .B1(n90295), .B2(n87148), .A(n91135), .ZN(n91134) );
  OAI21_X1 U76685 ( .B1(n91136), .B2(n105659), .A(n91137), .ZN(n91135) );
  OAI21_X1 U76686 ( .B1(n91138), .B2(n91139), .A(n90302), .ZN(n91137) );
  OAI21_X1 U76687 ( .B1(n102092), .B2(n90303), .A(n91140), .ZN(n91139) );
  AOI22_X1 U76688 ( .A1(n90305), .A2(n110844), .B1(n90306), .B2(n74267), .ZN(
        n91140) );
  NAND2_X1 U76689 ( .A1(n91141), .A2(n91142), .ZN(n91138) );
  AOI22_X1 U76690 ( .A1(n90309), .A2(n110849), .B1(n105653), .B2(n110846), 
        .ZN(n91142) );
  AOI22_X1 U76691 ( .A1(n90311), .A2(n74265), .B1(n90312), .B2(n110845), .ZN(
        n91141) );
  NOR4_X1 U76692 ( .A1(n91143), .A2(n91144), .A3(n91145), .A4(n91146), .ZN(
        n91136) );
  NAND2_X1 U76693 ( .A1(n91147), .A2(n91148), .ZN(n91146) );
  NOR4_X1 U76694 ( .A1(n91149), .A2(n91150), .A3(n91151), .A4(n91152), .ZN(
        n91148) );
  NAND2_X1 U76695 ( .A1(n91153), .A2(n91154), .ZN(n91152) );
  AOI22_X1 U76696 ( .A1(n90325), .A2(n110825), .B1(n90326), .B2(n110826), .ZN(
        n91154) );
  AOI22_X1 U76697 ( .A1(n90327), .A2(n110834), .B1(n90328), .B2(n110832), .ZN(
        n91153) );
  NAND2_X1 U76698 ( .A1(n91155), .A2(n91156), .ZN(n91151) );
  AOI22_X1 U76699 ( .A1(n90331), .A2(n74134), .B1(n90332), .B2(n110829), .ZN(
        n91156) );
  AOI22_X1 U76700 ( .A1(n90333), .A2(n74238), .B1(n90334), .B2(n110752), .ZN(
        n91155) );
  NAND2_X1 U76701 ( .A1(n91157), .A2(n91158), .ZN(n91150) );
  AOI22_X1 U76702 ( .A1(n90337), .A2(n110756), .B1(n90338), .B2(n74138), .ZN(
        n91158) );
  AOI22_X1 U76703 ( .A1(n90339), .A2(n110830), .B1(n90340), .B2(n110827), .ZN(
        n91157) );
  NAND2_X1 U76704 ( .A1(n91159), .A2(n91160), .ZN(n91149) );
  AOI22_X1 U76705 ( .A1(n90343), .A2(n110754), .B1(n90344), .B2(n110758), .ZN(
        n91160) );
  AOI22_X1 U76706 ( .A1(n90345), .A2(n110757), .B1(n90346), .B2(n74140), .ZN(
        n91159) );
  NOR4_X1 U76707 ( .A1(n91161), .A2(n91162), .A3(n91163), .A4(n91164), .ZN(
        n91147) );
  NAND2_X1 U76708 ( .A1(n91165), .A2(n91166), .ZN(n91164) );
  AOI22_X1 U76709 ( .A1(n90353), .A2(n110835), .B1(n90354), .B2(n110838), .ZN(
        n91166) );
  AOI22_X1 U76710 ( .A1(n90355), .A2(n110839), .B1(n90356), .B2(n110841), .ZN(
        n91165) );
  NAND2_X1 U76711 ( .A1(n91167), .A2(n91168), .ZN(n91163) );
  AOI22_X1 U76712 ( .A1(n90359), .A2(n110840), .B1(n90360), .B2(n110836), .ZN(
        n91168) );
  AOI22_X1 U76713 ( .A1(n90361), .A2(n110842), .B1(n90362), .B2(n110837), .ZN(
        n91167) );
  NAND2_X1 U76714 ( .A1(n91169), .A2(n91170), .ZN(n91162) );
  AOI22_X1 U76715 ( .A1(n90365), .A2(n74248), .B1(n90366), .B2(n74247), .ZN(
        n91170) );
  AOI22_X1 U76716 ( .A1(n90367), .A2(n74250), .B1(n90368), .B2(n110843), .ZN(
        n91169) );
  NAND2_X1 U76717 ( .A1(n91171), .A2(n91172), .ZN(n91161) );
  AOI22_X1 U76718 ( .A1(n90371), .A2(n110828), .B1(n90372), .B2(n110833), .ZN(
        n91172) );
  AOI22_X1 U76719 ( .A1(n90373), .A2(n74245), .B1(n90374), .B2(n110831), .ZN(
        n91171) );
  NAND2_X1 U76720 ( .A1(n91173), .A2(n91174), .ZN(n91145) );
  NOR4_X1 U76721 ( .A1(n91175), .A2(n91176), .A3(n91177), .A4(n91178), .ZN(
        n91174) );
  NAND2_X1 U76722 ( .A1(n91179), .A2(n91180), .ZN(n91178) );
  AOI22_X1 U76723 ( .A1(n90383), .A2(n110767), .B1(n90384), .B2(n110769), .ZN(
        n91180) );
  AOI22_X1 U76724 ( .A1(n90385), .A2(n74163), .B1(n90386), .B2(n110768), .ZN(
        n91179) );
  NAND2_X1 U76725 ( .A1(n91181), .A2(n91182), .ZN(n91177) );
  AOI22_X1 U76726 ( .A1(n90389), .A2(n74167), .B1(n90390), .B2(n74169), .ZN(
        n91182) );
  AOI22_X1 U76727 ( .A1(n90391), .A2(n110774), .B1(n90392), .B2(n110775), .ZN(
        n91181) );
  NAND2_X1 U76728 ( .A1(n91183), .A2(n91184), .ZN(n91176) );
  AOI22_X1 U76729 ( .A1(n90395), .A2(n110772), .B1(n90396), .B2(n110773), .ZN(
        n91184) );
  AOI22_X1 U76730 ( .A1(n90397), .A2(n110776), .B1(n90398), .B2(n74162), .ZN(
        n91183) );
  NAND2_X1 U76731 ( .A1(n91185), .A2(n91186), .ZN(n91175) );
  AOI22_X1 U76732 ( .A1(n90401), .A2(n110781), .B1(n90402), .B2(n74174), .ZN(
        n91186) );
  AOI22_X1 U76733 ( .A1(n90403), .A2(n110780), .B1(n90404), .B2(n74172), .ZN(
        n91185) );
  NOR4_X1 U76734 ( .A1(n91187), .A2(n91188), .A3(n91189), .A4(n91190), .ZN(
        n91173) );
  NAND2_X1 U76735 ( .A1(n91191), .A2(n91192), .ZN(n91190) );
  AOI22_X1 U76736 ( .A1(n90411), .A2(n110762), .B1(n90412), .B2(n110753), .ZN(
        n91192) );
  AOI22_X1 U76737 ( .A1(n90413), .A2(n110755), .B1(n90414), .B2(n74146), .ZN(
        n91191) );
  NAND2_X1 U76738 ( .A1(n91193), .A2(n91194), .ZN(n91189) );
  AOI22_X1 U76739 ( .A1(n90417), .A2(n110760), .B1(n90418), .B2(n110764), .ZN(
        n91194) );
  AOI22_X1 U76740 ( .A1(n90419), .A2(n110766), .B1(n90420), .B2(n110763), .ZN(
        n91193) );
  NAND2_X1 U76741 ( .A1(n91195), .A2(n91196), .ZN(n91188) );
  AOI22_X1 U76742 ( .A1(n90423), .A2(n74155), .B1(n90424), .B2(n110759), .ZN(
        n91196) );
  AOI22_X1 U76743 ( .A1(n90425), .A2(n110761), .B1(n90426), .B2(n110765), .ZN(
        n91195) );
  NAND2_X1 U76744 ( .A1(n91197), .A2(n91198), .ZN(n91187) );
  AOI22_X1 U76745 ( .A1(n90429), .A2(n110771), .B1(n90430), .B2(n74159), .ZN(
        n91198) );
  AOI22_X1 U76746 ( .A1(n90431), .A2(n74157), .B1(n90432), .B2(n110770), .ZN(
        n91197) );
  NAND2_X1 U76747 ( .A1(n91199), .A2(n91200), .ZN(n91144) );
  NOR4_X1 U76748 ( .A1(n91201), .A2(n91202), .A3(n91203), .A4(n91204), .ZN(
        n91200) );
  NAND2_X1 U76749 ( .A1(n91205), .A2(n91206), .ZN(n91204) );
  AOI22_X1 U76750 ( .A1(n90441), .A2(n74197), .B1(n90442), .B2(n110791), .ZN(
        n91206) );
  AOI22_X1 U76751 ( .A1(n90443), .A2(n110795), .B1(n90444), .B2(n110794), .ZN(
        n91205) );
  NAND2_X1 U76752 ( .A1(n91207), .A2(n91208), .ZN(n91203) );
  AOI22_X1 U76753 ( .A1(n90447), .A2(n110799), .B1(n90448), .B2(n110798), .ZN(
        n91208) );
  AOI22_X1 U76754 ( .A1(n90449), .A2(n110790), .B1(n90450), .B2(n110792), .ZN(
        n91207) );
  NAND2_X1 U76755 ( .A1(n91209), .A2(n91210), .ZN(n91202) );
  AOI22_X1 U76756 ( .A1(n90453), .A2(n110800), .B1(n90454), .B2(n74196), .ZN(
        n91210) );
  AOI22_X1 U76757 ( .A1(n90455), .A2(n74201), .B1(n90456), .B2(n74203), .ZN(
        n91209) );
  NAND2_X1 U76758 ( .A1(n91211), .A2(n91212), .ZN(n91201) );
  AOI22_X1 U76759 ( .A1(n90459), .A2(n74206), .B1(n90460), .B2(n74209), .ZN(
        n91212) );
  AOI22_X1 U76760 ( .A1(n90461), .A2(n110796), .B1(n90462), .B2(n110797), .ZN(
        n91211) );
  NOR4_X1 U76761 ( .A1(n91213), .A2(n91214), .A3(n91215), .A4(n91216), .ZN(
        n91199) );
  NAND2_X1 U76762 ( .A1(n91217), .A2(n91218), .ZN(n91216) );
  AOI22_X1 U76763 ( .A1(n90469), .A2(n110779), .B1(n90470), .B2(n110784), .ZN(
        n91218) );
  AOI22_X1 U76764 ( .A1(n90471), .A2(n110778), .B1(n90472), .B2(n74177), .ZN(
        n91217) );
  NAND2_X1 U76765 ( .A1(n91219), .A2(n91220), .ZN(n91215) );
  AOI22_X1 U76766 ( .A1(n90475), .A2(n74186), .B1(n90476), .B2(n110786), .ZN(
        n91220) );
  AOI22_X1 U76767 ( .A1(n90477), .A2(n110787), .B1(n90478), .B2(n110777), .ZN(
        n91219) );
  NAND2_X1 U76768 ( .A1(n91221), .A2(n91222), .ZN(n91214) );
  AOI22_X1 U76769 ( .A1(n90481), .A2(n110785), .B1(n90482), .B2(n110789), .ZN(
        n91222) );
  AOI22_X1 U76770 ( .A1(n90483), .A2(n110783), .B1(n90484), .B2(n110788), .ZN(
        n91221) );
  NAND2_X1 U76771 ( .A1(n91223), .A2(n91224), .ZN(n91213) );
  AOI22_X1 U76772 ( .A1(n90487), .A2(n74191), .B1(n90488), .B2(n110793), .ZN(
        n91224) );
  AOI22_X1 U76773 ( .A1(n90489), .A2(n74189), .B1(n90490), .B2(n110782), .ZN(
        n91223) );
  NAND2_X1 U76774 ( .A1(n91225), .A2(n91226), .ZN(n91143) );
  NOR4_X1 U76775 ( .A1(n91227), .A2(n91228), .A3(n91229), .A4(n91230), .ZN(
        n91226) );
  NAND2_X1 U76776 ( .A1(n91231), .A2(n91232), .ZN(n91230) );
  AOI22_X1 U76777 ( .A1(n90499), .A2(n110817), .B1(n90500), .B2(n110816), .ZN(
        n91232) );
  AOI22_X1 U76778 ( .A1(n90501), .A2(n74225), .B1(n90502), .B2(n110814), .ZN(
        n91231) );
  NAND2_X1 U76779 ( .A1(n91233), .A2(n91234), .ZN(n91229) );
  AOI22_X1 U76780 ( .A1(n90505), .A2(n110812), .B1(n90506), .B2(n110815), .ZN(
        n91234) );
  AOI22_X1 U76781 ( .A1(n90507), .A2(n74231), .B1(n90508), .B2(n110813), .ZN(
        n91233) );
  NAND2_X1 U76782 ( .A1(n91235), .A2(n91236), .ZN(n91228) );
  AOI22_X1 U76783 ( .A1(n105650), .A2(n110822), .B1(n90512), .B2(n74237), .ZN(
        n91236) );
  AOI22_X1 U76784 ( .A1(n90513), .A2(n110820), .B1(n90514), .B2(n110821), .ZN(
        n91235) );
  NAND2_X1 U76785 ( .A1(n91237), .A2(n91238), .ZN(n91227) );
  AOI22_X1 U76786 ( .A1(n90517), .A2(n74229), .B1(n90518), .B2(n110819), .ZN(
        n91238) );
  AOI22_X1 U76787 ( .A1(n90519), .A2(n110823), .B1(n105644), .B2(n110818), 
        .ZN(n91237) );
  NOR4_X1 U76788 ( .A1(n91239), .A2(n91240), .A3(n91241), .A4(n91242), .ZN(
        n91225) );
  NAND2_X1 U76789 ( .A1(n91243), .A2(n91244), .ZN(n91242) );
  AOI22_X1 U76790 ( .A1(n90527), .A2(n110802), .B1(n90528), .B2(n110804), .ZN(
        n91244) );
  AOI22_X1 U76791 ( .A1(n90529), .A2(n74210), .B1(n90530), .B2(n74208), .ZN(
        n91243) );
  NAND2_X1 U76792 ( .A1(n91245), .A2(n91246), .ZN(n91241) );
  AOI22_X1 U76793 ( .A1(n90533), .A2(n110809), .B1(n90534), .B2(n110801), .ZN(
        n91246) );
  AOI22_X1 U76794 ( .A1(n90535), .A2(n110803), .B1(n90536), .B2(n110806), .ZN(
        n91245) );
  NAND2_X1 U76795 ( .A1(n91247), .A2(n91248), .ZN(n91240) );
  AOI22_X1 U76796 ( .A1(n90539), .A2(n110805), .B1(n90540), .B2(n74218), .ZN(
        n91248) );
  AOI22_X1 U76797 ( .A1(n90541), .A2(n110811), .B1(n90542), .B2(n110808), .ZN(
        n91247) );
  NAND2_X1 U76798 ( .A1(n91249), .A2(n91250), .ZN(n91239) );
  AOI22_X1 U76799 ( .A1(n90545), .A2(n74226), .B1(n90546), .B2(n74212), .ZN(
        n91250) );
  AOI22_X1 U76800 ( .A1(n90547), .A2(n110807), .B1(n90548), .B2(n110810), .ZN(
        n91249) );
  AOI21_X1 U76801 ( .B1(n90295), .B2(n87266), .A(n91252), .ZN(n91251) );
  OAI21_X1 U76802 ( .B1(n91253), .B2(n105659), .A(n91254), .ZN(n91252) );
  OAI21_X1 U76803 ( .B1(n91255), .B2(n91256), .A(n90302), .ZN(n91254) );
  OAI21_X1 U76804 ( .B1(n102075), .B2(n90303), .A(n91257), .ZN(n91256) );
  AOI22_X1 U76805 ( .A1(n90305), .A2(n110945), .B1(n90306), .B2(n74407), .ZN(
        n91257) );
  NAND2_X1 U76806 ( .A1(n91258), .A2(n91259), .ZN(n91255) );
  AOI22_X1 U76807 ( .A1(n90309), .A2(n110950), .B1(n105653), .B2(n110947), 
        .ZN(n91259) );
  AOI22_X1 U76808 ( .A1(n90311), .A2(n74405), .B1(n90312), .B2(n110946), .ZN(
        n91258) );
  NOR4_X1 U76809 ( .A1(n91260), .A2(n91261), .A3(n91262), .A4(n91263), .ZN(
        n91253) );
  NAND2_X1 U76810 ( .A1(n91264), .A2(n91265), .ZN(n91263) );
  NOR4_X1 U76811 ( .A1(n91266), .A2(n91267), .A3(n91268), .A4(n91269), .ZN(
        n91265) );
  NAND2_X1 U76812 ( .A1(n91270), .A2(n91271), .ZN(n91269) );
  AOI22_X1 U76813 ( .A1(n90325), .A2(n110926), .B1(n90326), .B2(n110927), .ZN(
        n91271) );
  AOI22_X1 U76814 ( .A1(n90327), .A2(n110935), .B1(n90328), .B2(n110933), .ZN(
        n91270) );
  NAND2_X1 U76815 ( .A1(n91272), .A2(n91273), .ZN(n91268) );
  AOI22_X1 U76816 ( .A1(n90331), .A2(n74274), .B1(n90332), .B2(n110930), .ZN(
        n91273) );
  AOI22_X1 U76817 ( .A1(n90333), .A2(n74378), .B1(n90334), .B2(n110853), .ZN(
        n91272) );
  NAND2_X1 U76818 ( .A1(n91274), .A2(n91275), .ZN(n91267) );
  AOI22_X1 U76819 ( .A1(n90337), .A2(n110857), .B1(n90338), .B2(n74278), .ZN(
        n91275) );
  AOI22_X1 U76820 ( .A1(n90339), .A2(n110931), .B1(n90340), .B2(n110928), .ZN(
        n91274) );
  NAND2_X1 U76821 ( .A1(n91276), .A2(n91277), .ZN(n91266) );
  AOI22_X1 U76822 ( .A1(n90343), .A2(n110855), .B1(n90344), .B2(n110859), .ZN(
        n91277) );
  AOI22_X1 U76823 ( .A1(n90345), .A2(n110858), .B1(n90346), .B2(n74280), .ZN(
        n91276) );
  NOR4_X1 U76824 ( .A1(n91278), .A2(n91279), .A3(n91280), .A4(n91281), .ZN(
        n91264) );
  NAND2_X1 U76825 ( .A1(n91282), .A2(n91283), .ZN(n91281) );
  AOI22_X1 U76826 ( .A1(n90353), .A2(n110936), .B1(n90354), .B2(n110939), .ZN(
        n91283) );
  AOI22_X1 U76827 ( .A1(n90355), .A2(n110940), .B1(n90356), .B2(n110942), .ZN(
        n91282) );
  NAND2_X1 U76828 ( .A1(n91284), .A2(n91285), .ZN(n91280) );
  AOI22_X1 U76829 ( .A1(n90359), .A2(n110941), .B1(n90360), .B2(n110937), .ZN(
        n91285) );
  AOI22_X1 U76830 ( .A1(n90361), .A2(n110943), .B1(n90362), .B2(n110938), .ZN(
        n91284) );
  NAND2_X1 U76831 ( .A1(n91286), .A2(n91287), .ZN(n91279) );
  AOI22_X1 U76832 ( .A1(n90365), .A2(n74388), .B1(n90366), .B2(n74387), .ZN(
        n91287) );
  AOI22_X1 U76833 ( .A1(n90367), .A2(n74390), .B1(n90368), .B2(n110944), .ZN(
        n91286) );
  NAND2_X1 U76834 ( .A1(n91288), .A2(n91289), .ZN(n91278) );
  AOI22_X1 U76835 ( .A1(n90371), .A2(n110929), .B1(n90372), .B2(n110934), .ZN(
        n91289) );
  AOI22_X1 U76836 ( .A1(n90373), .A2(n74385), .B1(n90374), .B2(n110932), .ZN(
        n91288) );
  NAND2_X1 U76837 ( .A1(n91290), .A2(n91291), .ZN(n91262) );
  NOR4_X1 U76838 ( .A1(n91292), .A2(n91293), .A3(n91294), .A4(n91295), .ZN(
        n91291) );
  NAND2_X1 U76839 ( .A1(n91296), .A2(n91297), .ZN(n91295) );
  AOI22_X1 U76840 ( .A1(n90383), .A2(n110868), .B1(n90384), .B2(n110870), .ZN(
        n91297) );
  AOI22_X1 U76841 ( .A1(n90385), .A2(n74303), .B1(n90386), .B2(n110869), .ZN(
        n91296) );
  NAND2_X1 U76842 ( .A1(n91298), .A2(n91299), .ZN(n91294) );
  AOI22_X1 U76843 ( .A1(n90389), .A2(n74307), .B1(n90390), .B2(n74309), .ZN(
        n91299) );
  AOI22_X1 U76844 ( .A1(n90391), .A2(n110875), .B1(n90392), .B2(n110876), .ZN(
        n91298) );
  NAND2_X1 U76845 ( .A1(n91300), .A2(n91301), .ZN(n91293) );
  AOI22_X1 U76846 ( .A1(n90395), .A2(n110873), .B1(n90396), .B2(n110874), .ZN(
        n91301) );
  AOI22_X1 U76847 ( .A1(n90397), .A2(n110877), .B1(n90398), .B2(n74302), .ZN(
        n91300) );
  NAND2_X1 U76848 ( .A1(n91302), .A2(n91303), .ZN(n91292) );
  AOI22_X1 U76849 ( .A1(n90401), .A2(n110882), .B1(n90402), .B2(n74314), .ZN(
        n91303) );
  AOI22_X1 U76850 ( .A1(n90403), .A2(n110881), .B1(n90404), .B2(n74312), .ZN(
        n91302) );
  NOR4_X1 U76851 ( .A1(n91304), .A2(n91305), .A3(n91306), .A4(n91307), .ZN(
        n91290) );
  NAND2_X1 U76852 ( .A1(n91308), .A2(n91309), .ZN(n91307) );
  AOI22_X1 U76853 ( .A1(n90411), .A2(n110863), .B1(n90412), .B2(n110854), .ZN(
        n91309) );
  AOI22_X1 U76854 ( .A1(n90413), .A2(n110856), .B1(n90414), .B2(n74286), .ZN(
        n91308) );
  NAND2_X1 U76855 ( .A1(n91310), .A2(n91311), .ZN(n91306) );
  AOI22_X1 U76856 ( .A1(n90417), .A2(n110861), .B1(n90418), .B2(n110865), .ZN(
        n91311) );
  AOI22_X1 U76857 ( .A1(n90419), .A2(n110867), .B1(n90420), .B2(n110864), .ZN(
        n91310) );
  NAND2_X1 U76858 ( .A1(n91312), .A2(n91313), .ZN(n91305) );
  AOI22_X1 U76859 ( .A1(n90423), .A2(n74295), .B1(n90424), .B2(n110860), .ZN(
        n91313) );
  AOI22_X1 U76860 ( .A1(n90425), .A2(n110862), .B1(n90426), .B2(n110866), .ZN(
        n91312) );
  NAND2_X1 U76861 ( .A1(n91314), .A2(n91315), .ZN(n91304) );
  AOI22_X1 U76862 ( .A1(n90429), .A2(n110872), .B1(n90430), .B2(n74299), .ZN(
        n91315) );
  AOI22_X1 U76863 ( .A1(n90431), .A2(n74297), .B1(n90432), .B2(n110871), .ZN(
        n91314) );
  NAND2_X1 U76864 ( .A1(n91316), .A2(n91317), .ZN(n91261) );
  NOR4_X1 U76865 ( .A1(n91318), .A2(n91319), .A3(n91320), .A4(n91321), .ZN(
        n91317) );
  NAND2_X1 U76866 ( .A1(n91322), .A2(n91323), .ZN(n91321) );
  AOI22_X1 U76867 ( .A1(n90441), .A2(n74337), .B1(n90442), .B2(n110891), .ZN(
        n91323) );
  AOI22_X1 U76868 ( .A1(n90443), .A2(n110894), .B1(n90444), .B2(n110893), .ZN(
        n91322) );
  NAND2_X1 U76869 ( .A1(n91324), .A2(n91325), .ZN(n91320) );
  AOI22_X1 U76870 ( .A1(n90447), .A2(n110897), .B1(n90448), .B2(n110896), .ZN(
        n91325) );
  AOI22_X1 U76871 ( .A1(n90449), .A2(n110890), .B1(n90450), .B2(n111016), .ZN(
        n91324) );
  NAND2_X1 U76872 ( .A1(n91326), .A2(n91327), .ZN(n91319) );
  AOI22_X1 U76873 ( .A1(n90453), .A2(n74342), .B1(n90454), .B2(n74336), .ZN(
        n91327) );
  AOI22_X1 U76874 ( .A1(n90455), .A2(n74341), .B1(n90456), .B2(n74343), .ZN(
        n91326) );
  NAND2_X1 U76875 ( .A1(n91328), .A2(n91329), .ZN(n91318) );
  AOI22_X1 U76876 ( .A1(n90459), .A2(n111037), .B1(n90460), .B2(n74349), .ZN(
        n91329) );
  AOI22_X1 U76877 ( .A1(n90461), .A2(n110895), .B1(n90462), .B2(n74338), .ZN(
        n91328) );
  NOR4_X1 U76878 ( .A1(n91330), .A2(n91331), .A3(n91332), .A4(n91333), .ZN(
        n91316) );
  NAND2_X1 U76879 ( .A1(n91334), .A2(n91335), .ZN(n91333) );
  AOI22_X1 U76880 ( .A1(n90469), .A2(n110880), .B1(n90470), .B2(n110884), .ZN(
        n91335) );
  AOI22_X1 U76881 ( .A1(n90471), .A2(n110879), .B1(n90472), .B2(n74317), .ZN(
        n91334) );
  NAND2_X1 U76882 ( .A1(n91336), .A2(n91337), .ZN(n91332) );
  AOI22_X1 U76883 ( .A1(n90475), .A2(n74326), .B1(n90476), .B2(n110886), .ZN(
        n91337) );
  AOI22_X1 U76884 ( .A1(n90477), .A2(n110887), .B1(n90478), .B2(n110878), .ZN(
        n91336) );
  NAND2_X1 U76885 ( .A1(n91338), .A2(n91339), .ZN(n91331) );
  AOI22_X1 U76886 ( .A1(n90481), .A2(n110885), .B1(n90482), .B2(n110889), .ZN(
        n91339) );
  AOI22_X1 U76887 ( .A1(n90483), .A2(n74319), .B1(n90484), .B2(n110888), .ZN(
        n91338) );
  NAND2_X1 U76888 ( .A1(n91340), .A2(n91341), .ZN(n91330) );
  AOI22_X1 U76889 ( .A1(n90487), .A2(n74331), .B1(n90488), .B2(n110892), .ZN(
        n91341) );
  AOI22_X1 U76890 ( .A1(n90489), .A2(n74329), .B1(n90490), .B2(n110883), .ZN(
        n91340) );
  NAND2_X1 U76891 ( .A1(n91342), .A2(n91343), .ZN(n91260) );
  NOR4_X1 U76892 ( .A1(n91344), .A2(n91345), .A3(n91346), .A4(n91347), .ZN(
        n91343) );
  NAND2_X1 U76893 ( .A1(n91348), .A2(n91349), .ZN(n91347) );
  AOI22_X1 U76894 ( .A1(n90499), .A2(n110917), .B1(n90500), .B2(n110916), .ZN(
        n91349) );
  AOI22_X1 U76895 ( .A1(n90501), .A2(n74365), .B1(n90502), .B2(n110914), .ZN(
        n91348) );
  NAND2_X1 U76896 ( .A1(n91350), .A2(n91351), .ZN(n91346) );
  AOI22_X1 U76897 ( .A1(n90505), .A2(n110912), .B1(n90506), .B2(n110915), .ZN(
        n91351) );
  AOI22_X1 U76898 ( .A1(n90507), .A2(n74371), .B1(n90508), .B2(n110913), .ZN(
        n91350) );
  NAND2_X1 U76899 ( .A1(n91352), .A2(n91353), .ZN(n91345) );
  AOI22_X1 U76900 ( .A1(n105650), .A2(n110923), .B1(n90512), .B2(n74377), .ZN(
        n91353) );
  AOI22_X1 U76901 ( .A1(n90513), .A2(n110921), .B1(n90514), .B2(n110922), .ZN(
        n91352) );
  NAND2_X1 U76902 ( .A1(n91354), .A2(n91355), .ZN(n91344) );
  AOI22_X1 U76903 ( .A1(n90517), .A2(n110918), .B1(n90518), .B2(n110920), .ZN(
        n91355) );
  AOI22_X1 U76904 ( .A1(n90519), .A2(n110924), .B1(n105644), .B2(n110919), 
        .ZN(n91354) );
  NOR4_X1 U76905 ( .A1(n91356), .A2(n91357), .A3(n91358), .A4(n91359), .ZN(
        n91342) );
  NAND2_X1 U76906 ( .A1(n91360), .A2(n91361), .ZN(n91359) );
  AOI22_X1 U76907 ( .A1(n90527), .A2(n110899), .B1(n90528), .B2(n110902), .ZN(
        n91361) );
  AOI22_X1 U76908 ( .A1(n90529), .A2(n110901), .B1(n90530), .B2(n74348), .ZN(
        n91360) );
  NAND2_X1 U76909 ( .A1(n91362), .A2(n91363), .ZN(n91358) );
  AOI22_X1 U76910 ( .A1(n90533), .A2(n110908), .B1(n90534), .B2(n110898), .ZN(
        n91363) );
  AOI22_X1 U76911 ( .A1(n90535), .A2(n110900), .B1(n90536), .B2(n110905), .ZN(
        n91362) );
  NAND2_X1 U76912 ( .A1(n91364), .A2(n91365), .ZN(n91357) );
  AOI22_X1 U76913 ( .A1(n90539), .A2(n110904), .B1(n90540), .B2(n110909), .ZN(
        n91365) );
  AOI22_X1 U76914 ( .A1(n90541), .A2(n110911), .B1(n90542), .B2(n110907), .ZN(
        n91364) );
  NAND2_X1 U76915 ( .A1(n91366), .A2(n91367), .ZN(n91356) );
  AOI22_X1 U76916 ( .A1(n90545), .A2(n74366), .B1(n90546), .B2(n110903), .ZN(
        n91367) );
  AOI22_X1 U76917 ( .A1(n90547), .A2(n110906), .B1(n90548), .B2(n110910), .ZN(
        n91366) );
  AOI21_X1 U76918 ( .B1(n90295), .B2(n87384), .A(n91369), .ZN(n91368) );
  OAI21_X1 U76919 ( .B1(n91370), .B2(n105659), .A(n91371), .ZN(n91369) );
  OAI21_X1 U76920 ( .B1(n91372), .B2(n91373), .A(n90302), .ZN(n91371) );
  OAI21_X1 U76921 ( .B1(n102057), .B2(n90303), .A(n91374), .ZN(n91373) );
  AOI22_X1 U76922 ( .A1(n90305), .A2(n110538), .B1(n90306), .B2(n73843), .ZN(
        n91374) );
  NAND2_X1 U76923 ( .A1(n91375), .A2(n91376), .ZN(n91372) );
  AOI22_X1 U76924 ( .A1(n90309), .A2(n110543), .B1(n105653), .B2(n110540), 
        .ZN(n91376) );
  AOI22_X1 U76925 ( .A1(n90311), .A2(n73841), .B1(n90312), .B2(n110539), .ZN(
        n91375) );
  NOR4_X1 U76926 ( .A1(n91377), .A2(n91378), .A3(n91379), .A4(n91380), .ZN(
        n91370) );
  NAND2_X1 U76927 ( .A1(n91381), .A2(n91382), .ZN(n91380) );
  NOR4_X1 U76928 ( .A1(n91383), .A2(n91384), .A3(n91385), .A4(n91386), .ZN(
        n91382) );
  NAND2_X1 U76929 ( .A1(n91387), .A2(n91388), .ZN(n91386) );
  AOI22_X1 U76930 ( .A1(n90325), .A2(n110519), .B1(n90326), .B2(n110520), .ZN(
        n91388) );
  AOI22_X1 U76931 ( .A1(n90327), .A2(n110528), .B1(n90328), .B2(n110526), .ZN(
        n91387) );
  NAND2_X1 U76932 ( .A1(n91389), .A2(n91390), .ZN(n91385) );
  AOI22_X1 U76933 ( .A1(n90331), .A2(n73710), .B1(n90332), .B2(n110523), .ZN(
        n91390) );
  AOI22_X1 U76934 ( .A1(n90333), .A2(n73814), .B1(n90334), .B2(n110448), .ZN(
        n91389) );
  NAND2_X1 U76935 ( .A1(n91391), .A2(n91392), .ZN(n91384) );
  AOI22_X1 U76936 ( .A1(n90337), .A2(n110452), .B1(n90338), .B2(n73714), .ZN(
        n91392) );
  AOI22_X1 U76937 ( .A1(n90339), .A2(n110524), .B1(n90340), .B2(n110521), .ZN(
        n91391) );
  NAND2_X1 U76938 ( .A1(n91393), .A2(n91394), .ZN(n91383) );
  AOI22_X1 U76939 ( .A1(n90343), .A2(n110450), .B1(n90344), .B2(n110454), .ZN(
        n91394) );
  AOI22_X1 U76940 ( .A1(n90345), .A2(n110453), .B1(n90346), .B2(n73716), .ZN(
        n91393) );
  NOR4_X1 U76941 ( .A1(n91395), .A2(n91396), .A3(n91397), .A4(n91398), .ZN(
        n91381) );
  NAND2_X1 U76942 ( .A1(n91399), .A2(n91400), .ZN(n91398) );
  AOI22_X1 U76943 ( .A1(n90353), .A2(n110529), .B1(n90354), .B2(n110532), .ZN(
        n91400) );
  AOI22_X1 U76944 ( .A1(n90355), .A2(n110533), .B1(n90356), .B2(n110535), .ZN(
        n91399) );
  NAND2_X1 U76945 ( .A1(n91401), .A2(n91402), .ZN(n91397) );
  AOI22_X1 U76946 ( .A1(n90359), .A2(n110534), .B1(n90360), .B2(n110530), .ZN(
        n91402) );
  AOI22_X1 U76947 ( .A1(n90361), .A2(n110536), .B1(n90362), .B2(n110531), .ZN(
        n91401) );
  NAND2_X1 U76948 ( .A1(n91403), .A2(n91404), .ZN(n91396) );
  AOI22_X1 U76949 ( .A1(n90365), .A2(n73824), .B1(n90366), .B2(n73823), .ZN(
        n91404) );
  AOI22_X1 U76950 ( .A1(n90367), .A2(n73826), .B1(n90368), .B2(n110537), .ZN(
        n91403) );
  NAND2_X1 U76951 ( .A1(n91405), .A2(n91406), .ZN(n91395) );
  AOI22_X1 U76952 ( .A1(n90371), .A2(n110522), .B1(n90372), .B2(n110527), .ZN(
        n91406) );
  AOI22_X1 U76953 ( .A1(n90373), .A2(n73821), .B1(n90374), .B2(n110525), .ZN(
        n91405) );
  NAND2_X1 U76954 ( .A1(n91407), .A2(n91408), .ZN(n91379) );
  NOR4_X1 U76955 ( .A1(n91409), .A2(n91410), .A3(n91411), .A4(n91412), .ZN(
        n91408) );
  NAND2_X1 U76956 ( .A1(n91413), .A2(n91414), .ZN(n91412) );
  AOI22_X1 U76957 ( .A1(n90383), .A2(n110463), .B1(n90384), .B2(n110465), .ZN(
        n91414) );
  AOI22_X1 U76958 ( .A1(n90385), .A2(n73739), .B1(n90386), .B2(n110464), .ZN(
        n91413) );
  NAND2_X1 U76959 ( .A1(n91415), .A2(n91416), .ZN(n91411) );
  AOI22_X1 U76960 ( .A1(n90389), .A2(n73743), .B1(n90390), .B2(n73745), .ZN(
        n91416) );
  AOI22_X1 U76961 ( .A1(n90391), .A2(n110470), .B1(n90392), .B2(n110471), .ZN(
        n91415) );
  NAND2_X1 U76962 ( .A1(n91417), .A2(n91418), .ZN(n91410) );
  AOI22_X1 U76963 ( .A1(n90395), .A2(n110468), .B1(n90396), .B2(n110469), .ZN(
        n91418) );
  AOI22_X1 U76964 ( .A1(n90397), .A2(n73744), .B1(n90398), .B2(n73738), .ZN(
        n91417) );
  NAND2_X1 U76965 ( .A1(n91419), .A2(n91420), .ZN(n91409) );
  AOI22_X1 U76966 ( .A1(n90401), .A2(n110476), .B1(n90402), .B2(n73750), .ZN(
        n91420) );
  AOI22_X1 U76967 ( .A1(n90403), .A2(n110475), .B1(n90404), .B2(n73748), .ZN(
        n91419) );
  NOR4_X1 U76968 ( .A1(n91421), .A2(n91422), .A3(n91423), .A4(n91424), .ZN(
        n91407) );
  NAND2_X1 U76969 ( .A1(n91425), .A2(n91426), .ZN(n91424) );
  AOI22_X1 U76970 ( .A1(n90411), .A2(n110458), .B1(n90412), .B2(n110449), .ZN(
        n91426) );
  AOI22_X1 U76971 ( .A1(n90413), .A2(n110451), .B1(n90414), .B2(n73722), .ZN(
        n91425) );
  NAND2_X1 U76972 ( .A1(n91427), .A2(n91428), .ZN(n91423) );
  AOI22_X1 U76973 ( .A1(n90417), .A2(n110456), .B1(n90418), .B2(n110460), .ZN(
        n91428) );
  AOI22_X1 U76974 ( .A1(n90419), .A2(n110462), .B1(n90420), .B2(n110459), .ZN(
        n91427) );
  NAND2_X1 U76975 ( .A1(n91429), .A2(n91430), .ZN(n91422) );
  AOI22_X1 U76976 ( .A1(n90423), .A2(n73731), .B1(n90424), .B2(n110455), .ZN(
        n91430) );
  AOI22_X1 U76977 ( .A1(n90425), .A2(n110457), .B1(n90426), .B2(n110461), .ZN(
        n91429) );
  NAND2_X1 U76978 ( .A1(n91431), .A2(n91432), .ZN(n91421) );
  AOI22_X1 U76979 ( .A1(n90429), .A2(n110467), .B1(n90430), .B2(n73735), .ZN(
        n91432) );
  AOI22_X1 U76980 ( .A1(n90431), .A2(n73733), .B1(n90432), .B2(n110466), .ZN(
        n91431) );
  NAND2_X1 U76981 ( .A1(n91433), .A2(n91434), .ZN(n91378) );
  NOR4_X1 U76982 ( .A1(n91435), .A2(n91436), .A3(n91437), .A4(n91438), .ZN(
        n91434) );
  NAND2_X1 U76983 ( .A1(n91439), .A2(n91440), .ZN(n91438) );
  AOI22_X1 U76984 ( .A1(n90441), .A2(n73773), .B1(n90442), .B2(n110485), .ZN(
        n91440) );
  AOI22_X1 U76985 ( .A1(n90443), .A2(n110488), .B1(n90444), .B2(n110487), .ZN(
        n91439) );
  NAND2_X1 U76986 ( .A1(n91441), .A2(n91442), .ZN(n91437) );
  AOI22_X1 U76987 ( .A1(n90447), .A2(n110492), .B1(n90448), .B2(n110491), .ZN(
        n91442) );
  AOI22_X1 U76988 ( .A1(n90449), .A2(n110484), .B1(n90450), .B2(n111017), .ZN(
        n91441) );
  NAND2_X1 U76989 ( .A1(n91443), .A2(n91444), .ZN(n91436) );
  AOI22_X1 U76990 ( .A1(n90453), .A2(n110493), .B1(n90454), .B2(n73772), .ZN(
        n91444) );
  AOI22_X1 U76991 ( .A1(n90455), .A2(n73777), .B1(n90456), .B2(n73779), .ZN(
        n91443) );
  NAND2_X1 U76992 ( .A1(n91445), .A2(n91446), .ZN(n91435) );
  AOI22_X1 U76993 ( .A1(n90459), .A2(n111036), .B1(n90460), .B2(n73785), .ZN(
        n91446) );
  AOI22_X1 U76994 ( .A1(n90461), .A2(n110489), .B1(n90462), .B2(n110490), .ZN(
        n91445) );
  NOR4_X1 U76995 ( .A1(n91447), .A2(n91448), .A3(n91449), .A4(n91450), .ZN(
        n91433) );
  NAND2_X1 U76996 ( .A1(n91451), .A2(n91452), .ZN(n91450) );
  AOI22_X1 U76997 ( .A1(n90469), .A2(n110474), .B1(n90470), .B2(n110479), .ZN(
        n91452) );
  AOI22_X1 U76998 ( .A1(n90471), .A2(n110473), .B1(n90472), .B2(n73753), .ZN(
        n91451) );
  NAND2_X1 U76999 ( .A1(n91453), .A2(n91454), .ZN(n91449) );
  AOI22_X1 U77000 ( .A1(n90475), .A2(n73762), .B1(n90476), .B2(n110480), .ZN(
        n91454) );
  AOI22_X1 U77001 ( .A1(n90477), .A2(n110481), .B1(n90478), .B2(n110472), .ZN(
        n91453) );
  NAND2_X1 U77002 ( .A1(n91455), .A2(n91456), .ZN(n91448) );
  AOI22_X1 U77003 ( .A1(n90481), .A2(n73757), .B1(n90482), .B2(n110483), .ZN(
        n91456) );
  AOI22_X1 U77004 ( .A1(n90483), .A2(n110478), .B1(n90484), .B2(n110482), .ZN(
        n91455) );
  NAND2_X1 U77005 ( .A1(n91457), .A2(n91458), .ZN(n91447) );
  AOI22_X1 U77006 ( .A1(n90487), .A2(n73767), .B1(n90488), .B2(n110486), .ZN(
        n91458) );
  AOI22_X1 U77007 ( .A1(n90489), .A2(n73765), .B1(n90490), .B2(n110477), .ZN(
        n91457) );
  NAND2_X1 U77008 ( .A1(n91459), .A2(n91460), .ZN(n91377) );
  NOR4_X1 U77009 ( .A1(n91461), .A2(n91462), .A3(n91463), .A4(n91464), .ZN(
        n91460) );
  NAND2_X1 U77010 ( .A1(n91465), .A2(n91466), .ZN(n91464) );
  AOI22_X1 U77011 ( .A1(n90499), .A2(n110512), .B1(n90500), .B2(n110511), .ZN(
        n91466) );
  AOI22_X1 U77012 ( .A1(n90501), .A2(n73801), .B1(n90502), .B2(n110509), .ZN(
        n91465) );
  NAND2_X1 U77013 ( .A1(n91467), .A2(n91468), .ZN(n91463) );
  AOI22_X1 U77014 ( .A1(n90505), .A2(n110507), .B1(n90506), .B2(n110510), .ZN(
        n91468) );
  AOI22_X1 U77015 ( .A1(n90507), .A2(n73807), .B1(n90508), .B2(n110508), .ZN(
        n91467) );
  NAND2_X1 U77016 ( .A1(n91469), .A2(n91470), .ZN(n91462) );
  AOI22_X1 U77017 ( .A1(n105650), .A2(n110517), .B1(n90512), .B2(n73813), .ZN(
        n91470) );
  AOI22_X1 U77018 ( .A1(n90513), .A2(n110515), .B1(n90514), .B2(n110516), .ZN(
        n91469) );
  NAND2_X1 U77019 ( .A1(n91471), .A2(n91472), .ZN(n91461) );
  AOI22_X1 U77020 ( .A1(n90517), .A2(n73805), .B1(n90518), .B2(n110514), .ZN(
        n91472) );
  AOI22_X1 U77021 ( .A1(n90519), .A2(n73812), .B1(n90520), .B2(n110513), .ZN(
        n91471) );
  NOR4_X1 U77022 ( .A1(n91473), .A2(n91474), .A3(n91475), .A4(n91476), .ZN(
        n91459) );
  NAND2_X1 U77023 ( .A1(n91477), .A2(n91478), .ZN(n91476) );
  AOI22_X1 U77024 ( .A1(n90527), .A2(n110494), .B1(n90528), .B2(n110497), .ZN(
        n91478) );
  AOI22_X1 U77025 ( .A1(n90529), .A2(n110496), .B1(n90530), .B2(n73784), .ZN(
        n91477) );
  NAND2_X1 U77026 ( .A1(n91479), .A2(n91480), .ZN(n91475) );
  AOI22_X1 U77027 ( .A1(n90533), .A2(n110503), .B1(n90534), .B2(n73780), .ZN(
        n91480) );
  AOI22_X1 U77028 ( .A1(n90535), .A2(n110495), .B1(n90536), .B2(n110500), .ZN(
        n91479) );
  NAND2_X1 U77029 ( .A1(n91481), .A2(n91482), .ZN(n91474) );
  AOI22_X1 U77030 ( .A1(n90539), .A2(n110499), .B1(n90540), .B2(n110504), .ZN(
        n91482) );
  AOI22_X1 U77031 ( .A1(n90541), .A2(n110506), .B1(n90542), .B2(n110502), .ZN(
        n91481) );
  NAND2_X1 U77032 ( .A1(n91483), .A2(n91484), .ZN(n91473) );
  AOI22_X1 U77033 ( .A1(n90545), .A2(n73802), .B1(n90546), .B2(n110498), .ZN(
        n91484) );
  AOI22_X1 U77034 ( .A1(n90547), .A2(n110501), .B1(n90548), .B2(n110505), .ZN(
        n91483) );
  AOI21_X1 U77035 ( .B1(n90295), .B2(n87502), .A(n91486), .ZN(n91485) );
  OAI21_X1 U77036 ( .B1(n91487), .B2(n105659), .A(n91488), .ZN(n91486) );
  OAI21_X1 U77037 ( .B1(n91489), .B2(n91490), .A(n90302), .ZN(n91488) );
  OAI21_X1 U77038 ( .B1(n102041), .B2(n90303), .A(n91491), .ZN(n91490) );
  AOI22_X1 U77039 ( .A1(n90305), .A2(n110323), .B1(n90306), .B2(n73547), .ZN(
        n91491) );
  NAND2_X1 U77040 ( .A1(n91492), .A2(n91493), .ZN(n91489) );
  AOI22_X1 U77041 ( .A1(n90309), .A2(n110328), .B1(n105653), .B2(n110325), 
        .ZN(n91493) );
  AOI22_X1 U77042 ( .A1(n90311), .A2(n73545), .B1(n90312), .B2(n110324), .ZN(
        n91492) );
  NOR4_X1 U77043 ( .A1(n91494), .A2(n91495), .A3(n91496), .A4(n91497), .ZN(
        n91487) );
  NAND2_X1 U77044 ( .A1(n91498), .A2(n91499), .ZN(n91497) );
  NOR4_X1 U77045 ( .A1(n91500), .A2(n91501), .A3(n91502), .A4(n91503), .ZN(
        n91499) );
  NAND2_X1 U77046 ( .A1(n91504), .A2(n91505), .ZN(n91503) );
  AOI22_X1 U77047 ( .A1(n90325), .A2(n110304), .B1(n90326), .B2(n110305), .ZN(
        n91505) );
  AOI22_X1 U77048 ( .A1(n90327), .A2(n110313), .B1(n90328), .B2(n110311), .ZN(
        n91504) );
  NAND2_X1 U77049 ( .A1(n91506), .A2(n91507), .ZN(n91502) );
  AOI22_X1 U77050 ( .A1(n90331), .A2(n73414), .B1(n90332), .B2(n110308), .ZN(
        n91507) );
  AOI22_X1 U77051 ( .A1(n90333), .A2(n73518), .B1(n90334), .B2(n110231), .ZN(
        n91506) );
  NAND2_X1 U77052 ( .A1(n91508), .A2(n91509), .ZN(n91501) );
  AOI22_X1 U77053 ( .A1(n90337), .A2(n110234), .B1(n90338), .B2(n73418), .ZN(
        n91509) );
  AOI22_X1 U77054 ( .A1(n90339), .A2(n110309), .B1(n90340), .B2(n110306), .ZN(
        n91508) );
  NAND2_X1 U77055 ( .A1(n91510), .A2(n91511), .ZN(n91500) );
  AOI22_X1 U77056 ( .A1(n90343), .A2(n110232), .B1(n90344), .B2(n110236), .ZN(
        n91511) );
  AOI22_X1 U77057 ( .A1(n90345), .A2(n110235), .B1(n90346), .B2(n73420), .ZN(
        n91510) );
  NOR4_X1 U77058 ( .A1(n91512), .A2(n91513), .A3(n91514), .A4(n91515), .ZN(
        n91498) );
  NAND2_X1 U77059 ( .A1(n91516), .A2(n91517), .ZN(n91515) );
  AOI22_X1 U77060 ( .A1(n90353), .A2(n110314), .B1(n90354), .B2(n110317), .ZN(
        n91517) );
  AOI22_X1 U77061 ( .A1(n90355), .A2(n110318), .B1(n90356), .B2(n110320), .ZN(
        n91516) );
  NAND2_X1 U77062 ( .A1(n91518), .A2(n91519), .ZN(n91514) );
  AOI22_X1 U77063 ( .A1(n90359), .A2(n110319), .B1(n90360), .B2(n110315), .ZN(
        n91519) );
  AOI22_X1 U77064 ( .A1(n90361), .A2(n110321), .B1(n90362), .B2(n110316), .ZN(
        n91518) );
  NAND2_X1 U77065 ( .A1(n91520), .A2(n91521), .ZN(n91513) );
  AOI22_X1 U77066 ( .A1(n90365), .A2(n73528), .B1(n90366), .B2(n73527), .ZN(
        n91521) );
  AOI22_X1 U77067 ( .A1(n90367), .A2(n73530), .B1(n90368), .B2(n110322), .ZN(
        n91520) );
  NAND2_X1 U77068 ( .A1(n91522), .A2(n91523), .ZN(n91512) );
  AOI22_X1 U77069 ( .A1(n90371), .A2(n110307), .B1(n90372), .B2(n110312), .ZN(
        n91523) );
  AOI22_X1 U77070 ( .A1(n90373), .A2(n73525), .B1(n90374), .B2(n110310), .ZN(
        n91522) );
  NAND2_X1 U77071 ( .A1(n91524), .A2(n91525), .ZN(n91496) );
  NOR4_X1 U77072 ( .A1(n91526), .A2(n91527), .A3(n91528), .A4(n91529), .ZN(
        n91525) );
  NAND2_X1 U77073 ( .A1(n91530), .A2(n91531), .ZN(n91529) );
  AOI22_X1 U77074 ( .A1(n90383), .A2(n110245), .B1(n90384), .B2(n110247), .ZN(
        n91531) );
  AOI22_X1 U77075 ( .A1(n90385), .A2(n73443), .B1(n90386), .B2(n110246), .ZN(
        n91530) );
  NAND2_X1 U77076 ( .A1(n91532), .A2(n91533), .ZN(n91528) );
  AOI22_X1 U77077 ( .A1(n90389), .A2(n73447), .B1(n90390), .B2(n73449), .ZN(
        n91533) );
  AOI22_X1 U77078 ( .A1(n90391), .A2(n110252), .B1(n90392), .B2(n110253), .ZN(
        n91532) );
  NAND2_X1 U77079 ( .A1(n91534), .A2(n91535), .ZN(n91527) );
  AOI22_X1 U77080 ( .A1(n90395), .A2(n110250), .B1(n90396), .B2(n110251), .ZN(
        n91535) );
  AOI22_X1 U77081 ( .A1(n90397), .A2(n73448), .B1(n90398), .B2(n73442), .ZN(
        n91534) );
  NAND2_X1 U77082 ( .A1(n91536), .A2(n91537), .ZN(n91526) );
  AOI22_X1 U77083 ( .A1(n90401), .A2(n110258), .B1(n90402), .B2(n73454), .ZN(
        n91537) );
  AOI22_X1 U77084 ( .A1(n90403), .A2(n110257), .B1(n90404), .B2(n73452), .ZN(
        n91536) );
  NOR4_X1 U77085 ( .A1(n91538), .A2(n91539), .A3(n91540), .A4(n91541), .ZN(
        n91524) );
  NAND2_X1 U77086 ( .A1(n91542), .A2(n91543), .ZN(n91541) );
  AOI22_X1 U77087 ( .A1(n90411), .A2(n110240), .B1(n90412), .B2(n111020), .ZN(
        n91543) );
  AOI22_X1 U77088 ( .A1(n90413), .A2(n110233), .B1(n90414), .B2(n73426), .ZN(
        n91542) );
  NAND2_X1 U77089 ( .A1(n91544), .A2(n91545), .ZN(n91540) );
  AOI22_X1 U77090 ( .A1(n90417), .A2(n110238), .B1(n90418), .B2(n110242), .ZN(
        n91545) );
  AOI22_X1 U77091 ( .A1(n90419), .A2(n110244), .B1(n90420), .B2(n110241), .ZN(
        n91544) );
  NAND2_X1 U77092 ( .A1(n91546), .A2(n91547), .ZN(n91539) );
  AOI22_X1 U77093 ( .A1(n90423), .A2(n73435), .B1(n90424), .B2(n110237), .ZN(
        n91547) );
  AOI22_X1 U77094 ( .A1(n90425), .A2(n110239), .B1(n90426), .B2(n110243), .ZN(
        n91546) );
  NAND2_X1 U77095 ( .A1(n91548), .A2(n91549), .ZN(n91538) );
  AOI22_X1 U77096 ( .A1(n90429), .A2(n110249), .B1(n90430), .B2(n73439), .ZN(
        n91549) );
  AOI22_X1 U77097 ( .A1(n90431), .A2(n73437), .B1(n90432), .B2(n110248), .ZN(
        n91548) );
  NAND2_X1 U77098 ( .A1(n91550), .A2(n91551), .ZN(n91495) );
  NOR4_X1 U77099 ( .A1(n91552), .A2(n91553), .A3(n91554), .A4(n91555), .ZN(
        n91551) );
  NAND2_X1 U77100 ( .A1(n91556), .A2(n91557), .ZN(n91555) );
  AOI22_X1 U77101 ( .A1(n90441), .A2(n73477), .B1(n90442), .B2(n110267), .ZN(
        n91557) );
  AOI22_X1 U77102 ( .A1(n90443), .A2(n110271), .B1(n90444), .B2(n110270), .ZN(
        n91556) );
  NAND2_X1 U77103 ( .A1(n91558), .A2(n91559), .ZN(n91554) );
  AOI22_X1 U77104 ( .A1(n90447), .A2(n110275), .B1(n90448), .B2(n110274), .ZN(
        n91559) );
  AOI22_X1 U77105 ( .A1(n90449), .A2(n110266), .B1(n90450), .B2(n110268), .ZN(
        n91558) );
  NAND2_X1 U77106 ( .A1(n91560), .A2(n91561), .ZN(n91553) );
  AOI22_X1 U77107 ( .A1(n90453), .A2(n110276), .B1(n90454), .B2(n73476), .ZN(
        n91561) );
  AOI22_X1 U77108 ( .A1(n90455), .A2(n73481), .B1(n90456), .B2(n73483), .ZN(
        n91560) );
  NAND2_X1 U77109 ( .A1(n91562), .A2(n91563), .ZN(n91552) );
  AOI22_X1 U77110 ( .A1(n90459), .A2(n110278), .B1(n90460), .B2(n73489), .ZN(
        n91563) );
  AOI22_X1 U77111 ( .A1(n90461), .A2(n110272), .B1(n90462), .B2(n110273), .ZN(
        n91562) );
  NOR4_X1 U77112 ( .A1(n91564), .A2(n91565), .A3(n91566), .A4(n91567), .ZN(
        n91550) );
  NAND2_X1 U77113 ( .A1(n91568), .A2(n91569), .ZN(n91567) );
  AOI22_X1 U77114 ( .A1(n90469), .A2(n110256), .B1(n90470), .B2(n110261), .ZN(
        n91569) );
  AOI22_X1 U77115 ( .A1(n90471), .A2(n110255), .B1(n90472), .B2(n73457), .ZN(
        n91568) );
  NAND2_X1 U77116 ( .A1(n91570), .A2(n91571), .ZN(n91566) );
  AOI22_X1 U77117 ( .A1(n90475), .A2(n73466), .B1(n90476), .B2(n110262), .ZN(
        n91571) );
  AOI22_X1 U77118 ( .A1(n90477), .A2(n110263), .B1(n90478), .B2(n110254), .ZN(
        n91570) );
  NAND2_X1 U77119 ( .A1(n91572), .A2(n91573), .ZN(n91565) );
  AOI22_X1 U77120 ( .A1(n90481), .A2(n73461), .B1(n90482), .B2(n110265), .ZN(
        n91573) );
  AOI22_X1 U77121 ( .A1(n90483), .A2(n110260), .B1(n90484), .B2(n110264), .ZN(
        n91572) );
  NAND2_X1 U77122 ( .A1(n91574), .A2(n91575), .ZN(n91564) );
  AOI22_X1 U77123 ( .A1(n90487), .A2(n73471), .B1(n90488), .B2(n110269), .ZN(
        n91575) );
  AOI22_X1 U77124 ( .A1(n90489), .A2(n73469), .B1(n90490), .B2(n110259), .ZN(
        n91574) );
  NAND2_X1 U77125 ( .A1(n91576), .A2(n91577), .ZN(n91494) );
  NOR4_X1 U77126 ( .A1(n91578), .A2(n91579), .A3(n91580), .A4(n91581), .ZN(
        n91577) );
  NAND2_X1 U77127 ( .A1(n91582), .A2(n91583), .ZN(n91581) );
  AOI22_X1 U77128 ( .A1(n90499), .A2(n110295), .B1(n90500), .B2(n110294), .ZN(
        n91583) );
  AOI22_X1 U77129 ( .A1(n90501), .A2(n73505), .B1(n90502), .B2(n110292), .ZN(
        n91582) );
  NAND2_X1 U77130 ( .A1(n91584), .A2(n91585), .ZN(n91580) );
  AOI22_X1 U77131 ( .A1(n90505), .A2(n110290), .B1(n90506), .B2(n110293), .ZN(
        n91585) );
  AOI22_X1 U77132 ( .A1(n90507), .A2(n73511), .B1(n90508), .B2(n110291), .ZN(
        n91584) );
  NAND2_X1 U77133 ( .A1(n91586), .A2(n91587), .ZN(n91579) );
  AOI22_X1 U77134 ( .A1(n105650), .A2(n110301), .B1(n90512), .B2(n73517), .ZN(
        n91587) );
  AOI22_X1 U77135 ( .A1(n90513), .A2(n110299), .B1(n90514), .B2(n110300), .ZN(
        n91586) );
  NAND2_X1 U77136 ( .A1(n91588), .A2(n91589), .ZN(n91578) );
  AOI22_X1 U77137 ( .A1(n90517), .A2(n110296), .B1(n90518), .B2(n110298), .ZN(
        n91589) );
  AOI22_X1 U77138 ( .A1(n90519), .A2(n110302), .B1(n90520), .B2(n110297), .ZN(
        n91588) );
  NOR4_X1 U77139 ( .A1(n91590), .A2(n91591), .A3(n91592), .A4(n91593), .ZN(
        n91576) );
  NAND2_X1 U77140 ( .A1(n91594), .A2(n91595), .ZN(n91593) );
  AOI22_X1 U77141 ( .A1(n90527), .A2(n110277), .B1(n90528), .B2(n110280), .ZN(
        n91595) );
  AOI22_X1 U77142 ( .A1(n90529), .A2(n111039), .B1(n90530), .B2(n73488), .ZN(
        n91594) );
  NAND2_X1 U77143 ( .A1(n91596), .A2(n91597), .ZN(n91592) );
  AOI22_X1 U77144 ( .A1(n90533), .A2(n110286), .B1(n90534), .B2(n73484), .ZN(
        n91597) );
  AOI22_X1 U77145 ( .A1(n90535), .A2(n110279), .B1(n90536), .B2(n110283), .ZN(
        n91596) );
  NAND2_X1 U77146 ( .A1(n91598), .A2(n91599), .ZN(n91591) );
  AOI22_X1 U77147 ( .A1(n90539), .A2(n110282), .B1(n90540), .B2(n110287), .ZN(
        n91599) );
  AOI22_X1 U77148 ( .A1(n90541), .A2(n110289), .B1(n90542), .B2(n110285), .ZN(
        n91598) );
  NAND2_X1 U77149 ( .A1(n91600), .A2(n91601), .ZN(n91590) );
  AOI22_X1 U77150 ( .A1(n90545), .A2(n73506), .B1(n90546), .B2(n110281), .ZN(
        n91601) );
  AOI22_X1 U77151 ( .A1(n90547), .A2(n110284), .B1(n90548), .B2(n110288), .ZN(
        n91600) );
  AOI21_X1 U77152 ( .B1(n90295), .B2(n87620), .A(n91603), .ZN(n91602) );
  OAI21_X1 U77153 ( .B1(n91604), .B2(n105659), .A(n91605), .ZN(n91603) );
  OAI21_X1 U77154 ( .B1(n91606), .B2(n91607), .A(n90302), .ZN(n91605) );
  OAI21_X1 U77155 ( .B1(n102024), .B2(n90303), .A(n91608), .ZN(n91607) );
  AOI22_X1 U77156 ( .A1(n90305), .A2(n110643), .B1(n90306), .B2(n73984), .ZN(
        n91608) );
  NAND2_X1 U77157 ( .A1(n91609), .A2(n91610), .ZN(n91606) );
  AOI22_X1 U77158 ( .A1(n90309), .A2(n110648), .B1(n105653), .B2(n110645), 
        .ZN(n91610) );
  AOI22_X1 U77159 ( .A1(n90311), .A2(n73982), .B1(n90312), .B2(n110644), .ZN(
        n91609) );
  NOR4_X1 U77160 ( .A1(n91611), .A2(n91612), .A3(n91613), .A4(n91614), .ZN(
        n91604) );
  NAND2_X1 U77161 ( .A1(n91615), .A2(n91616), .ZN(n91614) );
  NOR4_X1 U77162 ( .A1(n91617), .A2(n91618), .A3(n91619), .A4(n91620), .ZN(
        n91616) );
  NAND2_X1 U77163 ( .A1(n91621), .A2(n91622), .ZN(n91620) );
  AOI22_X1 U77164 ( .A1(n90325), .A2(n110624), .B1(n90326), .B2(n110625), .ZN(
        n91622) );
  AOI22_X1 U77165 ( .A1(n90327), .A2(n110633), .B1(n90328), .B2(n110631), .ZN(
        n91621) );
  NAND2_X1 U77166 ( .A1(n91623), .A2(n91624), .ZN(n91619) );
  AOI22_X1 U77167 ( .A1(n90331), .A2(n73851), .B1(n90332), .B2(n110628), .ZN(
        n91624) );
  AOI22_X1 U77168 ( .A1(n90333), .A2(n73955), .B1(n90334), .B2(n110548), .ZN(
        n91623) );
  NAND2_X1 U77169 ( .A1(n91625), .A2(n91626), .ZN(n91618) );
  AOI22_X1 U77170 ( .A1(n90337), .A2(n110551), .B1(n90338), .B2(n73855), .ZN(
        n91626) );
  AOI22_X1 U77171 ( .A1(n90339), .A2(n110629), .B1(n90340), .B2(n110626), .ZN(
        n91625) );
  NAND2_X1 U77172 ( .A1(n91627), .A2(n91628), .ZN(n91617) );
  AOI22_X1 U77173 ( .A1(n90343), .A2(n110549), .B1(n90344), .B2(n110553), .ZN(
        n91628) );
  AOI22_X1 U77174 ( .A1(n90345), .A2(n110552), .B1(n90346), .B2(n73857), .ZN(
        n91627) );
  NOR4_X1 U77175 ( .A1(n91629), .A2(n91630), .A3(n91631), .A4(n91632), .ZN(
        n91615) );
  NAND2_X1 U77176 ( .A1(n91633), .A2(n91634), .ZN(n91632) );
  AOI22_X1 U77177 ( .A1(n90353), .A2(n110634), .B1(n90354), .B2(n110637), .ZN(
        n91634) );
  AOI22_X1 U77178 ( .A1(n90355), .A2(n110638), .B1(n90356), .B2(n110640), .ZN(
        n91633) );
  NAND2_X1 U77179 ( .A1(n91635), .A2(n91636), .ZN(n91631) );
  AOI22_X1 U77180 ( .A1(n90359), .A2(n110639), .B1(n90360), .B2(n110635), .ZN(
        n91636) );
  AOI22_X1 U77181 ( .A1(n90361), .A2(n110641), .B1(n90362), .B2(n110636), .ZN(
        n91635) );
  NAND2_X1 U77182 ( .A1(n91637), .A2(n91638), .ZN(n91630) );
  AOI22_X1 U77183 ( .A1(n90365), .A2(n73965), .B1(n90366), .B2(n73964), .ZN(
        n91638) );
  AOI22_X1 U77184 ( .A1(n90367), .A2(n73967), .B1(n90368), .B2(n110642), .ZN(
        n91637) );
  NAND2_X1 U77185 ( .A1(n91639), .A2(n91640), .ZN(n91629) );
  AOI22_X1 U77186 ( .A1(n90371), .A2(n110627), .B1(n90372), .B2(n110632), .ZN(
        n91640) );
  AOI22_X1 U77187 ( .A1(n90373), .A2(n73962), .B1(n90374), .B2(n110630), .ZN(
        n91639) );
  NAND2_X1 U77188 ( .A1(n91641), .A2(n91642), .ZN(n91613) );
  NOR4_X1 U77189 ( .A1(n91643), .A2(n91644), .A3(n91645), .A4(n91646), .ZN(
        n91642) );
  NAND2_X1 U77190 ( .A1(n91647), .A2(n91648), .ZN(n91646) );
  AOI22_X1 U77191 ( .A1(n90383), .A2(n110562), .B1(n90384), .B2(n110564), .ZN(
        n91648) );
  AOI22_X1 U77192 ( .A1(n90385), .A2(n73880), .B1(n90386), .B2(n110563), .ZN(
        n91647) );
  NAND2_X1 U77193 ( .A1(n91649), .A2(n91650), .ZN(n91645) );
  AOI22_X1 U77194 ( .A1(n90389), .A2(n73884), .B1(n90390), .B2(n73886), .ZN(
        n91650) );
  AOI22_X1 U77195 ( .A1(n90391), .A2(n110569), .B1(n90392), .B2(n110570), .ZN(
        n91649) );
  NAND2_X1 U77196 ( .A1(n91651), .A2(n91652), .ZN(n91644) );
  AOI22_X1 U77197 ( .A1(n90395), .A2(n110567), .B1(n90396), .B2(n110568), .ZN(
        n91652) );
  AOI22_X1 U77198 ( .A1(n90397), .A2(n73885), .B1(n90398), .B2(n73879), .ZN(
        n91651) );
  NAND2_X1 U77199 ( .A1(n91653), .A2(n91654), .ZN(n91643) );
  AOI22_X1 U77200 ( .A1(n90401), .A2(n110575), .B1(n90402), .B2(n73891), .ZN(
        n91654) );
  AOI22_X1 U77201 ( .A1(n90403), .A2(n110574), .B1(n90404), .B2(n73889), .ZN(
        n91653) );
  NOR4_X1 U77202 ( .A1(n91655), .A2(n91656), .A3(n91657), .A4(n91658), .ZN(
        n91641) );
  NAND2_X1 U77203 ( .A1(n91659), .A2(n91660), .ZN(n91658) );
  AOI22_X1 U77204 ( .A1(n90411), .A2(n110557), .B1(n90412), .B2(n111018), .ZN(
        n91660) );
  AOI22_X1 U77205 ( .A1(n90413), .A2(n110550), .B1(n90414), .B2(n73863), .ZN(
        n91659) );
  NAND2_X1 U77206 ( .A1(n91661), .A2(n91662), .ZN(n91657) );
  AOI22_X1 U77207 ( .A1(n90417), .A2(n110555), .B1(n90418), .B2(n110559), .ZN(
        n91662) );
  AOI22_X1 U77208 ( .A1(n90419), .A2(n110561), .B1(n90420), .B2(n110558), .ZN(
        n91661) );
  NAND2_X1 U77209 ( .A1(n91663), .A2(n91664), .ZN(n91656) );
  AOI22_X1 U77210 ( .A1(n90423), .A2(n73872), .B1(n90424), .B2(n110554), .ZN(
        n91664) );
  AOI22_X1 U77211 ( .A1(n90425), .A2(n110556), .B1(n90426), .B2(n110560), .ZN(
        n91663) );
  NAND2_X1 U77212 ( .A1(n91665), .A2(n91666), .ZN(n91655) );
  AOI22_X1 U77213 ( .A1(n90429), .A2(n110566), .B1(n90430), .B2(n73876), .ZN(
        n91666) );
  AOI22_X1 U77214 ( .A1(n90431), .A2(n73874), .B1(n90432), .B2(n110565), .ZN(
        n91665) );
  NAND2_X1 U77215 ( .A1(n91667), .A2(n91668), .ZN(n91612) );
  NOR4_X1 U77216 ( .A1(n91669), .A2(n91670), .A3(n91671), .A4(n91672), .ZN(
        n91668) );
  NAND2_X1 U77217 ( .A1(n91673), .A2(n91674), .ZN(n91672) );
  AOI22_X1 U77218 ( .A1(n90441), .A2(n73914), .B1(n90442), .B2(n110585), .ZN(
        n91674) );
  AOI22_X1 U77219 ( .A1(n90443), .A2(n110589), .B1(n90444), .B2(n110588), .ZN(
        n91673) );
  NAND2_X1 U77220 ( .A1(n91675), .A2(n91676), .ZN(n91671) );
  AOI22_X1 U77221 ( .A1(n90447), .A2(n110593), .B1(n90448), .B2(n110592), .ZN(
        n91676) );
  AOI22_X1 U77222 ( .A1(n90449), .A2(n110584), .B1(n90450), .B2(n110586), .ZN(
        n91675) );
  NAND2_X1 U77223 ( .A1(n91677), .A2(n91678), .ZN(n91670) );
  AOI22_X1 U77224 ( .A1(n90453), .A2(n110594), .B1(n90454), .B2(n73913), .ZN(
        n91678) );
  AOI22_X1 U77225 ( .A1(n90455), .A2(n73918), .B1(n90456), .B2(n73920), .ZN(
        n91677) );
  NAND2_X1 U77226 ( .A1(n91679), .A2(n91680), .ZN(n91669) );
  AOI22_X1 U77227 ( .A1(n90459), .A2(n110597), .B1(n90460), .B2(n73926), .ZN(
        n91680) );
  AOI22_X1 U77228 ( .A1(n90461), .A2(n110590), .B1(n90462), .B2(n110591), .ZN(
        n91679) );
  NOR4_X1 U77229 ( .A1(n91681), .A2(n91682), .A3(n91683), .A4(n91684), .ZN(
        n91667) );
  NAND2_X1 U77230 ( .A1(n91685), .A2(n91686), .ZN(n91684) );
  AOI22_X1 U77231 ( .A1(n90469), .A2(n110573), .B1(n90470), .B2(n110578), .ZN(
        n91686) );
  AOI22_X1 U77232 ( .A1(n90471), .A2(n110572), .B1(n90472), .B2(n73894), .ZN(
        n91685) );
  NAND2_X1 U77233 ( .A1(n91687), .A2(n91688), .ZN(n91683) );
  AOI22_X1 U77234 ( .A1(n90475), .A2(n73903), .B1(n90476), .B2(n110580), .ZN(
        n91688) );
  AOI22_X1 U77235 ( .A1(n90477), .A2(n110581), .B1(n90478), .B2(n110571), .ZN(
        n91687) );
  NAND2_X1 U77236 ( .A1(n91689), .A2(n91690), .ZN(n91682) );
  AOI22_X1 U77237 ( .A1(n90481), .A2(n110579), .B1(n90482), .B2(n110583), .ZN(
        n91690) );
  AOI22_X1 U77238 ( .A1(n90483), .A2(n110577), .B1(n90484), .B2(n110582), .ZN(
        n91689) );
  NAND2_X1 U77239 ( .A1(n91691), .A2(n91692), .ZN(n91681) );
  AOI22_X1 U77240 ( .A1(n90487), .A2(n73908), .B1(n90488), .B2(n110587), .ZN(
        n91692) );
  AOI22_X1 U77241 ( .A1(n90489), .A2(n73906), .B1(n90490), .B2(n110576), .ZN(
        n91691) );
  NAND2_X1 U77242 ( .A1(n91693), .A2(n91694), .ZN(n91611) );
  NOR4_X1 U77243 ( .A1(n91695), .A2(n91696), .A3(n91697), .A4(n91698), .ZN(
        n91694) );
  NAND2_X1 U77244 ( .A1(n91699), .A2(n91700), .ZN(n91698) );
  AOI22_X1 U77245 ( .A1(n90499), .A2(n110615), .B1(n90500), .B2(n110614), .ZN(
        n91700) );
  AOI22_X1 U77246 ( .A1(n90501), .A2(n73942), .B1(n90502), .B2(n110612), .ZN(
        n91699) );
  NAND2_X1 U77247 ( .A1(n91701), .A2(n91702), .ZN(n91697) );
  AOI22_X1 U77248 ( .A1(n90505), .A2(n110610), .B1(n90506), .B2(n110613), .ZN(
        n91702) );
  AOI22_X1 U77249 ( .A1(n90507), .A2(n110618), .B1(n90508), .B2(n110611), .ZN(
        n91701) );
  NAND2_X1 U77250 ( .A1(n91703), .A2(n91704), .ZN(n91696) );
  AOI22_X1 U77251 ( .A1(n105650), .A2(n110622), .B1(n90512), .B2(n73954), .ZN(
        n91704) );
  AOI22_X1 U77252 ( .A1(n90513), .A2(n110620), .B1(n90514), .B2(n110621), .ZN(
        n91703) );
  NAND2_X1 U77253 ( .A1(n91705), .A2(n91706), .ZN(n91695) );
  AOI22_X1 U77254 ( .A1(n90517), .A2(n110616), .B1(n90518), .B2(n110619), .ZN(
        n91706) );
  AOI22_X1 U77255 ( .A1(n90519), .A2(n73953), .B1(n90520), .B2(n110617), .ZN(
        n91705) );
  NOR4_X1 U77256 ( .A1(n91707), .A2(n91708), .A3(n91709), .A4(n91710), .ZN(
        n91693) );
  NAND2_X1 U77257 ( .A1(n91711), .A2(n91712), .ZN(n91710) );
  AOI22_X1 U77258 ( .A1(n90527), .A2(n110596), .B1(n90528), .B2(n110600), .ZN(
        n91712) );
  AOI22_X1 U77259 ( .A1(n90529), .A2(n110599), .B1(n90530), .B2(n73925), .ZN(
        n91711) );
  NAND2_X1 U77260 ( .A1(n91713), .A2(n91714), .ZN(n91709) );
  AOI22_X1 U77261 ( .A1(n90533), .A2(n110606), .B1(n90534), .B2(n110595), .ZN(
        n91714) );
  AOI22_X1 U77262 ( .A1(n90535), .A2(n110598), .B1(n90536), .B2(n110603), .ZN(
        n91713) );
  NAND2_X1 U77263 ( .A1(n91715), .A2(n91716), .ZN(n91708) );
  AOI22_X1 U77264 ( .A1(n90539), .A2(n110602), .B1(n90540), .B2(n110607), .ZN(
        n91716) );
  AOI22_X1 U77265 ( .A1(n90541), .A2(n110609), .B1(n90542), .B2(n110605), .ZN(
        n91715) );
  NAND2_X1 U77266 ( .A1(n91717), .A2(n91718), .ZN(n91707) );
  AOI22_X1 U77267 ( .A1(n90545), .A2(n73943), .B1(n90546), .B2(n110601), .ZN(
        n91718) );
  AOI22_X1 U77268 ( .A1(n90547), .A2(n110604), .B1(n90548), .B2(n110608), .ZN(
        n91717) );
  AOI21_X1 U77269 ( .B1(n90295), .B2(n87738), .A(n91720), .ZN(n91719) );
  OAI21_X1 U77270 ( .B1(n91721), .B2(n105659), .A(n91722), .ZN(n91720) );
  OAI21_X1 U77271 ( .B1(n91723), .B2(n91724), .A(n105658), .ZN(n91722) );
  OAI21_X1 U77272 ( .B1(n102006), .B2(n90303), .A(n91725), .ZN(n91724) );
  AOI22_X1 U77273 ( .A1(n105656), .A2(n110432), .B1(n90306), .B2(n73696), .ZN(
        n91725) );
  NAND2_X1 U77274 ( .A1(n91726), .A2(n91727), .ZN(n91723) );
  AOI22_X1 U77275 ( .A1(n105654), .A2(n110437), .B1(n105653), .B2(n110434), 
        .ZN(n91727) );
  AOI22_X1 U77276 ( .A1(n90311), .A2(n73694), .B1(n90312), .B2(n110433), .ZN(
        n91726) );
  NOR4_X1 U77277 ( .A1(n91728), .A2(n91729), .A3(n91730), .A4(n91731), .ZN(
        n91721) );
  NAND2_X1 U77278 ( .A1(n91732), .A2(n91733), .ZN(n91731) );
  NOR4_X1 U77279 ( .A1(n91734), .A2(n91735), .A3(n91736), .A4(n91737), .ZN(
        n91733) );
  NAND2_X1 U77280 ( .A1(n91738), .A2(n91739), .ZN(n91737) );
  AOI22_X1 U77281 ( .A1(n90325), .A2(n110413), .B1(n90326), .B2(n110414), .ZN(
        n91739) );
  AOI22_X1 U77282 ( .A1(n90327), .A2(n110422), .B1(n90328), .B2(n110420), .ZN(
        n91738) );
  NAND2_X1 U77283 ( .A1(n91740), .A2(n91741), .ZN(n91736) );
  AOI22_X1 U77284 ( .A1(n90331), .A2(n73563), .B1(n90332), .B2(n110417), .ZN(
        n91741) );
  AOI22_X1 U77285 ( .A1(n90333), .A2(n73667), .B1(n90334), .B2(n110339), .ZN(
        n91740) );
  NAND2_X1 U77286 ( .A1(n91742), .A2(n91743), .ZN(n91735) );
  AOI22_X1 U77287 ( .A1(n90337), .A2(n110342), .B1(n90338), .B2(n73567), .ZN(
        n91743) );
  AOI22_X1 U77288 ( .A1(n90339), .A2(n110418), .B1(n90340), .B2(n110415), .ZN(
        n91742) );
  NAND2_X1 U77289 ( .A1(n91744), .A2(n91745), .ZN(n91734) );
  AOI22_X1 U77290 ( .A1(n90343), .A2(n110340), .B1(n90344), .B2(n110344), .ZN(
        n91745) );
  AOI22_X1 U77291 ( .A1(n90345), .A2(n110343), .B1(n90346), .B2(n73569), .ZN(
        n91744) );
  NOR4_X1 U77292 ( .A1(n91746), .A2(n91747), .A3(n91748), .A4(n91749), .ZN(
        n91732) );
  NAND2_X1 U77293 ( .A1(n91750), .A2(n91751), .ZN(n91749) );
  AOI22_X1 U77294 ( .A1(n90353), .A2(n110423), .B1(n90354), .B2(n110426), .ZN(
        n91751) );
  AOI22_X1 U77295 ( .A1(n90355), .A2(n110427), .B1(n90356), .B2(n110429), .ZN(
        n91750) );
  NAND2_X1 U77296 ( .A1(n91752), .A2(n91753), .ZN(n91748) );
  AOI22_X1 U77297 ( .A1(n90359), .A2(n110428), .B1(n90360), .B2(n110424), .ZN(
        n91753) );
  AOI22_X1 U77298 ( .A1(n90361), .A2(n110430), .B1(n90362), .B2(n110425), .ZN(
        n91752) );
  NAND2_X1 U77299 ( .A1(n91754), .A2(n91755), .ZN(n91747) );
  AOI22_X1 U77300 ( .A1(n90365), .A2(n73677), .B1(n90366), .B2(n73676), .ZN(
        n91755) );
  AOI22_X1 U77301 ( .A1(n90367), .A2(n73679), .B1(n90368), .B2(n110431), .ZN(
        n91754) );
  NAND2_X1 U77302 ( .A1(n91756), .A2(n91757), .ZN(n91746) );
  AOI22_X1 U77303 ( .A1(n90371), .A2(n110416), .B1(n90372), .B2(n110421), .ZN(
        n91757) );
  AOI22_X1 U77304 ( .A1(n90373), .A2(n73674), .B1(n90374), .B2(n110419), .ZN(
        n91756) );
  NAND2_X1 U77305 ( .A1(n91758), .A2(n91759), .ZN(n91730) );
  NOR4_X1 U77306 ( .A1(n91760), .A2(n91761), .A3(n91762), .A4(n91763), .ZN(
        n91759) );
  NAND2_X1 U77307 ( .A1(n91764), .A2(n91765), .ZN(n91763) );
  AOI22_X1 U77308 ( .A1(n90383), .A2(n110353), .B1(n90384), .B2(n110355), .ZN(
        n91765) );
  AOI22_X1 U77309 ( .A1(n90385), .A2(n73592), .B1(n90386), .B2(n110354), .ZN(
        n91764) );
  NAND2_X1 U77310 ( .A1(n91766), .A2(n91767), .ZN(n91762) );
  AOI22_X1 U77311 ( .A1(n90389), .A2(n73596), .B1(n90390), .B2(n73598), .ZN(
        n91767) );
  AOI22_X1 U77312 ( .A1(n90391), .A2(n110360), .B1(n90392), .B2(n110361), .ZN(
        n91766) );
  NAND2_X1 U77313 ( .A1(n91768), .A2(n91769), .ZN(n91761) );
  AOI22_X1 U77314 ( .A1(n90395), .A2(n110358), .B1(n90396), .B2(n110359), .ZN(
        n91769) );
  AOI22_X1 U77315 ( .A1(n90397), .A2(n73597), .B1(n90398), .B2(n73591), .ZN(
        n91768) );
  NAND2_X1 U77316 ( .A1(n91770), .A2(n91771), .ZN(n91760) );
  AOI22_X1 U77317 ( .A1(n90401), .A2(n110366), .B1(n90402), .B2(n73603), .ZN(
        n91771) );
  AOI22_X1 U77318 ( .A1(n90403), .A2(n110365), .B1(n90404), .B2(n73601), .ZN(
        n91770) );
  NOR4_X1 U77319 ( .A1(n91772), .A2(n91773), .A3(n91774), .A4(n91775), .ZN(
        n91758) );
  NAND2_X1 U77320 ( .A1(n91776), .A2(n91777), .ZN(n91775) );
  AOI22_X1 U77321 ( .A1(n90411), .A2(n110348), .B1(n90412), .B2(n111019), .ZN(
        n91777) );
  AOI22_X1 U77322 ( .A1(n90413), .A2(n110341), .B1(n90414), .B2(n73575), .ZN(
        n91776) );
  NAND2_X1 U77323 ( .A1(n91778), .A2(n91779), .ZN(n91774) );
  AOI22_X1 U77324 ( .A1(n90417), .A2(n110346), .B1(n90418), .B2(n110350), .ZN(
        n91779) );
  AOI22_X1 U77325 ( .A1(n90419), .A2(n110352), .B1(n90420), .B2(n110349), .ZN(
        n91778) );
  NAND2_X1 U77326 ( .A1(n91780), .A2(n91781), .ZN(n91773) );
  AOI22_X1 U77327 ( .A1(n90423), .A2(n73584), .B1(n90424), .B2(n110345), .ZN(
        n91781) );
  AOI22_X1 U77328 ( .A1(n90425), .A2(n110347), .B1(n90426), .B2(n110351), .ZN(
        n91780) );
  NAND2_X1 U77329 ( .A1(n91782), .A2(n91783), .ZN(n91772) );
  AOI22_X1 U77330 ( .A1(n90429), .A2(n110357), .B1(n90430), .B2(n73588), .ZN(
        n91783) );
  AOI22_X1 U77331 ( .A1(n90431), .A2(n73586), .B1(n90432), .B2(n110356), .ZN(
        n91782) );
  NAND2_X1 U77332 ( .A1(n91784), .A2(n91785), .ZN(n91729) );
  NOR4_X1 U77333 ( .A1(n91786), .A2(n91787), .A3(n91788), .A4(n91789), .ZN(
        n91785) );
  NAND2_X1 U77334 ( .A1(n91790), .A2(n91791), .ZN(n91789) );
  AOI22_X1 U77335 ( .A1(n90441), .A2(n73626), .B1(n90442), .B2(n110376), .ZN(
        n91791) );
  AOI22_X1 U77336 ( .A1(n90443), .A2(n110380), .B1(n90444), .B2(n110379), .ZN(
        n91790) );
  NAND2_X1 U77337 ( .A1(n91792), .A2(n91793), .ZN(n91788) );
  AOI22_X1 U77338 ( .A1(n90447), .A2(n110383), .B1(n90448), .B2(n110382), .ZN(
        n91793) );
  AOI22_X1 U77339 ( .A1(n90449), .A2(n110375), .B1(n90450), .B2(n110377), .ZN(
        n91792) );
  NAND2_X1 U77340 ( .A1(n91794), .A2(n91795), .ZN(n91787) );
  AOI22_X1 U77341 ( .A1(n90453), .A2(n110384), .B1(n90454), .B2(n73625), .ZN(
        n91795) );
  AOI22_X1 U77342 ( .A1(n90455), .A2(n73630), .B1(n90456), .B2(n73632), .ZN(
        n91794) );
  NAND2_X1 U77343 ( .A1(n91796), .A2(n91797), .ZN(n91786) );
  AOI22_X1 U77344 ( .A1(n90459), .A2(n110387), .B1(n90460), .B2(n73638), .ZN(
        n91797) );
  AOI22_X1 U77345 ( .A1(n90461), .A2(n110381), .B1(n90462), .B2(n73627), .ZN(
        n91796) );
  NOR4_X1 U77346 ( .A1(n91798), .A2(n91799), .A3(n91800), .A4(n91801), .ZN(
        n91784) );
  NAND2_X1 U77347 ( .A1(n91802), .A2(n91803), .ZN(n91801) );
  AOI22_X1 U77348 ( .A1(n90469), .A2(n110364), .B1(n90470), .B2(n110369), .ZN(
        n91803) );
  AOI22_X1 U77349 ( .A1(n90471), .A2(n110363), .B1(n90472), .B2(n73606), .ZN(
        n91802) );
  NAND2_X1 U77350 ( .A1(n91804), .A2(n91805), .ZN(n91800) );
  AOI22_X1 U77351 ( .A1(n90475), .A2(n73615), .B1(n90476), .B2(n110371), .ZN(
        n91805) );
  AOI22_X1 U77352 ( .A1(n90477), .A2(n110372), .B1(n90478), .B2(n110362), .ZN(
        n91804) );
  NAND2_X1 U77353 ( .A1(n91806), .A2(n91807), .ZN(n91799) );
  AOI22_X1 U77354 ( .A1(n90481), .A2(n110370), .B1(n90482), .B2(n110374), .ZN(
        n91807) );
  AOI22_X1 U77355 ( .A1(n90483), .A2(n110368), .B1(n90484), .B2(n110373), .ZN(
        n91806) );
  NAND2_X1 U77356 ( .A1(n91808), .A2(n91809), .ZN(n91798) );
  AOI22_X1 U77357 ( .A1(n90487), .A2(n73620), .B1(n90488), .B2(n110378), .ZN(
        n91809) );
  AOI22_X1 U77358 ( .A1(n90489), .A2(n73618), .B1(n90490), .B2(n110367), .ZN(
        n91808) );
  NAND2_X1 U77359 ( .A1(n91810), .A2(n91811), .ZN(n91728) );
  NOR4_X1 U77360 ( .A1(n91812), .A2(n91813), .A3(n91814), .A4(n91815), .ZN(
        n91811) );
  NAND2_X1 U77361 ( .A1(n91816), .A2(n91817), .ZN(n91815) );
  AOI22_X1 U77362 ( .A1(n90499), .A2(n110404), .B1(n90500), .B2(n110403), .ZN(
        n91817) );
  AOI22_X1 U77363 ( .A1(n90501), .A2(n73654), .B1(n90502), .B2(n110401), .ZN(
        n91816) );
  NAND2_X1 U77364 ( .A1(n91818), .A2(n91819), .ZN(n91814) );
  AOI22_X1 U77365 ( .A1(n90505), .A2(n110399), .B1(n90506), .B2(n110402), .ZN(
        n91819) );
  AOI22_X1 U77366 ( .A1(n105651), .A2(n73660), .B1(n90508), .B2(n110400), .ZN(
        n91818) );
  NAND2_X1 U77367 ( .A1(n91820), .A2(n91821), .ZN(n91813) );
  AOI22_X1 U77368 ( .A1(n105650), .A2(n110410), .B1(n90512), .B2(n73666), .ZN(
        n91821) );
  AOI22_X1 U77369 ( .A1(n105648), .A2(n110408), .B1(n90514), .B2(n110409), 
        .ZN(n91820) );
  NAND2_X1 U77370 ( .A1(n91822), .A2(n91823), .ZN(n91812) );
  AOI22_X1 U77371 ( .A1(n90517), .A2(n110405), .B1(n90518), .B2(n110407), .ZN(
        n91823) );
  AOI22_X1 U77372 ( .A1(n105645), .A2(n110411), .B1(n90520), .B2(n110406), 
        .ZN(n91822) );
  NOR4_X1 U77373 ( .A1(n91824), .A2(n91825), .A3(n91826), .A4(n91827), .ZN(
        n91810) );
  NAND2_X1 U77374 ( .A1(n91828), .A2(n91829), .ZN(n91827) );
  AOI22_X1 U77375 ( .A1(n90527), .A2(n110386), .B1(n90528), .B2(n110389), .ZN(
        n91829) );
  AOI22_X1 U77376 ( .A1(n90529), .A2(n111038), .B1(n90530), .B2(n73637), .ZN(
        n91828) );
  NAND2_X1 U77377 ( .A1(n91830), .A2(n91831), .ZN(n91826) );
  AOI22_X1 U77378 ( .A1(n90533), .A2(n110395), .B1(n90534), .B2(n110385), .ZN(
        n91831) );
  AOI22_X1 U77379 ( .A1(n90535), .A2(n110388), .B1(n90536), .B2(n110392), .ZN(
        n91830) );
  NAND2_X1 U77380 ( .A1(n91832), .A2(n91833), .ZN(n91825) );
  AOI22_X1 U77381 ( .A1(n90539), .A2(n110391), .B1(n90540), .B2(n110396), .ZN(
        n91833) );
  AOI22_X1 U77382 ( .A1(n90541), .A2(n110398), .B1(n90542), .B2(n110394), .ZN(
        n91832) );
  NAND2_X1 U77383 ( .A1(n91834), .A2(n91835), .ZN(n91824) );
  AOI22_X1 U77384 ( .A1(n90545), .A2(n73655), .B1(n90546), .B2(n110390), .ZN(
        n91835) );
  AOI22_X1 U77385 ( .A1(n90547), .A2(n110393), .B1(n90548), .B2(n110397), .ZN(
        n91834) );
  AOI21_X1 U77386 ( .B1(n90295), .B2(n87856), .A(n91837), .ZN(n91836) );
  OAI21_X1 U77387 ( .B1(n91838), .B2(n105659), .A(n91839), .ZN(n91837) );
  OAI21_X1 U77388 ( .B1(n91840), .B2(n91841), .A(n105658), .ZN(n91839) );
  OAI21_X1 U77389 ( .B1(n101988), .B2(n105657), .A(n91842), .ZN(n91841) );
  AOI22_X1 U77390 ( .A1(n105656), .A2(n110110), .B1(n105655), .B2(n73258), 
        .ZN(n91842) );
  NAND2_X1 U77391 ( .A1(n91843), .A2(n91844), .ZN(n91840) );
  AOI22_X1 U77392 ( .A1(n105654), .A2(n110115), .B1(n105653), .B2(n110112), 
        .ZN(n91844) );
  AOI22_X1 U77393 ( .A1(n90311), .A2(n73256), .B1(n105652), .B2(n110111), .ZN(
        n91843) );
  NOR4_X1 U77394 ( .A1(n91845), .A2(n91846), .A3(n91847), .A4(n91848), .ZN(
        n91838) );
  NAND2_X1 U77395 ( .A1(n91849), .A2(n91850), .ZN(n91848) );
  NOR4_X1 U77396 ( .A1(n91851), .A2(n91852), .A3(n91853), .A4(n91854), .ZN(
        n91850) );
  NAND2_X1 U77397 ( .A1(n91855), .A2(n91856), .ZN(n91854) );
  AOI22_X1 U77398 ( .A1(n90325), .A2(n110091), .B1(n90326), .B2(n110092), .ZN(
        n91856) );
  AOI22_X1 U77399 ( .A1(n90327), .A2(n110100), .B1(n90328), .B2(n110098), .ZN(
        n91855) );
  NAND2_X1 U77400 ( .A1(n91857), .A2(n91858), .ZN(n91853) );
  AOI22_X1 U77401 ( .A1(n90331), .A2(n73125), .B1(n90332), .B2(n110095), .ZN(
        n91858) );
  AOI22_X1 U77402 ( .A1(n90333), .A2(n73229), .B1(n90334), .B2(n110013), .ZN(
        n91857) );
  NAND2_X1 U77403 ( .A1(n91859), .A2(n91860), .ZN(n91852) );
  AOI22_X1 U77404 ( .A1(n90337), .A2(n110017), .B1(n90338), .B2(n73129), .ZN(
        n91860) );
  AOI22_X1 U77405 ( .A1(n90339), .A2(n110096), .B1(n90340), .B2(n110093), .ZN(
        n91859) );
  NAND2_X1 U77406 ( .A1(n91861), .A2(n91862), .ZN(n91851) );
  AOI22_X1 U77407 ( .A1(n90343), .A2(n110015), .B1(n90344), .B2(n110019), .ZN(
        n91862) );
  AOI22_X1 U77408 ( .A1(n90345), .A2(n110018), .B1(n90346), .B2(n73131), .ZN(
        n91861) );
  NOR4_X1 U77409 ( .A1(n91863), .A2(n91864), .A3(n91865), .A4(n91866), .ZN(
        n91849) );
  NAND2_X1 U77410 ( .A1(n91867), .A2(n91868), .ZN(n91866) );
  AOI22_X1 U77411 ( .A1(n90353), .A2(n110101), .B1(n90354), .B2(n110104), .ZN(
        n91868) );
  AOI22_X1 U77412 ( .A1(n90355), .A2(n110105), .B1(n90356), .B2(n110107), .ZN(
        n91867) );
  NAND2_X1 U77413 ( .A1(n91869), .A2(n91870), .ZN(n91865) );
  AOI22_X1 U77414 ( .A1(n90359), .A2(n110106), .B1(n90360), .B2(n110102), .ZN(
        n91870) );
  AOI22_X1 U77415 ( .A1(n90361), .A2(n110108), .B1(n90362), .B2(n110103), .ZN(
        n91869) );
  NAND2_X1 U77416 ( .A1(n91871), .A2(n91872), .ZN(n91864) );
  AOI22_X1 U77417 ( .A1(n90365), .A2(n73239), .B1(n90366), .B2(n73238), .ZN(
        n91872) );
  AOI22_X1 U77418 ( .A1(n90367), .A2(n73241), .B1(n90368), .B2(n110109), .ZN(
        n91871) );
  NAND2_X1 U77419 ( .A1(n91873), .A2(n91874), .ZN(n91863) );
  AOI22_X1 U77420 ( .A1(n90371), .A2(n110094), .B1(n90372), .B2(n110099), .ZN(
        n91874) );
  AOI22_X1 U77421 ( .A1(n90373), .A2(n73236), .B1(n90374), .B2(n110097), .ZN(
        n91873) );
  NAND2_X1 U77422 ( .A1(n91875), .A2(n91876), .ZN(n91847) );
  NOR4_X1 U77423 ( .A1(n91877), .A2(n91878), .A3(n91879), .A4(n91880), .ZN(
        n91876) );
  NAND2_X1 U77424 ( .A1(n91881), .A2(n91882), .ZN(n91880) );
  AOI22_X1 U77425 ( .A1(n90383), .A2(n110028), .B1(n90384), .B2(n110030), .ZN(
        n91882) );
  AOI22_X1 U77426 ( .A1(n90385), .A2(n73154), .B1(n90386), .B2(n110029), .ZN(
        n91881) );
  NAND2_X1 U77427 ( .A1(n91883), .A2(n91884), .ZN(n91879) );
  AOI22_X1 U77428 ( .A1(n90389), .A2(n73158), .B1(n90390), .B2(n73160), .ZN(
        n91884) );
  AOI22_X1 U77429 ( .A1(n90391), .A2(n110036), .B1(n90392), .B2(n110037), .ZN(
        n91883) );
  NAND2_X1 U77430 ( .A1(n91885), .A2(n91886), .ZN(n91878) );
  AOI22_X1 U77431 ( .A1(n90395), .A2(n110033), .B1(n90396), .B2(n110035), .ZN(
        n91886) );
  AOI22_X1 U77432 ( .A1(n90397), .A2(n73159), .B1(n90398), .B2(n110034), .ZN(
        n91885) );
  NAND2_X1 U77433 ( .A1(n91887), .A2(n91888), .ZN(n91877) );
  AOI22_X1 U77434 ( .A1(n90401), .A2(n110042), .B1(n90402), .B2(n73165), .ZN(
        n91888) );
  AOI22_X1 U77435 ( .A1(n90403), .A2(n110041), .B1(n90404), .B2(n73163), .ZN(
        n91887) );
  NOR4_X1 U77436 ( .A1(n91889), .A2(n91890), .A3(n91891), .A4(n91892), .ZN(
        n91875) );
  NAND2_X1 U77437 ( .A1(n91893), .A2(n91894), .ZN(n91892) );
  AOI22_X1 U77438 ( .A1(n90411), .A2(n110023), .B1(n90412), .B2(n110014), .ZN(
        n91894) );
  AOI22_X1 U77439 ( .A1(n90413), .A2(n110016), .B1(n90414), .B2(n73137), .ZN(
        n91893) );
  NAND2_X1 U77440 ( .A1(n91895), .A2(n91896), .ZN(n91891) );
  AOI22_X1 U77441 ( .A1(n90417), .A2(n110021), .B1(n90418), .B2(n110025), .ZN(
        n91896) );
  AOI22_X1 U77442 ( .A1(n90419), .A2(n110027), .B1(n90420), .B2(n110024), .ZN(
        n91895) );
  NAND2_X1 U77443 ( .A1(n91897), .A2(n91898), .ZN(n91890) );
  AOI22_X1 U77444 ( .A1(n90423), .A2(n73146), .B1(n90424), .B2(n110020), .ZN(
        n91898) );
  AOI22_X1 U77445 ( .A1(n90425), .A2(n110022), .B1(n90426), .B2(n110026), .ZN(
        n91897) );
  NAND2_X1 U77446 ( .A1(n91899), .A2(n91900), .ZN(n91889) );
  AOI22_X1 U77447 ( .A1(n90429), .A2(n110032), .B1(n90430), .B2(n73150), .ZN(
        n91900) );
  AOI22_X1 U77448 ( .A1(n90431), .A2(n73148), .B1(n90432), .B2(n110031), .ZN(
        n91899) );
  NAND2_X1 U77449 ( .A1(n91901), .A2(n91902), .ZN(n91846) );
  NOR4_X1 U77450 ( .A1(n91903), .A2(n91904), .A3(n91905), .A4(n91906), .ZN(
        n91902) );
  NAND2_X1 U77451 ( .A1(n91907), .A2(n91908), .ZN(n91906) );
  AOI22_X1 U77452 ( .A1(n90441), .A2(n73188), .B1(n90442), .B2(n110052), .ZN(
        n91908) );
  AOI22_X1 U77453 ( .A1(n90443), .A2(n110056), .B1(n90444), .B2(n110055), .ZN(
        n91907) );
  NAND2_X1 U77454 ( .A1(n91909), .A2(n91910), .ZN(n91905) );
  AOI22_X1 U77455 ( .A1(n90447), .A2(n110061), .B1(n90448), .B2(n110060), .ZN(
        n91910) );
  AOI22_X1 U77456 ( .A1(n90449), .A2(n110051), .B1(n90450), .B2(n110053), .ZN(
        n91909) );
  NAND2_X1 U77457 ( .A1(n91911), .A2(n91912), .ZN(n91904) );
  AOI22_X1 U77458 ( .A1(n90453), .A2(n110062), .B1(n90454), .B2(n110058), .ZN(
        n91912) );
  AOI22_X1 U77459 ( .A1(n90455), .A2(n73192), .B1(n90456), .B2(n73194), .ZN(
        n91911) );
  NAND2_X1 U77460 ( .A1(n91913), .A2(n91914), .ZN(n91903) );
  AOI22_X1 U77461 ( .A1(n90459), .A2(n110065), .B1(n90460), .B2(n73200), .ZN(
        n91914) );
  AOI22_X1 U77462 ( .A1(n90461), .A2(n110057), .B1(n90462), .B2(n110059), .ZN(
        n91913) );
  NOR4_X1 U77463 ( .A1(n91915), .A2(n91916), .A3(n91917), .A4(n91918), .ZN(
        n91901) );
  NAND2_X1 U77464 ( .A1(n91919), .A2(n91920), .ZN(n91918) );
  AOI22_X1 U77465 ( .A1(n90469), .A2(n110040), .B1(n90470), .B2(n110045), .ZN(
        n91920) );
  AOI22_X1 U77466 ( .A1(n90471), .A2(n110039), .B1(n90472), .B2(n73168), .ZN(
        n91919) );
  NAND2_X1 U77467 ( .A1(n91921), .A2(n91922), .ZN(n91917) );
  AOI22_X1 U77468 ( .A1(n90475), .A2(n73177), .B1(n90476), .B2(n110047), .ZN(
        n91922) );
  AOI22_X1 U77469 ( .A1(n90477), .A2(n110048), .B1(n90478), .B2(n110038), .ZN(
        n91921) );
  NAND2_X1 U77470 ( .A1(n91923), .A2(n91924), .ZN(n91916) );
  AOI22_X1 U77471 ( .A1(n90481), .A2(n110046), .B1(n90482), .B2(n110050), .ZN(
        n91924) );
  AOI22_X1 U77472 ( .A1(n90483), .A2(n110044), .B1(n90484), .B2(n110049), .ZN(
        n91923) );
  NAND2_X1 U77473 ( .A1(n91925), .A2(n91926), .ZN(n91915) );
  AOI22_X1 U77474 ( .A1(n90487), .A2(n73182), .B1(n90488), .B2(n110054), .ZN(
        n91926) );
  AOI22_X1 U77475 ( .A1(n90489), .A2(n73180), .B1(n90490), .B2(n110043), .ZN(
        n91925) );
  NAND2_X1 U77476 ( .A1(n91927), .A2(n91928), .ZN(n91845) );
  NOR4_X1 U77477 ( .A1(n91929), .A2(n91930), .A3(n91931), .A4(n91932), .ZN(
        n91928) );
  NAND2_X1 U77478 ( .A1(n91933), .A2(n91934), .ZN(n91932) );
  AOI22_X1 U77479 ( .A1(n90499), .A2(n110082), .B1(n90500), .B2(n110081), .ZN(
        n91934) );
  AOI22_X1 U77480 ( .A1(n90501), .A2(n73216), .B1(n90502), .B2(n110079), .ZN(
        n91933) );
  NAND2_X1 U77481 ( .A1(n91935), .A2(n91936), .ZN(n91931) );
  AOI22_X1 U77482 ( .A1(n90505), .A2(n110077), .B1(n90506), .B2(n110080), .ZN(
        n91936) );
  AOI22_X1 U77483 ( .A1(n105651), .A2(n73222), .B1(n90508), .B2(n110078), .ZN(
        n91935) );
  NAND2_X1 U77484 ( .A1(n91937), .A2(n91938), .ZN(n91930) );
  AOI22_X1 U77485 ( .A1(n105650), .A2(n110088), .B1(n105649), .B2(n73228), 
        .ZN(n91938) );
  AOI22_X1 U77486 ( .A1(n105648), .A2(n110086), .B1(n105647), .B2(n110087), 
        .ZN(n91937) );
  NAND2_X1 U77487 ( .A1(n91939), .A2(n91940), .ZN(n91929) );
  AOI22_X1 U77488 ( .A1(n90517), .A2(n110083), .B1(n105646), .B2(n110085), 
        .ZN(n91940) );
  AOI22_X1 U77489 ( .A1(n105645), .A2(n110089), .B1(n90520), .B2(n110084), 
        .ZN(n91939) );
  NOR4_X1 U77490 ( .A1(n91941), .A2(n91942), .A3(n91943), .A4(n91944), .ZN(
        n91927) );
  NAND2_X1 U77491 ( .A1(n91945), .A2(n91946), .ZN(n91944) );
  AOI22_X1 U77492 ( .A1(n90527), .A2(n110064), .B1(n90528), .B2(n110067), .ZN(
        n91946) );
  AOI22_X1 U77493 ( .A1(n90529), .A2(n111040), .B1(n90530), .B2(n73199), .ZN(
        n91945) );
  NAND2_X1 U77494 ( .A1(n91947), .A2(n91948), .ZN(n91943) );
  AOI22_X1 U77495 ( .A1(n90533), .A2(n110073), .B1(n90534), .B2(n110063), .ZN(
        n91948) );
  AOI22_X1 U77496 ( .A1(n90535), .A2(n110066), .B1(n90536), .B2(n110070), .ZN(
        n91947) );
  NAND2_X1 U77497 ( .A1(n91949), .A2(n91950), .ZN(n91942) );
  AOI22_X1 U77498 ( .A1(n90539), .A2(n110069), .B1(n90540), .B2(n110074), .ZN(
        n91950) );
  AOI22_X1 U77499 ( .A1(n90541), .A2(n110076), .B1(n90542), .B2(n110072), .ZN(
        n91949) );
  NAND2_X1 U77500 ( .A1(n91951), .A2(n91952), .ZN(n91941) );
  AOI22_X1 U77501 ( .A1(n90545), .A2(n73217), .B1(n90546), .B2(n110068), .ZN(
        n91952) );
  AOI22_X1 U77502 ( .A1(n90547), .A2(n110071), .B1(n90548), .B2(n110075), .ZN(
        n91951) );
  AOI21_X1 U77503 ( .B1(n90295), .B2(n87974), .A(n91954), .ZN(n91953) );
  OAI21_X1 U77504 ( .B1(n91955), .B2(n105659), .A(n91956), .ZN(n91954) );
  OAI21_X1 U77505 ( .B1(n91957), .B2(n91958), .A(n105658), .ZN(n91956) );
  OAI21_X1 U77506 ( .B1(n101972), .B2(n90303), .A(n91959), .ZN(n91958) );
  AOI22_X1 U77507 ( .A1(n105656), .A2(n110217), .B1(n105655), .B2(n73400), 
        .ZN(n91959) );
  NAND2_X1 U77508 ( .A1(n91960), .A2(n91961), .ZN(n91957) );
  AOI22_X1 U77509 ( .A1(n105654), .A2(n110222), .B1(n105653), .B2(n110219), 
        .ZN(n91961) );
  AOI22_X1 U77510 ( .A1(n90311), .A2(n73398), .B1(n105652), .B2(n110218), .ZN(
        n91960) );
  NOR4_X1 U77511 ( .A1(n91962), .A2(n91963), .A3(n91964), .A4(n91965), .ZN(
        n91955) );
  NAND2_X1 U77512 ( .A1(n91966), .A2(n91967), .ZN(n91965) );
  NOR4_X1 U77513 ( .A1(n91968), .A2(n91969), .A3(n91970), .A4(n91971), .ZN(
        n91967) );
  NAND2_X1 U77514 ( .A1(n91972), .A2(n91973), .ZN(n91971) );
  AOI22_X1 U77515 ( .A1(n90325), .A2(n110198), .B1(n90326), .B2(n110199), .ZN(
        n91973) );
  AOI22_X1 U77516 ( .A1(n90327), .A2(n110207), .B1(n90328), .B2(n110205), .ZN(
        n91972) );
  NAND2_X1 U77517 ( .A1(n91974), .A2(n91975), .ZN(n91970) );
  AOI22_X1 U77518 ( .A1(n90331), .A2(n73267), .B1(n90332), .B2(n110202), .ZN(
        n91975) );
  AOI22_X1 U77519 ( .A1(n90333), .A2(n73371), .B1(n90334), .B2(n110121), .ZN(
        n91974) );
  NAND2_X1 U77520 ( .A1(n91976), .A2(n91977), .ZN(n91969) );
  AOI22_X1 U77521 ( .A1(n90337), .A2(n110124), .B1(n90338), .B2(n73271), .ZN(
        n91977) );
  AOI22_X1 U77522 ( .A1(n90339), .A2(n110203), .B1(n90340), .B2(n110200), .ZN(
        n91976) );
  NAND2_X1 U77523 ( .A1(n91978), .A2(n91979), .ZN(n91968) );
  AOI22_X1 U77524 ( .A1(n90343), .A2(n110122), .B1(n90344), .B2(n110126), .ZN(
        n91979) );
  AOI22_X1 U77525 ( .A1(n90345), .A2(n110125), .B1(n90346), .B2(n73273), .ZN(
        n91978) );
  NOR4_X1 U77526 ( .A1(n91980), .A2(n91981), .A3(n91982), .A4(n91983), .ZN(
        n91966) );
  NAND2_X1 U77527 ( .A1(n91984), .A2(n91985), .ZN(n91983) );
  AOI22_X1 U77528 ( .A1(n90353), .A2(n110208), .B1(n90354), .B2(n110211), .ZN(
        n91985) );
  AOI22_X1 U77529 ( .A1(n90355), .A2(n110212), .B1(n90356), .B2(n110214), .ZN(
        n91984) );
  NAND2_X1 U77530 ( .A1(n91986), .A2(n91987), .ZN(n91982) );
  AOI22_X1 U77531 ( .A1(n90359), .A2(n110213), .B1(n90360), .B2(n110209), .ZN(
        n91987) );
  AOI22_X1 U77532 ( .A1(n90361), .A2(n110215), .B1(n90362), .B2(n110210), .ZN(
        n91986) );
  NAND2_X1 U77533 ( .A1(n91988), .A2(n91989), .ZN(n91981) );
  AOI22_X1 U77534 ( .A1(n90365), .A2(n73381), .B1(n90366), .B2(n73380), .ZN(
        n91989) );
  AOI22_X1 U77535 ( .A1(n90367), .A2(n73383), .B1(n90368), .B2(n110216), .ZN(
        n91988) );
  NAND2_X1 U77536 ( .A1(n91990), .A2(n91991), .ZN(n91980) );
  AOI22_X1 U77537 ( .A1(n90371), .A2(n110201), .B1(n90372), .B2(n110206), .ZN(
        n91991) );
  AOI22_X1 U77538 ( .A1(n90373), .A2(n73378), .B1(n90374), .B2(n110204), .ZN(
        n91990) );
  NAND2_X1 U77539 ( .A1(n91992), .A2(n91993), .ZN(n91964) );
  NOR4_X1 U77540 ( .A1(n91994), .A2(n91995), .A3(n91996), .A4(n91997), .ZN(
        n91993) );
  NAND2_X1 U77541 ( .A1(n91998), .A2(n91999), .ZN(n91997) );
  AOI22_X1 U77542 ( .A1(n90383), .A2(n110135), .B1(n90384), .B2(n110137), .ZN(
        n91999) );
  AOI22_X1 U77543 ( .A1(n90385), .A2(n73296), .B1(n90386), .B2(n110136), .ZN(
        n91998) );
  NAND2_X1 U77544 ( .A1(n92000), .A2(n92001), .ZN(n91996) );
  AOI22_X1 U77545 ( .A1(n90389), .A2(n73300), .B1(n90390), .B2(n73302), .ZN(
        n92001) );
  AOI22_X1 U77546 ( .A1(n90391), .A2(n110143), .B1(n90392), .B2(n110144), .ZN(
        n92000) );
  NAND2_X1 U77547 ( .A1(n92002), .A2(n92003), .ZN(n91995) );
  AOI22_X1 U77548 ( .A1(n90395), .A2(n110140), .B1(n90396), .B2(n110142), .ZN(
        n92003) );
  AOI22_X1 U77549 ( .A1(n90397), .A2(n73301), .B1(n90398), .B2(n110141), .ZN(
        n92002) );
  NAND2_X1 U77550 ( .A1(n92004), .A2(n92005), .ZN(n91994) );
  AOI22_X1 U77551 ( .A1(n90401), .A2(n110149), .B1(n90402), .B2(n73307), .ZN(
        n92005) );
  AOI22_X1 U77552 ( .A1(n90403), .A2(n110148), .B1(n90404), .B2(n73305), .ZN(
        n92004) );
  NOR4_X1 U77553 ( .A1(n92006), .A2(n92007), .A3(n92008), .A4(n92009), .ZN(
        n91992) );
  NAND2_X1 U77554 ( .A1(n92010), .A2(n92011), .ZN(n92009) );
  AOI22_X1 U77555 ( .A1(n90411), .A2(n110130), .B1(n90412), .B2(n111021), .ZN(
        n92011) );
  AOI22_X1 U77556 ( .A1(n90413), .A2(n110123), .B1(n90414), .B2(n73279), .ZN(
        n92010) );
  NAND2_X1 U77557 ( .A1(n92012), .A2(n92013), .ZN(n92008) );
  AOI22_X1 U77558 ( .A1(n90417), .A2(n110128), .B1(n90418), .B2(n110132), .ZN(
        n92013) );
  AOI22_X1 U77559 ( .A1(n90419), .A2(n110134), .B1(n90420), .B2(n110131), .ZN(
        n92012) );
  NAND2_X1 U77560 ( .A1(n92014), .A2(n92015), .ZN(n92007) );
  AOI22_X1 U77561 ( .A1(n90423), .A2(n73288), .B1(n90424), .B2(n110127), .ZN(
        n92015) );
  AOI22_X1 U77562 ( .A1(n90425), .A2(n110129), .B1(n90426), .B2(n110133), .ZN(
        n92014) );
  NAND2_X1 U77563 ( .A1(n92016), .A2(n92017), .ZN(n92006) );
  AOI22_X1 U77564 ( .A1(n90429), .A2(n110139), .B1(n90430), .B2(n73292), .ZN(
        n92017) );
  AOI22_X1 U77565 ( .A1(n90431), .A2(n73290), .B1(n90432), .B2(n110138), .ZN(
        n92016) );
  NAND2_X1 U77566 ( .A1(n92018), .A2(n92019), .ZN(n91963) );
  NOR4_X1 U77567 ( .A1(n92020), .A2(n92021), .A3(n92022), .A4(n92023), .ZN(
        n92019) );
  NAND2_X1 U77568 ( .A1(n92024), .A2(n92025), .ZN(n92023) );
  AOI22_X1 U77569 ( .A1(n90441), .A2(n73330), .B1(n90442), .B2(n110159), .ZN(
        n92025) );
  AOI22_X1 U77570 ( .A1(n90443), .A2(n110163), .B1(n90444), .B2(n110162), .ZN(
        n92024) );
  NAND2_X1 U77571 ( .A1(n92026), .A2(n92027), .ZN(n92022) );
  AOI22_X1 U77572 ( .A1(n90447), .A2(n110168), .B1(n90448), .B2(n110167), .ZN(
        n92027) );
  AOI22_X1 U77573 ( .A1(n90449), .A2(n110158), .B1(n90450), .B2(n110160), .ZN(
        n92026) );
  NAND2_X1 U77574 ( .A1(n92028), .A2(n92029), .ZN(n92021) );
  AOI22_X1 U77575 ( .A1(n90453), .A2(n110169), .B1(n90454), .B2(n110165), .ZN(
        n92029) );
  AOI22_X1 U77576 ( .A1(n90455), .A2(n73334), .B1(n90456), .B2(n73336), .ZN(
        n92028) );
  NAND2_X1 U77577 ( .A1(n92030), .A2(n92031), .ZN(n92020) );
  AOI22_X1 U77578 ( .A1(n90459), .A2(n110172), .B1(n90460), .B2(n73342), .ZN(
        n92031) );
  AOI22_X1 U77579 ( .A1(n90461), .A2(n110164), .B1(n90462), .B2(n110166), .ZN(
        n92030) );
  NOR4_X1 U77580 ( .A1(n92032), .A2(n92033), .A3(n92034), .A4(n92035), .ZN(
        n92018) );
  NAND2_X1 U77581 ( .A1(n92036), .A2(n92037), .ZN(n92035) );
  AOI22_X1 U77582 ( .A1(n90469), .A2(n110147), .B1(n90470), .B2(n110152), .ZN(
        n92037) );
  AOI22_X1 U77583 ( .A1(n90471), .A2(n110146), .B1(n90472), .B2(n73310), .ZN(
        n92036) );
  NAND2_X1 U77584 ( .A1(n92038), .A2(n92039), .ZN(n92034) );
  AOI22_X1 U77585 ( .A1(n90475), .A2(n73319), .B1(n90476), .B2(n110154), .ZN(
        n92039) );
  AOI22_X1 U77586 ( .A1(n90477), .A2(n110155), .B1(n90478), .B2(n110145), .ZN(
        n92038) );
  NAND2_X1 U77587 ( .A1(n92040), .A2(n92041), .ZN(n92033) );
  AOI22_X1 U77588 ( .A1(n90481), .A2(n110153), .B1(n90482), .B2(n110157), .ZN(
        n92041) );
  AOI22_X1 U77589 ( .A1(n90483), .A2(n110151), .B1(n90484), .B2(n110156), .ZN(
        n92040) );
  NAND2_X1 U77590 ( .A1(n92042), .A2(n92043), .ZN(n92032) );
  AOI22_X1 U77591 ( .A1(n90487), .A2(n73324), .B1(n90488), .B2(n110161), .ZN(
        n92043) );
  AOI22_X1 U77592 ( .A1(n90489), .A2(n73322), .B1(n90490), .B2(n110150), .ZN(
        n92042) );
  NAND2_X1 U77593 ( .A1(n92044), .A2(n92045), .ZN(n91962) );
  NOR4_X1 U77594 ( .A1(n92046), .A2(n92047), .A3(n92048), .A4(n92049), .ZN(
        n92045) );
  NAND2_X1 U77595 ( .A1(n92050), .A2(n92051), .ZN(n92049) );
  AOI22_X1 U77596 ( .A1(n90499), .A2(n110189), .B1(n90500), .B2(n110188), .ZN(
        n92051) );
  AOI22_X1 U77597 ( .A1(n90501), .A2(n73358), .B1(n90502), .B2(n110186), .ZN(
        n92050) );
  NAND2_X1 U77598 ( .A1(n92052), .A2(n92053), .ZN(n92048) );
  AOI22_X1 U77599 ( .A1(n90505), .A2(n110184), .B1(n90506), .B2(n110187), .ZN(
        n92053) );
  AOI22_X1 U77600 ( .A1(n105651), .A2(n73364), .B1(n90508), .B2(n110185), .ZN(
        n92052) );
  NAND2_X1 U77601 ( .A1(n92054), .A2(n92055), .ZN(n92047) );
  AOI22_X1 U77602 ( .A1(n105650), .A2(n110195), .B1(n105649), .B2(n73370), 
        .ZN(n92055) );
  AOI22_X1 U77603 ( .A1(n105648), .A2(n110193), .B1(n105647), .B2(n110194), 
        .ZN(n92054) );
  NAND2_X1 U77604 ( .A1(n92056), .A2(n92057), .ZN(n92046) );
  AOI22_X1 U77605 ( .A1(n90517), .A2(n110190), .B1(n105646), .B2(n110192), 
        .ZN(n92057) );
  AOI22_X1 U77606 ( .A1(n105645), .A2(n110196), .B1(n90520), .B2(n110191), 
        .ZN(n92056) );
  NOR4_X1 U77607 ( .A1(n92058), .A2(n92059), .A3(n92060), .A4(n92061), .ZN(
        n92044) );
  NAND2_X1 U77608 ( .A1(n92062), .A2(n92063), .ZN(n92061) );
  AOI22_X1 U77609 ( .A1(n90527), .A2(n110171), .B1(n90528), .B2(n110174), .ZN(
        n92063) );
  AOI22_X1 U77610 ( .A1(n90529), .A2(n111035), .B1(n90530), .B2(n73341), .ZN(
        n92062) );
  NAND2_X1 U77611 ( .A1(n92064), .A2(n92065), .ZN(n92060) );
  AOI22_X1 U77612 ( .A1(n90533), .A2(n110180), .B1(n90534), .B2(n110170), .ZN(
        n92065) );
  AOI22_X1 U77613 ( .A1(n90535), .A2(n110173), .B1(n90536), .B2(n110177), .ZN(
        n92064) );
  NAND2_X1 U77614 ( .A1(n92066), .A2(n92067), .ZN(n92059) );
  AOI22_X1 U77615 ( .A1(n90539), .A2(n110176), .B1(n90540), .B2(n110181), .ZN(
        n92067) );
  AOI22_X1 U77616 ( .A1(n90541), .A2(n110183), .B1(n90542), .B2(n110179), .ZN(
        n92066) );
  NAND2_X1 U77617 ( .A1(n92068), .A2(n92069), .ZN(n92058) );
  AOI22_X1 U77618 ( .A1(n90545), .A2(n73359), .B1(n90546), .B2(n110175), .ZN(
        n92069) );
  AOI22_X1 U77619 ( .A1(n90547), .A2(n110178), .B1(n90548), .B2(n110182), .ZN(
        n92068) );
  AOI21_X1 U77620 ( .B1(n90295), .B2(n88092), .A(n92071), .ZN(n92070) );
  OAI21_X1 U77621 ( .B1(n92072), .B2(n105659), .A(n92073), .ZN(n92071) );
  OAI21_X1 U77622 ( .B1(n92074), .B2(n92075), .A(n105658), .ZN(n92073) );
  OAI21_X1 U77623 ( .B1(n101956), .B2(n105657), .A(n92076), .ZN(n92075) );
  AOI22_X1 U77624 ( .A1(n105656), .A2(n110002), .B1(n105655), .B2(n73116), 
        .ZN(n92076) );
  NAND2_X1 U77625 ( .A1(n92077), .A2(n92078), .ZN(n92074) );
  AOI22_X1 U77626 ( .A1(n105654), .A2(n110007), .B1(n105653), .B2(n110004), 
        .ZN(n92078) );
  AOI22_X1 U77627 ( .A1(n90311), .A2(n73114), .B1(n105652), .B2(n110003), .ZN(
        n92077) );
  NOR4_X1 U77628 ( .A1(n92079), .A2(n92080), .A3(n92081), .A4(n92082), .ZN(
        n92072) );
  NAND2_X1 U77629 ( .A1(n92083), .A2(n92084), .ZN(n92082) );
  NOR4_X1 U77630 ( .A1(n92085), .A2(n92086), .A3(n92087), .A4(n92088), .ZN(
        n92084) );
  NAND2_X1 U77631 ( .A1(n92089), .A2(n92090), .ZN(n92088) );
  AOI22_X1 U77632 ( .A1(n90325), .A2(n109983), .B1(n90326), .B2(n109984), .ZN(
        n92090) );
  AOI22_X1 U77633 ( .A1(n90327), .A2(n109992), .B1(n90328), .B2(n109990), .ZN(
        n92089) );
  NAND2_X1 U77634 ( .A1(n92091), .A2(n92092), .ZN(n92087) );
  AOI22_X1 U77635 ( .A1(n90331), .A2(n72983), .B1(n90332), .B2(n109987), .ZN(
        n92092) );
  AOI22_X1 U77636 ( .A1(n90333), .A2(n73087), .B1(n90334), .B2(n109904), .ZN(
        n92091) );
  NAND2_X1 U77637 ( .A1(n92093), .A2(n92094), .ZN(n92086) );
  AOI22_X1 U77638 ( .A1(n90337), .A2(n109908), .B1(n90338), .B2(n72987), .ZN(
        n92094) );
  AOI22_X1 U77639 ( .A1(n90339), .A2(n109988), .B1(n90340), .B2(n109985), .ZN(
        n92093) );
  NAND2_X1 U77640 ( .A1(n92095), .A2(n92096), .ZN(n92085) );
  AOI22_X1 U77641 ( .A1(n90343), .A2(n109906), .B1(n90344), .B2(n109910), .ZN(
        n92096) );
  AOI22_X1 U77642 ( .A1(n90345), .A2(n109909), .B1(n90346), .B2(n72989), .ZN(
        n92095) );
  NOR4_X1 U77643 ( .A1(n92097), .A2(n92098), .A3(n92099), .A4(n92100), .ZN(
        n92083) );
  NAND2_X1 U77644 ( .A1(n92101), .A2(n92102), .ZN(n92100) );
  AOI22_X1 U77645 ( .A1(n90353), .A2(n109993), .B1(n90354), .B2(n109996), .ZN(
        n92102) );
  AOI22_X1 U77646 ( .A1(n90355), .A2(n109997), .B1(n90356), .B2(n109999), .ZN(
        n92101) );
  NAND2_X1 U77647 ( .A1(n92103), .A2(n92104), .ZN(n92099) );
  AOI22_X1 U77648 ( .A1(n90359), .A2(n109998), .B1(n90360), .B2(n109994), .ZN(
        n92104) );
  AOI22_X1 U77649 ( .A1(n90361), .A2(n110000), .B1(n90362), .B2(n109995), .ZN(
        n92103) );
  NAND2_X1 U77650 ( .A1(n92105), .A2(n92106), .ZN(n92098) );
  AOI22_X1 U77651 ( .A1(n90365), .A2(n73097), .B1(n90366), .B2(n73096), .ZN(
        n92106) );
  AOI22_X1 U77652 ( .A1(n90367), .A2(n73099), .B1(n90368), .B2(n110001), .ZN(
        n92105) );
  NAND2_X1 U77653 ( .A1(n92107), .A2(n92108), .ZN(n92097) );
  AOI22_X1 U77654 ( .A1(n90371), .A2(n109986), .B1(n90372), .B2(n109991), .ZN(
        n92108) );
  AOI22_X1 U77655 ( .A1(n90373), .A2(n73094), .B1(n90374), .B2(n109989), .ZN(
        n92107) );
  NAND2_X1 U77656 ( .A1(n92109), .A2(n92110), .ZN(n92081) );
  NOR4_X1 U77657 ( .A1(n92111), .A2(n92112), .A3(n92113), .A4(n92114), .ZN(
        n92110) );
  NAND2_X1 U77658 ( .A1(n92115), .A2(n92116), .ZN(n92114) );
  AOI22_X1 U77659 ( .A1(n90383), .A2(n109919), .B1(n90384), .B2(n109921), .ZN(
        n92116) );
  AOI22_X1 U77660 ( .A1(n90385), .A2(n73012), .B1(n90386), .B2(n109920), .ZN(
        n92115) );
  NAND2_X1 U77661 ( .A1(n92117), .A2(n92118), .ZN(n92113) );
  AOI22_X1 U77662 ( .A1(n90389), .A2(n73016), .B1(n90390), .B2(n73018), .ZN(
        n92118) );
  AOI22_X1 U77663 ( .A1(n90391), .A2(n109927), .B1(n90392), .B2(n109928), .ZN(
        n92117) );
  NAND2_X1 U77664 ( .A1(n92119), .A2(n92120), .ZN(n92112) );
  AOI22_X1 U77665 ( .A1(n90395), .A2(n109924), .B1(n90396), .B2(n109926), .ZN(
        n92120) );
  AOI22_X1 U77666 ( .A1(n90397), .A2(n73017), .B1(n90398), .B2(n109925), .ZN(
        n92119) );
  NAND2_X1 U77667 ( .A1(n92121), .A2(n92122), .ZN(n92111) );
  AOI22_X1 U77668 ( .A1(n90401), .A2(n109933), .B1(n90402), .B2(n73023), .ZN(
        n92122) );
  AOI22_X1 U77669 ( .A1(n90403), .A2(n109932), .B1(n90404), .B2(n73021), .ZN(
        n92121) );
  NOR4_X1 U77670 ( .A1(n92123), .A2(n92124), .A3(n92125), .A4(n92126), .ZN(
        n92109) );
  NAND2_X1 U77671 ( .A1(n92127), .A2(n92128), .ZN(n92126) );
  AOI22_X1 U77672 ( .A1(n90411), .A2(n109914), .B1(n90412), .B2(n109905), .ZN(
        n92128) );
  AOI22_X1 U77673 ( .A1(n90413), .A2(n109907), .B1(n90414), .B2(n72995), .ZN(
        n92127) );
  NAND2_X1 U77674 ( .A1(n92129), .A2(n92130), .ZN(n92125) );
  AOI22_X1 U77675 ( .A1(n90417), .A2(n109912), .B1(n90418), .B2(n109916), .ZN(
        n92130) );
  AOI22_X1 U77676 ( .A1(n90419), .A2(n109918), .B1(n90420), .B2(n109915), .ZN(
        n92129) );
  NAND2_X1 U77677 ( .A1(n92131), .A2(n92132), .ZN(n92124) );
  AOI22_X1 U77678 ( .A1(n90423), .A2(n73004), .B1(n90424), .B2(n109911), .ZN(
        n92132) );
  AOI22_X1 U77679 ( .A1(n90425), .A2(n109913), .B1(n90426), .B2(n109917), .ZN(
        n92131) );
  NAND2_X1 U77680 ( .A1(n92133), .A2(n92134), .ZN(n92123) );
  AOI22_X1 U77681 ( .A1(n90429), .A2(n109923), .B1(n90430), .B2(n73008), .ZN(
        n92134) );
  AOI22_X1 U77682 ( .A1(n90431), .A2(n73006), .B1(n90432), .B2(n109922), .ZN(
        n92133) );
  NAND2_X1 U77683 ( .A1(n92135), .A2(n92136), .ZN(n92080) );
  NOR4_X1 U77684 ( .A1(n92137), .A2(n92138), .A3(n92139), .A4(n92140), .ZN(
        n92136) );
  NAND2_X1 U77685 ( .A1(n92141), .A2(n92142), .ZN(n92140) );
  AOI22_X1 U77686 ( .A1(n90441), .A2(n73046), .B1(n90442), .B2(n109943), .ZN(
        n92142) );
  AOI22_X1 U77687 ( .A1(n90443), .A2(n109947), .B1(n90444), .B2(n109946), .ZN(
        n92141) );
  NAND2_X1 U77688 ( .A1(n92143), .A2(n92144), .ZN(n92139) );
  AOI22_X1 U77689 ( .A1(n90447), .A2(n109952), .B1(n90448), .B2(n109951), .ZN(
        n92144) );
  AOI22_X1 U77690 ( .A1(n90449), .A2(n109942), .B1(n90450), .B2(n109944), .ZN(
        n92143) );
  NAND2_X1 U77691 ( .A1(n92145), .A2(n92146), .ZN(n92138) );
  AOI22_X1 U77692 ( .A1(n90453), .A2(n109953), .B1(n90454), .B2(n109949), .ZN(
        n92146) );
  AOI22_X1 U77693 ( .A1(n90455), .A2(n73050), .B1(n90456), .B2(n73052), .ZN(
        n92145) );
  NAND2_X1 U77694 ( .A1(n92147), .A2(n92148), .ZN(n92137) );
  AOI22_X1 U77695 ( .A1(n90459), .A2(n109956), .B1(n90460), .B2(n73058), .ZN(
        n92148) );
  AOI22_X1 U77696 ( .A1(n90461), .A2(n109948), .B1(n90462), .B2(n109950), .ZN(
        n92147) );
  NOR4_X1 U77697 ( .A1(n92149), .A2(n92150), .A3(n92151), .A4(n92152), .ZN(
        n92135) );
  NAND2_X1 U77698 ( .A1(n92153), .A2(n92154), .ZN(n92152) );
  AOI22_X1 U77699 ( .A1(n90469), .A2(n109931), .B1(n90470), .B2(n109936), .ZN(
        n92154) );
  AOI22_X1 U77700 ( .A1(n90471), .A2(n109930), .B1(n90472), .B2(n73026), .ZN(
        n92153) );
  NAND2_X1 U77701 ( .A1(n92155), .A2(n92156), .ZN(n92151) );
  AOI22_X1 U77702 ( .A1(n90475), .A2(n73035), .B1(n90476), .B2(n109938), .ZN(
        n92156) );
  AOI22_X1 U77703 ( .A1(n90477), .A2(n109939), .B1(n90478), .B2(n109929), .ZN(
        n92155) );
  NAND2_X1 U77704 ( .A1(n92157), .A2(n92158), .ZN(n92150) );
  AOI22_X1 U77705 ( .A1(n90481), .A2(n109937), .B1(n90482), .B2(n109941), .ZN(
        n92158) );
  AOI22_X1 U77706 ( .A1(n90483), .A2(n109935), .B1(n90484), .B2(n109940), .ZN(
        n92157) );
  NAND2_X1 U77707 ( .A1(n92159), .A2(n92160), .ZN(n92149) );
  AOI22_X1 U77708 ( .A1(n90487), .A2(n73040), .B1(n90488), .B2(n109945), .ZN(
        n92160) );
  AOI22_X1 U77709 ( .A1(n90489), .A2(n73038), .B1(n90490), .B2(n109934), .ZN(
        n92159) );
  NAND2_X1 U77710 ( .A1(n92161), .A2(n92162), .ZN(n92079) );
  NOR4_X1 U77711 ( .A1(n92163), .A2(n92164), .A3(n92165), .A4(n92166), .ZN(
        n92162) );
  NAND2_X1 U77712 ( .A1(n92167), .A2(n92168), .ZN(n92166) );
  AOI22_X1 U77713 ( .A1(n90499), .A2(n109974), .B1(n90500), .B2(n109973), .ZN(
        n92168) );
  AOI22_X1 U77714 ( .A1(n90501), .A2(n73074), .B1(n90502), .B2(n109971), .ZN(
        n92167) );
  NAND2_X1 U77715 ( .A1(n92169), .A2(n92170), .ZN(n92165) );
  AOI22_X1 U77716 ( .A1(n90505), .A2(n109969), .B1(n90506), .B2(n109972), .ZN(
        n92170) );
  AOI22_X1 U77717 ( .A1(n105651), .A2(n73080), .B1(n90508), .B2(n109970), .ZN(
        n92169) );
  NAND2_X1 U77718 ( .A1(n92171), .A2(n92172), .ZN(n92164) );
  AOI22_X1 U77719 ( .A1(n105650), .A2(n109980), .B1(n105649), .B2(n73086), 
        .ZN(n92172) );
  AOI22_X1 U77720 ( .A1(n105648), .A2(n109978), .B1(n105647), .B2(n109979), 
        .ZN(n92171) );
  NAND2_X1 U77721 ( .A1(n92173), .A2(n92174), .ZN(n92163) );
  AOI22_X1 U77722 ( .A1(n90517), .A2(n109975), .B1(n105646), .B2(n109977), 
        .ZN(n92174) );
  AOI22_X1 U77723 ( .A1(n105645), .A2(n109981), .B1(n90520), .B2(n109976), 
        .ZN(n92173) );
  NOR4_X1 U77724 ( .A1(n92175), .A2(n92176), .A3(n92177), .A4(n92178), .ZN(
        n92161) );
  NAND2_X1 U77725 ( .A1(n92179), .A2(n92180), .ZN(n92178) );
  AOI22_X1 U77726 ( .A1(n90527), .A2(n109955), .B1(n90528), .B2(n109959), .ZN(
        n92180) );
  AOI22_X1 U77727 ( .A1(n90529), .A2(n109958), .B1(n90530), .B2(n73057), .ZN(
        n92179) );
  NAND2_X1 U77728 ( .A1(n92181), .A2(n92182), .ZN(n92177) );
  AOI22_X1 U77729 ( .A1(n90533), .A2(n109965), .B1(n90534), .B2(n109954), .ZN(
        n92182) );
  AOI22_X1 U77730 ( .A1(n90535), .A2(n109957), .B1(n90536), .B2(n109962), .ZN(
        n92181) );
  NAND2_X1 U77731 ( .A1(n92183), .A2(n92184), .ZN(n92176) );
  AOI22_X1 U77732 ( .A1(n90539), .A2(n109961), .B1(n90540), .B2(n109966), .ZN(
        n92184) );
  AOI22_X1 U77733 ( .A1(n90541), .A2(n109968), .B1(n90542), .B2(n109964), .ZN(
        n92183) );
  NAND2_X1 U77734 ( .A1(n92185), .A2(n92186), .ZN(n92175) );
  AOI22_X1 U77735 ( .A1(n90545), .A2(n73075), .B1(n90546), .B2(n109960), .ZN(
        n92186) );
  AOI22_X1 U77736 ( .A1(n90547), .A2(n109963), .B1(n90548), .B2(n109967), .ZN(
        n92185) );
  AOI21_X1 U77737 ( .B1(n90295), .B2(n88210), .A(n92188), .ZN(n92187) );
  OAI21_X1 U77738 ( .B1(n92189), .B2(n105659), .A(n92190), .ZN(n92188) );
  OAI21_X1 U77739 ( .B1(n92191), .B2(n92192), .A(n105658), .ZN(n92190) );
  OAI21_X1 U77740 ( .B1(n101940), .B2(n90303), .A(n92193), .ZN(n92192) );
  AOI22_X1 U77741 ( .A1(n105656), .A2(n109885), .B1(n105655), .B2(n72966), 
        .ZN(n92193) );
  NAND2_X1 U77742 ( .A1(n92194), .A2(n92195), .ZN(n92191) );
  AOI22_X1 U77743 ( .A1(n105654), .A2(n109890), .B1(n105653), .B2(n109887), 
        .ZN(n92195) );
  AOI22_X1 U77744 ( .A1(n90311), .A2(n72964), .B1(n105652), .B2(n109886), .ZN(
        n92194) );
  NOR4_X1 U77745 ( .A1(n92196), .A2(n92197), .A3(n92198), .A4(n92199), .ZN(
        n92189) );
  NAND2_X1 U77746 ( .A1(n92200), .A2(n92201), .ZN(n92199) );
  NOR4_X1 U77747 ( .A1(n92202), .A2(n92203), .A3(n92204), .A4(n92205), .ZN(
        n92201) );
  NAND2_X1 U77748 ( .A1(n92206), .A2(n92207), .ZN(n92205) );
  AOI22_X1 U77749 ( .A1(n90325), .A2(n109866), .B1(n90326), .B2(n109867), .ZN(
        n92207) );
  AOI22_X1 U77750 ( .A1(n90327), .A2(n109875), .B1(n90328), .B2(n109873), .ZN(
        n92206) );
  NAND2_X1 U77751 ( .A1(n92208), .A2(n92209), .ZN(n92204) );
  AOI22_X1 U77752 ( .A1(n90331), .A2(n72833), .B1(n90332), .B2(n109870), .ZN(
        n92209) );
  AOI22_X1 U77753 ( .A1(n90333), .A2(n72937), .B1(n90334), .B2(n109786), .ZN(
        n92208) );
  NAND2_X1 U77754 ( .A1(n92210), .A2(n92211), .ZN(n92203) );
  AOI22_X1 U77755 ( .A1(n90337), .A2(n109790), .B1(n90338), .B2(n72837), .ZN(
        n92211) );
  AOI22_X1 U77756 ( .A1(n90339), .A2(n109871), .B1(n90340), .B2(n109868), .ZN(
        n92210) );
  NAND2_X1 U77757 ( .A1(n92212), .A2(n92213), .ZN(n92202) );
  AOI22_X1 U77758 ( .A1(n90343), .A2(n109788), .B1(n90344), .B2(n109792), .ZN(
        n92213) );
  AOI22_X1 U77759 ( .A1(n90345), .A2(n109791), .B1(n90346), .B2(n72839), .ZN(
        n92212) );
  NOR4_X1 U77760 ( .A1(n92214), .A2(n92215), .A3(n92216), .A4(n92217), .ZN(
        n92200) );
  NAND2_X1 U77761 ( .A1(n92218), .A2(n92219), .ZN(n92217) );
  AOI22_X1 U77762 ( .A1(n90353), .A2(n109876), .B1(n90354), .B2(n109879), .ZN(
        n92219) );
  AOI22_X1 U77763 ( .A1(n90355), .A2(n109880), .B1(n90356), .B2(n109882), .ZN(
        n92218) );
  NAND2_X1 U77764 ( .A1(n92220), .A2(n92221), .ZN(n92216) );
  AOI22_X1 U77765 ( .A1(n90359), .A2(n109881), .B1(n90360), .B2(n109877), .ZN(
        n92221) );
  AOI22_X1 U77766 ( .A1(n90361), .A2(n109883), .B1(n90362), .B2(n109878), .ZN(
        n92220) );
  NAND2_X1 U77767 ( .A1(n92222), .A2(n92223), .ZN(n92215) );
  AOI22_X1 U77768 ( .A1(n90365), .A2(n72947), .B1(n90366), .B2(n72946), .ZN(
        n92223) );
  AOI22_X1 U77769 ( .A1(n90367), .A2(n72949), .B1(n90368), .B2(n109884), .ZN(
        n92222) );
  NAND2_X1 U77770 ( .A1(n92224), .A2(n92225), .ZN(n92214) );
  AOI22_X1 U77771 ( .A1(n90371), .A2(n109869), .B1(n90372), .B2(n109874), .ZN(
        n92225) );
  AOI22_X1 U77772 ( .A1(n90373), .A2(n72944), .B1(n90374), .B2(n109872), .ZN(
        n92224) );
  NAND2_X1 U77773 ( .A1(n92226), .A2(n92227), .ZN(n92198) );
  NOR4_X1 U77774 ( .A1(n92228), .A2(n92229), .A3(n92230), .A4(n92231), .ZN(
        n92227) );
  NAND2_X1 U77775 ( .A1(n92232), .A2(n92233), .ZN(n92231) );
  AOI22_X1 U77776 ( .A1(n90383), .A2(n109801), .B1(n90384), .B2(n109803), .ZN(
        n92233) );
  AOI22_X1 U77777 ( .A1(n90385), .A2(n72862), .B1(n90386), .B2(n109802), .ZN(
        n92232) );
  NAND2_X1 U77778 ( .A1(n92234), .A2(n92235), .ZN(n92230) );
  AOI22_X1 U77779 ( .A1(n90389), .A2(n72866), .B1(n90390), .B2(n72868), .ZN(
        n92235) );
  AOI22_X1 U77780 ( .A1(n90391), .A2(n109809), .B1(n90392), .B2(n109810), .ZN(
        n92234) );
  NAND2_X1 U77781 ( .A1(n92236), .A2(n92237), .ZN(n92229) );
  AOI22_X1 U77782 ( .A1(n90395), .A2(n109806), .B1(n90396), .B2(n109808), .ZN(
        n92237) );
  AOI22_X1 U77783 ( .A1(n90397), .A2(n109811), .B1(n90398), .B2(n109807), .ZN(
        n92236) );
  NAND2_X1 U77784 ( .A1(n92238), .A2(n92239), .ZN(n92228) );
  AOI22_X1 U77785 ( .A1(n90401), .A2(n109816), .B1(n90402), .B2(n72873), .ZN(
        n92239) );
  AOI22_X1 U77786 ( .A1(n90403), .A2(n109815), .B1(n90404), .B2(n72871), .ZN(
        n92238) );
  NOR4_X1 U77787 ( .A1(n92240), .A2(n92241), .A3(n92242), .A4(n92243), .ZN(
        n92226) );
  NAND2_X1 U77788 ( .A1(n92244), .A2(n92245), .ZN(n92243) );
  AOI22_X1 U77789 ( .A1(n90411), .A2(n109796), .B1(n90412), .B2(n109787), .ZN(
        n92245) );
  AOI22_X1 U77790 ( .A1(n90413), .A2(n109789), .B1(n90414), .B2(n72845), .ZN(
        n92244) );
  NAND2_X1 U77791 ( .A1(n92246), .A2(n92247), .ZN(n92242) );
  AOI22_X1 U77792 ( .A1(n90417), .A2(n109794), .B1(n90418), .B2(n109798), .ZN(
        n92247) );
  AOI22_X1 U77793 ( .A1(n90419), .A2(n109800), .B1(n90420), .B2(n109797), .ZN(
        n92246) );
  NAND2_X1 U77794 ( .A1(n92248), .A2(n92249), .ZN(n92241) );
  AOI22_X1 U77795 ( .A1(n90423), .A2(n72854), .B1(n90424), .B2(n109793), .ZN(
        n92249) );
  AOI22_X1 U77796 ( .A1(n90425), .A2(n109795), .B1(n90426), .B2(n109799), .ZN(
        n92248) );
  NAND2_X1 U77797 ( .A1(n92250), .A2(n92251), .ZN(n92240) );
  AOI22_X1 U77798 ( .A1(n90429), .A2(n109805), .B1(n90430), .B2(n72858), .ZN(
        n92251) );
  AOI22_X1 U77799 ( .A1(n90431), .A2(n72856), .B1(n90432), .B2(n109804), .ZN(
        n92250) );
  NAND2_X1 U77800 ( .A1(n92252), .A2(n92253), .ZN(n92197) );
  NOR4_X1 U77801 ( .A1(n92254), .A2(n92255), .A3(n92256), .A4(n92257), .ZN(
        n92253) );
  NAND2_X1 U77802 ( .A1(n92258), .A2(n92259), .ZN(n92257) );
  AOI22_X1 U77803 ( .A1(n90441), .A2(n72896), .B1(n90442), .B2(n109826), .ZN(
        n92259) );
  AOI22_X1 U77804 ( .A1(n90443), .A2(n109830), .B1(n90444), .B2(n109829), .ZN(
        n92258) );
  NAND2_X1 U77805 ( .A1(n92260), .A2(n92261), .ZN(n92256) );
  AOI22_X1 U77806 ( .A1(n90447), .A2(n109835), .B1(n90448), .B2(n109834), .ZN(
        n92261) );
  AOI22_X1 U77807 ( .A1(n90449), .A2(n109825), .B1(n90450), .B2(n109827), .ZN(
        n92260) );
  NAND2_X1 U77808 ( .A1(n92262), .A2(n92263), .ZN(n92255) );
  AOI22_X1 U77809 ( .A1(n90453), .A2(n109836), .B1(n90454), .B2(n109832), .ZN(
        n92263) );
  AOI22_X1 U77810 ( .A1(n90455), .A2(n72900), .B1(n90456), .B2(n72902), .ZN(
        n92262) );
  NAND2_X1 U77811 ( .A1(n92264), .A2(n92265), .ZN(n92254) );
  AOI22_X1 U77812 ( .A1(n90459), .A2(n109839), .B1(n90460), .B2(n72908), .ZN(
        n92265) );
  AOI22_X1 U77813 ( .A1(n90461), .A2(n109831), .B1(n90462), .B2(n109833), .ZN(
        n92264) );
  NOR4_X1 U77814 ( .A1(n92266), .A2(n92267), .A3(n92268), .A4(n92269), .ZN(
        n92252) );
  NAND2_X1 U77815 ( .A1(n92270), .A2(n92271), .ZN(n92269) );
  AOI22_X1 U77816 ( .A1(n90469), .A2(n109814), .B1(n90470), .B2(n109819), .ZN(
        n92271) );
  AOI22_X1 U77817 ( .A1(n90471), .A2(n109813), .B1(n90472), .B2(n72876), .ZN(
        n92270) );
  NAND2_X1 U77818 ( .A1(n92272), .A2(n92273), .ZN(n92268) );
  AOI22_X1 U77819 ( .A1(n90475), .A2(n72885), .B1(n90476), .B2(n109821), .ZN(
        n92273) );
  AOI22_X1 U77820 ( .A1(n90477), .A2(n109822), .B1(n90478), .B2(n109812), .ZN(
        n92272) );
  NAND2_X1 U77821 ( .A1(n92274), .A2(n92275), .ZN(n92267) );
  AOI22_X1 U77822 ( .A1(n90481), .A2(n109820), .B1(n90482), .B2(n109824), .ZN(
        n92275) );
  AOI22_X1 U77823 ( .A1(n90483), .A2(n109818), .B1(n90484), .B2(n109823), .ZN(
        n92274) );
  NAND2_X1 U77824 ( .A1(n92276), .A2(n92277), .ZN(n92266) );
  AOI22_X1 U77825 ( .A1(n90487), .A2(n72890), .B1(n90488), .B2(n109828), .ZN(
        n92277) );
  AOI22_X1 U77826 ( .A1(n90489), .A2(n72888), .B1(n90490), .B2(n109817), .ZN(
        n92276) );
  NAND2_X1 U77827 ( .A1(n92278), .A2(n92279), .ZN(n92196) );
  NOR4_X1 U77828 ( .A1(n92280), .A2(n92281), .A3(n92282), .A4(n92283), .ZN(
        n92279) );
  NAND2_X1 U77829 ( .A1(n92284), .A2(n92285), .ZN(n92283) );
  AOI22_X1 U77830 ( .A1(n90499), .A2(n109857), .B1(n90500), .B2(n109856), .ZN(
        n92285) );
  AOI22_X1 U77831 ( .A1(n90501), .A2(n72924), .B1(n90502), .B2(n109854), .ZN(
        n92284) );
  NAND2_X1 U77832 ( .A1(n92286), .A2(n92287), .ZN(n92282) );
  AOI22_X1 U77833 ( .A1(n90505), .A2(n109852), .B1(n90506), .B2(n109855), .ZN(
        n92287) );
  AOI22_X1 U77834 ( .A1(n105651), .A2(n72930), .B1(n90508), .B2(n109853), .ZN(
        n92286) );
  NAND2_X1 U77835 ( .A1(n92288), .A2(n92289), .ZN(n92281) );
  AOI22_X1 U77836 ( .A1(n105650), .A2(n109863), .B1(n105649), .B2(n72936), 
        .ZN(n92289) );
  AOI22_X1 U77837 ( .A1(n105648), .A2(n109861), .B1(n105647), .B2(n109862), 
        .ZN(n92288) );
  NAND2_X1 U77838 ( .A1(n92290), .A2(n92291), .ZN(n92280) );
  AOI22_X1 U77839 ( .A1(n90517), .A2(n109858), .B1(n105646), .B2(n109860), 
        .ZN(n92291) );
  AOI22_X1 U77840 ( .A1(n105645), .A2(n109864), .B1(n105644), .B2(n109859), 
        .ZN(n92290) );
  NOR4_X1 U77841 ( .A1(n92292), .A2(n92293), .A3(n92294), .A4(n92295), .ZN(
        n92278) );
  NAND2_X1 U77842 ( .A1(n92296), .A2(n92297), .ZN(n92295) );
  AOI22_X1 U77843 ( .A1(n90527), .A2(n109838), .B1(n90528), .B2(n109842), .ZN(
        n92297) );
  AOI22_X1 U77844 ( .A1(n90529), .A2(n109841), .B1(n90530), .B2(n72907), .ZN(
        n92296) );
  NAND2_X1 U77845 ( .A1(n92298), .A2(n92299), .ZN(n92294) );
  AOI22_X1 U77846 ( .A1(n90533), .A2(n109848), .B1(n90534), .B2(n109837), .ZN(
        n92299) );
  AOI22_X1 U77847 ( .A1(n90535), .A2(n109840), .B1(n90536), .B2(n109845), .ZN(
        n92298) );
  NAND2_X1 U77848 ( .A1(n92300), .A2(n92301), .ZN(n92293) );
  AOI22_X1 U77849 ( .A1(n90539), .A2(n109844), .B1(n90540), .B2(n109849), .ZN(
        n92301) );
  AOI22_X1 U77850 ( .A1(n90541), .A2(n109851), .B1(n90542), .B2(n109847), .ZN(
        n92300) );
  NAND2_X1 U77851 ( .A1(n92302), .A2(n92303), .ZN(n92292) );
  AOI22_X1 U77852 ( .A1(n90545), .A2(n72925), .B1(n90546), .B2(n109843), .ZN(
        n92303) );
  AOI22_X1 U77853 ( .A1(n90547), .A2(n109846), .B1(n90548), .B2(n109850), .ZN(
        n92302) );
  AOI21_X1 U77854 ( .B1(n90295), .B2(n88328), .A(n92305), .ZN(n92304) );
  OAI21_X1 U77855 ( .B1(n92306), .B2(n105659), .A(n92307), .ZN(n92305) );
  OAI21_X1 U77856 ( .B1(n92308), .B2(n92309), .A(n105658), .ZN(n92307) );
  OAI21_X1 U77857 ( .B1(n101924), .B2(n105657), .A(n92310), .ZN(n92309) );
  AOI22_X1 U77858 ( .A1(n105656), .A2(n108259), .B1(n105655), .B2(n70862), 
        .ZN(n92310) );
  NAND2_X1 U77859 ( .A1(n92311), .A2(n92312), .ZN(n92308) );
  AOI22_X1 U77860 ( .A1(n105654), .A2(n108264), .B1(n105653), .B2(n108261), 
        .ZN(n92312) );
  AOI22_X1 U77861 ( .A1(n90311), .A2(n70860), .B1(n105652), .B2(n108260), .ZN(
        n92311) );
  NOR4_X1 U77862 ( .A1(n92313), .A2(n92314), .A3(n92315), .A4(n92316), .ZN(
        n92306) );
  NAND2_X1 U77863 ( .A1(n92317), .A2(n92318), .ZN(n92316) );
  NOR4_X1 U77864 ( .A1(n92319), .A2(n92320), .A3(n92321), .A4(n92322), .ZN(
        n92318) );
  NAND2_X1 U77865 ( .A1(n92323), .A2(n92324), .ZN(n92322) );
  AOI22_X1 U77866 ( .A1(n90325), .A2(n108240), .B1(n90326), .B2(n108241), .ZN(
        n92324) );
  AOI22_X1 U77867 ( .A1(n90327), .A2(n108249), .B1(n90328), .B2(n108247), .ZN(
        n92323) );
  NAND2_X1 U77868 ( .A1(n92325), .A2(n92326), .ZN(n92321) );
  AOI22_X1 U77869 ( .A1(n90331), .A2(n70729), .B1(n90332), .B2(n108244), .ZN(
        n92326) );
  AOI22_X1 U77870 ( .A1(n90333), .A2(n70833), .B1(n90334), .B2(n108160), .ZN(
        n92325) );
  NAND2_X1 U77871 ( .A1(n92327), .A2(n92328), .ZN(n92320) );
  AOI22_X1 U77872 ( .A1(n90337), .A2(n108164), .B1(n90338), .B2(n70733), .ZN(
        n92328) );
  AOI22_X1 U77873 ( .A1(n90339), .A2(n108245), .B1(n90340), .B2(n108242), .ZN(
        n92327) );
  NAND2_X1 U77874 ( .A1(n92329), .A2(n92330), .ZN(n92319) );
  AOI22_X1 U77875 ( .A1(n90343), .A2(n108162), .B1(n90344), .B2(n108166), .ZN(
        n92330) );
  AOI22_X1 U77876 ( .A1(n90345), .A2(n108165), .B1(n90346), .B2(n70735), .ZN(
        n92329) );
  NOR4_X1 U77877 ( .A1(n92331), .A2(n92332), .A3(n92333), .A4(n92334), .ZN(
        n92317) );
  NAND2_X1 U77878 ( .A1(n92335), .A2(n92336), .ZN(n92334) );
  AOI22_X1 U77879 ( .A1(n90353), .A2(n108250), .B1(n90354), .B2(n108253), .ZN(
        n92336) );
  AOI22_X1 U77880 ( .A1(n90355), .A2(n108254), .B1(n90356), .B2(n108256), .ZN(
        n92335) );
  NAND2_X1 U77881 ( .A1(n92337), .A2(n92338), .ZN(n92333) );
  AOI22_X1 U77882 ( .A1(n90359), .A2(n108255), .B1(n90360), .B2(n108251), .ZN(
        n92338) );
  AOI22_X1 U77883 ( .A1(n90361), .A2(n108257), .B1(n90362), .B2(n108252), .ZN(
        n92337) );
  NAND2_X1 U77884 ( .A1(n92339), .A2(n92340), .ZN(n92332) );
  AOI22_X1 U77885 ( .A1(n90365), .A2(n70843), .B1(n90366), .B2(n70842), .ZN(
        n92340) );
  AOI22_X1 U77886 ( .A1(n90367), .A2(n70845), .B1(n90368), .B2(n108258), .ZN(
        n92339) );
  NAND2_X1 U77887 ( .A1(n92341), .A2(n92342), .ZN(n92331) );
  AOI22_X1 U77888 ( .A1(n90371), .A2(n108243), .B1(n90372), .B2(n108248), .ZN(
        n92342) );
  AOI22_X1 U77889 ( .A1(n90373), .A2(n70840), .B1(n90374), .B2(n108246), .ZN(
        n92341) );
  NAND2_X1 U77890 ( .A1(n92343), .A2(n92344), .ZN(n92315) );
  NOR4_X1 U77891 ( .A1(n92345), .A2(n92346), .A3(n92347), .A4(n92348), .ZN(
        n92344) );
  NAND2_X1 U77892 ( .A1(n92349), .A2(n92350), .ZN(n92348) );
  AOI22_X1 U77893 ( .A1(n90383), .A2(n108175), .B1(n90384), .B2(n108177), .ZN(
        n92350) );
  AOI22_X1 U77894 ( .A1(n90385), .A2(n70758), .B1(n90386), .B2(n108176), .ZN(
        n92349) );
  NAND2_X1 U77895 ( .A1(n92351), .A2(n92352), .ZN(n92347) );
  AOI22_X1 U77896 ( .A1(n90389), .A2(n70762), .B1(n90390), .B2(n70764), .ZN(
        n92352) );
  AOI22_X1 U77897 ( .A1(n90391), .A2(n108183), .B1(n90392), .B2(n108184), .ZN(
        n92351) );
  NAND2_X1 U77898 ( .A1(n92353), .A2(n92354), .ZN(n92346) );
  AOI22_X1 U77899 ( .A1(n90395), .A2(n108180), .B1(n90396), .B2(n108182), .ZN(
        n92354) );
  AOI22_X1 U77900 ( .A1(n90397), .A2(n108185), .B1(n90398), .B2(n108181), .ZN(
        n92353) );
  NAND2_X1 U77901 ( .A1(n92355), .A2(n92356), .ZN(n92345) );
  AOI22_X1 U77902 ( .A1(n90401), .A2(n108190), .B1(n90402), .B2(n70769), .ZN(
        n92356) );
  AOI22_X1 U77903 ( .A1(n90403), .A2(n108189), .B1(n90404), .B2(n70767), .ZN(
        n92355) );
  NOR4_X1 U77904 ( .A1(n92357), .A2(n92358), .A3(n92359), .A4(n92360), .ZN(
        n92343) );
  NAND2_X1 U77905 ( .A1(n92361), .A2(n92362), .ZN(n92360) );
  AOI22_X1 U77906 ( .A1(n90411), .A2(n108170), .B1(n90412), .B2(n108161), .ZN(
        n92362) );
  AOI22_X1 U77907 ( .A1(n90413), .A2(n108163), .B1(n90414), .B2(n70741), .ZN(
        n92361) );
  NAND2_X1 U77908 ( .A1(n92363), .A2(n92364), .ZN(n92359) );
  AOI22_X1 U77909 ( .A1(n90417), .A2(n108168), .B1(n90418), .B2(n108172), .ZN(
        n92364) );
  AOI22_X1 U77910 ( .A1(n90419), .A2(n108174), .B1(n90420), .B2(n108171), .ZN(
        n92363) );
  NAND2_X1 U77911 ( .A1(n92365), .A2(n92366), .ZN(n92358) );
  AOI22_X1 U77912 ( .A1(n90423), .A2(n70750), .B1(n90424), .B2(n108167), .ZN(
        n92366) );
  AOI22_X1 U77913 ( .A1(n90425), .A2(n108169), .B1(n90426), .B2(n108173), .ZN(
        n92365) );
  NAND2_X1 U77914 ( .A1(n92367), .A2(n92368), .ZN(n92357) );
  AOI22_X1 U77915 ( .A1(n90429), .A2(n108179), .B1(n90430), .B2(n70754), .ZN(
        n92368) );
  AOI22_X1 U77916 ( .A1(n90431), .A2(n70752), .B1(n90432), .B2(n108178), .ZN(
        n92367) );
  NAND2_X1 U77917 ( .A1(n92369), .A2(n92370), .ZN(n92314) );
  NOR4_X1 U77918 ( .A1(n92371), .A2(n92372), .A3(n92373), .A4(n92374), .ZN(
        n92370) );
  NAND2_X1 U77919 ( .A1(n92375), .A2(n92376), .ZN(n92374) );
  AOI22_X1 U77920 ( .A1(n90441), .A2(n70792), .B1(n90442), .B2(n108200), .ZN(
        n92376) );
  AOI22_X1 U77921 ( .A1(n90443), .A2(n108204), .B1(n90444), .B2(n108203), .ZN(
        n92375) );
  NAND2_X1 U77922 ( .A1(n92377), .A2(n92378), .ZN(n92373) );
  AOI22_X1 U77923 ( .A1(n90447), .A2(n108209), .B1(n90448), .B2(n108208), .ZN(
        n92378) );
  AOI22_X1 U77924 ( .A1(n90449), .A2(n108199), .B1(n90450), .B2(n108201), .ZN(
        n92377) );
  NAND2_X1 U77925 ( .A1(n92379), .A2(n92380), .ZN(n92372) );
  AOI22_X1 U77926 ( .A1(n90453), .A2(n108210), .B1(n90454), .B2(n108206), .ZN(
        n92380) );
  AOI22_X1 U77927 ( .A1(n90455), .A2(n70796), .B1(n90456), .B2(n70798), .ZN(
        n92379) );
  NAND2_X1 U77928 ( .A1(n92381), .A2(n92382), .ZN(n92371) );
  AOI22_X1 U77929 ( .A1(n90459), .A2(n108213), .B1(n90460), .B2(n70804), .ZN(
        n92382) );
  AOI22_X1 U77930 ( .A1(n90461), .A2(n108205), .B1(n90462), .B2(n108207), .ZN(
        n92381) );
  NOR4_X1 U77931 ( .A1(n92383), .A2(n92384), .A3(n92385), .A4(n92386), .ZN(
        n92369) );
  NAND2_X1 U77932 ( .A1(n92387), .A2(n92388), .ZN(n92386) );
  AOI22_X1 U77933 ( .A1(n90469), .A2(n108188), .B1(n90470), .B2(n108193), .ZN(
        n92388) );
  AOI22_X1 U77934 ( .A1(n90471), .A2(n108187), .B1(n90472), .B2(n70772), .ZN(
        n92387) );
  NAND2_X1 U77935 ( .A1(n92389), .A2(n92390), .ZN(n92385) );
  AOI22_X1 U77936 ( .A1(n90475), .A2(n70781), .B1(n90476), .B2(n108195), .ZN(
        n92390) );
  AOI22_X1 U77937 ( .A1(n90477), .A2(n108196), .B1(n90478), .B2(n108186), .ZN(
        n92389) );
  NAND2_X1 U77938 ( .A1(n92391), .A2(n92392), .ZN(n92384) );
  AOI22_X1 U77939 ( .A1(n90481), .A2(n108194), .B1(n90482), .B2(n108198), .ZN(
        n92392) );
  AOI22_X1 U77940 ( .A1(n90483), .A2(n108192), .B1(n90484), .B2(n108197), .ZN(
        n92391) );
  NAND2_X1 U77941 ( .A1(n92393), .A2(n92394), .ZN(n92383) );
  AOI22_X1 U77942 ( .A1(n90487), .A2(n70786), .B1(n90488), .B2(n108202), .ZN(
        n92394) );
  AOI22_X1 U77943 ( .A1(n90489), .A2(n70784), .B1(n90490), .B2(n108191), .ZN(
        n92393) );
  NAND2_X1 U77944 ( .A1(n92395), .A2(n92396), .ZN(n92313) );
  NOR4_X1 U77945 ( .A1(n92397), .A2(n92398), .A3(n92399), .A4(n92400), .ZN(
        n92396) );
  NAND2_X1 U77946 ( .A1(n92401), .A2(n92402), .ZN(n92400) );
  AOI22_X1 U77947 ( .A1(n90499), .A2(n108231), .B1(n90500), .B2(n108230), .ZN(
        n92402) );
  AOI22_X1 U77948 ( .A1(n90501), .A2(n70820), .B1(n90502), .B2(n108228), .ZN(
        n92401) );
  NAND2_X1 U77949 ( .A1(n92403), .A2(n92404), .ZN(n92399) );
  AOI22_X1 U77950 ( .A1(n90505), .A2(n108226), .B1(n90506), .B2(n108229), .ZN(
        n92404) );
  AOI22_X1 U77951 ( .A1(n105651), .A2(n70826), .B1(n90508), .B2(n108227), .ZN(
        n92403) );
  NAND2_X1 U77952 ( .A1(n92405), .A2(n92406), .ZN(n92398) );
  AOI22_X1 U77953 ( .A1(n105650), .A2(n108237), .B1(n105649), .B2(n70832), 
        .ZN(n92406) );
  AOI22_X1 U77954 ( .A1(n105648), .A2(n108235), .B1(n105647), .B2(n108236), 
        .ZN(n92405) );
  NAND2_X1 U77955 ( .A1(n92407), .A2(n92408), .ZN(n92397) );
  AOI22_X1 U77956 ( .A1(n90517), .A2(n108232), .B1(n105646), .B2(n108234), 
        .ZN(n92408) );
  AOI22_X1 U77957 ( .A1(n105645), .A2(n108238), .B1(n90520), .B2(n108233), 
        .ZN(n92407) );
  NOR4_X1 U77958 ( .A1(n92409), .A2(n92410), .A3(n92411), .A4(n92412), .ZN(
        n92395) );
  NAND2_X1 U77959 ( .A1(n92413), .A2(n92414), .ZN(n92412) );
  AOI22_X1 U77960 ( .A1(n90527), .A2(n108212), .B1(n90528), .B2(n108216), .ZN(
        n92414) );
  AOI22_X1 U77961 ( .A1(n90529), .A2(n108215), .B1(n90530), .B2(n70803), .ZN(
        n92413) );
  NAND2_X1 U77962 ( .A1(n92415), .A2(n92416), .ZN(n92411) );
  AOI22_X1 U77963 ( .A1(n90533), .A2(n108222), .B1(n90534), .B2(n108211), .ZN(
        n92416) );
  AOI22_X1 U77964 ( .A1(n90535), .A2(n108214), .B1(n90536), .B2(n108219), .ZN(
        n92415) );
  NAND2_X1 U77965 ( .A1(n92417), .A2(n92418), .ZN(n92410) );
  AOI22_X1 U77966 ( .A1(n90539), .A2(n108218), .B1(n90540), .B2(n108223), .ZN(
        n92418) );
  AOI22_X1 U77967 ( .A1(n90541), .A2(n108225), .B1(n90542), .B2(n108221), .ZN(
        n92417) );
  NAND2_X1 U77968 ( .A1(n92419), .A2(n92420), .ZN(n92409) );
  AOI22_X1 U77969 ( .A1(n90545), .A2(n70821), .B1(n90546), .B2(n108217), .ZN(
        n92420) );
  AOI22_X1 U77970 ( .A1(n90547), .A2(n108220), .B1(n90548), .B2(n108224), .ZN(
        n92419) );
  AOI21_X1 U77971 ( .B1(n90295), .B2(n88446), .A(n92422), .ZN(n92421) );
  OAI21_X1 U77972 ( .B1(n92423), .B2(n105659), .A(n92424), .ZN(n92422) );
  OAI21_X1 U77973 ( .B1(n92425), .B2(n92426), .A(n105658), .ZN(n92424) );
  OAI21_X1 U77974 ( .B1(n101908), .B2(n90303), .A(n92427), .ZN(n92426) );
  AOI22_X1 U77975 ( .A1(n105656), .A2(n108382), .B1(n105655), .B2(n71021), 
        .ZN(n92427) );
  NAND2_X1 U77976 ( .A1(n92428), .A2(n92429), .ZN(n92425) );
  AOI22_X1 U77977 ( .A1(n105654), .A2(n108387), .B1(n105653), .B2(n108384), 
        .ZN(n92429) );
  AOI22_X1 U77978 ( .A1(n90311), .A2(n71019), .B1(n105652), .B2(n108383), .ZN(
        n92428) );
  NOR4_X1 U77979 ( .A1(n92430), .A2(n92431), .A3(n92432), .A4(n92433), .ZN(
        n92423) );
  NAND2_X1 U77980 ( .A1(n92434), .A2(n92435), .ZN(n92433) );
  NOR4_X1 U77981 ( .A1(n92436), .A2(n92437), .A3(n92438), .A4(n92439), .ZN(
        n92435) );
  NAND2_X1 U77982 ( .A1(n92440), .A2(n92441), .ZN(n92439) );
  AOI22_X1 U77983 ( .A1(n90325), .A2(n108363), .B1(n90326), .B2(n108364), .ZN(
        n92441) );
  AOI22_X1 U77984 ( .A1(n90327), .A2(n108372), .B1(n90328), .B2(n108370), .ZN(
        n92440) );
  NAND2_X1 U77985 ( .A1(n92442), .A2(n92443), .ZN(n92438) );
  AOI22_X1 U77986 ( .A1(n90331), .A2(n70888), .B1(n90332), .B2(n108367), .ZN(
        n92443) );
  AOI22_X1 U77987 ( .A1(n90333), .A2(n70992), .B1(n90334), .B2(n108283), .ZN(
        n92442) );
  NAND2_X1 U77988 ( .A1(n92444), .A2(n92445), .ZN(n92437) );
  AOI22_X1 U77989 ( .A1(n90337), .A2(n108287), .B1(n90338), .B2(n70892), .ZN(
        n92445) );
  AOI22_X1 U77990 ( .A1(n90339), .A2(n108368), .B1(n90340), .B2(n108365), .ZN(
        n92444) );
  NAND2_X1 U77991 ( .A1(n92446), .A2(n92447), .ZN(n92436) );
  AOI22_X1 U77992 ( .A1(n90343), .A2(n108285), .B1(n90344), .B2(n108289), .ZN(
        n92447) );
  AOI22_X1 U77993 ( .A1(n90345), .A2(n108288), .B1(n90346), .B2(n70894), .ZN(
        n92446) );
  NOR4_X1 U77994 ( .A1(n92448), .A2(n92449), .A3(n92450), .A4(n92451), .ZN(
        n92434) );
  NAND2_X1 U77995 ( .A1(n92452), .A2(n92453), .ZN(n92451) );
  AOI22_X1 U77996 ( .A1(n90353), .A2(n108373), .B1(n90354), .B2(n108376), .ZN(
        n92453) );
  AOI22_X1 U77997 ( .A1(n90355), .A2(n108377), .B1(n90356), .B2(n108379), .ZN(
        n92452) );
  NAND2_X1 U77998 ( .A1(n92454), .A2(n92455), .ZN(n92450) );
  AOI22_X1 U77999 ( .A1(n90359), .A2(n108378), .B1(n90360), .B2(n108374), .ZN(
        n92455) );
  AOI22_X1 U78000 ( .A1(n90361), .A2(n108380), .B1(n90362), .B2(n108375), .ZN(
        n92454) );
  NAND2_X1 U78001 ( .A1(n92456), .A2(n92457), .ZN(n92449) );
  AOI22_X1 U78002 ( .A1(n90365), .A2(n71002), .B1(n90366), .B2(n71001), .ZN(
        n92457) );
  AOI22_X1 U78003 ( .A1(n90367), .A2(n71004), .B1(n90368), .B2(n108381), .ZN(
        n92456) );
  NAND2_X1 U78004 ( .A1(n92458), .A2(n92459), .ZN(n92448) );
  AOI22_X1 U78005 ( .A1(n90371), .A2(n108366), .B1(n90372), .B2(n108371), .ZN(
        n92459) );
  AOI22_X1 U78006 ( .A1(n90373), .A2(n70999), .B1(n90374), .B2(n108369), .ZN(
        n92458) );
  NAND2_X1 U78007 ( .A1(n92460), .A2(n92461), .ZN(n92432) );
  NOR4_X1 U78008 ( .A1(n92462), .A2(n92463), .A3(n92464), .A4(n92465), .ZN(
        n92461) );
  NAND2_X1 U78009 ( .A1(n92466), .A2(n92467), .ZN(n92465) );
  AOI22_X1 U78010 ( .A1(n90383), .A2(n108298), .B1(n90384), .B2(n108300), .ZN(
        n92467) );
  AOI22_X1 U78011 ( .A1(n90385), .A2(n70917), .B1(n90386), .B2(n108299), .ZN(
        n92466) );
  NAND2_X1 U78012 ( .A1(n92468), .A2(n92469), .ZN(n92464) );
  AOI22_X1 U78013 ( .A1(n90389), .A2(n70921), .B1(n90390), .B2(n70923), .ZN(
        n92469) );
  AOI22_X1 U78014 ( .A1(n90391), .A2(n108306), .B1(n90392), .B2(n108307), .ZN(
        n92468) );
  NAND2_X1 U78015 ( .A1(n92470), .A2(n92471), .ZN(n92463) );
  AOI22_X1 U78016 ( .A1(n90395), .A2(n108303), .B1(n90396), .B2(n108305), .ZN(
        n92471) );
  AOI22_X1 U78017 ( .A1(n90397), .A2(n108308), .B1(n90398), .B2(n108304), .ZN(
        n92470) );
  NAND2_X1 U78018 ( .A1(n92472), .A2(n92473), .ZN(n92462) );
  AOI22_X1 U78019 ( .A1(n90401), .A2(n108313), .B1(n90402), .B2(n70928), .ZN(
        n92473) );
  AOI22_X1 U78020 ( .A1(n90403), .A2(n108312), .B1(n90404), .B2(n70926), .ZN(
        n92472) );
  NOR4_X1 U78021 ( .A1(n92474), .A2(n92475), .A3(n92476), .A4(n92477), .ZN(
        n92460) );
  NAND2_X1 U78022 ( .A1(n92478), .A2(n92479), .ZN(n92477) );
  AOI22_X1 U78023 ( .A1(n90411), .A2(n108293), .B1(n90412), .B2(n108284), .ZN(
        n92479) );
  AOI22_X1 U78024 ( .A1(n90413), .A2(n108286), .B1(n90414), .B2(n70900), .ZN(
        n92478) );
  NAND2_X1 U78025 ( .A1(n92480), .A2(n92481), .ZN(n92476) );
  AOI22_X1 U78026 ( .A1(n90417), .A2(n108291), .B1(n90418), .B2(n108295), .ZN(
        n92481) );
  AOI22_X1 U78027 ( .A1(n90419), .A2(n108297), .B1(n90420), .B2(n108294), .ZN(
        n92480) );
  NAND2_X1 U78028 ( .A1(n92482), .A2(n92483), .ZN(n92475) );
  AOI22_X1 U78029 ( .A1(n90423), .A2(n70909), .B1(n90424), .B2(n108290), .ZN(
        n92483) );
  AOI22_X1 U78030 ( .A1(n90425), .A2(n108292), .B1(n90426), .B2(n108296), .ZN(
        n92482) );
  NAND2_X1 U78031 ( .A1(n92484), .A2(n92485), .ZN(n92474) );
  AOI22_X1 U78032 ( .A1(n90429), .A2(n108302), .B1(n90430), .B2(n70913), .ZN(
        n92485) );
  AOI22_X1 U78033 ( .A1(n90431), .A2(n70911), .B1(n90432), .B2(n108301), .ZN(
        n92484) );
  NAND2_X1 U78034 ( .A1(n92486), .A2(n92487), .ZN(n92431) );
  NOR4_X1 U78035 ( .A1(n92488), .A2(n92489), .A3(n92490), .A4(n92491), .ZN(
        n92487) );
  NAND2_X1 U78036 ( .A1(n92492), .A2(n92493), .ZN(n92491) );
  AOI22_X1 U78037 ( .A1(n90441), .A2(n70951), .B1(n90442), .B2(n108323), .ZN(
        n92493) );
  AOI22_X1 U78038 ( .A1(n90443), .A2(n108327), .B1(n90444), .B2(n108326), .ZN(
        n92492) );
  NAND2_X1 U78039 ( .A1(n92494), .A2(n92495), .ZN(n92490) );
  AOI22_X1 U78040 ( .A1(n90447), .A2(n108332), .B1(n90448), .B2(n108331), .ZN(
        n92495) );
  AOI22_X1 U78041 ( .A1(n90449), .A2(n108322), .B1(n90450), .B2(n108324), .ZN(
        n92494) );
  NAND2_X1 U78042 ( .A1(n92496), .A2(n92497), .ZN(n92489) );
  AOI22_X1 U78043 ( .A1(n90453), .A2(n108333), .B1(n90454), .B2(n108329), .ZN(
        n92497) );
  AOI22_X1 U78044 ( .A1(n90455), .A2(n70955), .B1(n90456), .B2(n70957), .ZN(
        n92496) );
  NAND2_X1 U78045 ( .A1(n92498), .A2(n92499), .ZN(n92488) );
  AOI22_X1 U78046 ( .A1(n90459), .A2(n108336), .B1(n90460), .B2(n70963), .ZN(
        n92499) );
  AOI22_X1 U78047 ( .A1(n90461), .A2(n108328), .B1(n90462), .B2(n108330), .ZN(
        n92498) );
  NOR4_X1 U78048 ( .A1(n92500), .A2(n92501), .A3(n92502), .A4(n92503), .ZN(
        n92486) );
  NAND2_X1 U78049 ( .A1(n92504), .A2(n92505), .ZN(n92503) );
  AOI22_X1 U78050 ( .A1(n90469), .A2(n108311), .B1(n90470), .B2(n108316), .ZN(
        n92505) );
  AOI22_X1 U78051 ( .A1(n90471), .A2(n108310), .B1(n90472), .B2(n70931), .ZN(
        n92504) );
  NAND2_X1 U78052 ( .A1(n92506), .A2(n92507), .ZN(n92502) );
  AOI22_X1 U78053 ( .A1(n90475), .A2(n70940), .B1(n90476), .B2(n108318), .ZN(
        n92507) );
  AOI22_X1 U78054 ( .A1(n90477), .A2(n108319), .B1(n90478), .B2(n108309), .ZN(
        n92506) );
  NAND2_X1 U78055 ( .A1(n92508), .A2(n92509), .ZN(n92501) );
  AOI22_X1 U78056 ( .A1(n90481), .A2(n108317), .B1(n90482), .B2(n108321), .ZN(
        n92509) );
  AOI22_X1 U78057 ( .A1(n90483), .A2(n108315), .B1(n90484), .B2(n108320), .ZN(
        n92508) );
  NAND2_X1 U78058 ( .A1(n92510), .A2(n92511), .ZN(n92500) );
  AOI22_X1 U78059 ( .A1(n90487), .A2(n70945), .B1(n90488), .B2(n108325), .ZN(
        n92511) );
  AOI22_X1 U78060 ( .A1(n90489), .A2(n70943), .B1(n90490), .B2(n108314), .ZN(
        n92510) );
  NAND2_X1 U78061 ( .A1(n92512), .A2(n92513), .ZN(n92430) );
  NOR4_X1 U78062 ( .A1(n92514), .A2(n92515), .A3(n92516), .A4(n92517), .ZN(
        n92513) );
  NAND2_X1 U78063 ( .A1(n92518), .A2(n92519), .ZN(n92517) );
  AOI22_X1 U78064 ( .A1(n90499), .A2(n108354), .B1(n90500), .B2(n108353), .ZN(
        n92519) );
  AOI22_X1 U78065 ( .A1(n90501), .A2(n70979), .B1(n90502), .B2(n108351), .ZN(
        n92518) );
  NAND2_X1 U78066 ( .A1(n92520), .A2(n92521), .ZN(n92516) );
  AOI22_X1 U78067 ( .A1(n90505), .A2(n108349), .B1(n90506), .B2(n108352), .ZN(
        n92521) );
  AOI22_X1 U78068 ( .A1(n105651), .A2(n70985), .B1(n90508), .B2(n108350), .ZN(
        n92520) );
  NAND2_X1 U78069 ( .A1(n92522), .A2(n92523), .ZN(n92515) );
  AOI22_X1 U78070 ( .A1(n105650), .A2(n108360), .B1(n105649), .B2(n70991), 
        .ZN(n92523) );
  AOI22_X1 U78071 ( .A1(n105648), .A2(n108358), .B1(n105647), .B2(n108359), 
        .ZN(n92522) );
  NAND2_X1 U78072 ( .A1(n92524), .A2(n92525), .ZN(n92514) );
  AOI22_X1 U78073 ( .A1(n90517), .A2(n108355), .B1(n105646), .B2(n108357), 
        .ZN(n92525) );
  AOI22_X1 U78074 ( .A1(n105645), .A2(n108361), .B1(n105644), .B2(n108356), 
        .ZN(n92524) );
  NOR4_X1 U78075 ( .A1(n92526), .A2(n92527), .A3(n92528), .A4(n92529), .ZN(
        n92512) );
  NAND2_X1 U78076 ( .A1(n92530), .A2(n92531), .ZN(n92529) );
  AOI22_X1 U78077 ( .A1(n90527), .A2(n108335), .B1(n90528), .B2(n108339), .ZN(
        n92531) );
  AOI22_X1 U78078 ( .A1(n90529), .A2(n108338), .B1(n90530), .B2(n70962), .ZN(
        n92530) );
  NAND2_X1 U78079 ( .A1(n92532), .A2(n92533), .ZN(n92528) );
  AOI22_X1 U78080 ( .A1(n90533), .A2(n108345), .B1(n90534), .B2(n108334), .ZN(
        n92533) );
  AOI22_X1 U78081 ( .A1(n90535), .A2(n108337), .B1(n90536), .B2(n108342), .ZN(
        n92532) );
  NAND2_X1 U78082 ( .A1(n92534), .A2(n92535), .ZN(n92527) );
  AOI22_X1 U78083 ( .A1(n90539), .A2(n108341), .B1(n90540), .B2(n108346), .ZN(
        n92535) );
  AOI22_X1 U78084 ( .A1(n90541), .A2(n108348), .B1(n90542), .B2(n108344), .ZN(
        n92534) );
  NAND2_X1 U78085 ( .A1(n92536), .A2(n92537), .ZN(n92526) );
  AOI22_X1 U78086 ( .A1(n90545), .A2(n70980), .B1(n90546), .B2(n108340), .ZN(
        n92537) );
  AOI22_X1 U78087 ( .A1(n90547), .A2(n108343), .B1(n90548), .B2(n108347), .ZN(
        n92536) );
  AOI21_X1 U78088 ( .B1(n90295), .B2(n88564), .A(n92539), .ZN(n92538) );
  OAI21_X1 U78089 ( .B1(n92540), .B2(n90298), .A(n92541), .ZN(n92539) );
  OAI21_X1 U78090 ( .B1(n92542), .B2(n92543), .A(n105658), .ZN(n92541) );
  OAI21_X1 U78091 ( .B1(n101892), .B2(n105657), .A(n92544), .ZN(n92543) );
  AOI22_X1 U78092 ( .A1(n105656), .A2(n108493), .B1(n105655), .B2(n71166), 
        .ZN(n92544) );
  NAND2_X1 U78093 ( .A1(n92545), .A2(n92546), .ZN(n92542) );
  AOI22_X1 U78094 ( .A1(n105654), .A2(n108498), .B1(n105653), .B2(n108495), 
        .ZN(n92546) );
  AOI22_X1 U78095 ( .A1(n90311), .A2(n71164), .B1(n105652), .B2(n108494), .ZN(
        n92545) );
  NOR4_X1 U78096 ( .A1(n92547), .A2(n92548), .A3(n92549), .A4(n92550), .ZN(
        n92540) );
  NAND2_X1 U78097 ( .A1(n92551), .A2(n92552), .ZN(n92550) );
  NOR4_X1 U78098 ( .A1(n92553), .A2(n92554), .A3(n92555), .A4(n92556), .ZN(
        n92552) );
  NAND2_X1 U78099 ( .A1(n92557), .A2(n92558), .ZN(n92556) );
  AOI22_X1 U78100 ( .A1(n90325), .A2(n108474), .B1(n90326), .B2(n108475), .ZN(
        n92558) );
  AOI22_X1 U78101 ( .A1(n90327), .A2(n108483), .B1(n90328), .B2(n108481), .ZN(
        n92557) );
  NAND2_X1 U78102 ( .A1(n92559), .A2(n92560), .ZN(n92555) );
  AOI22_X1 U78103 ( .A1(n90331), .A2(n71033), .B1(n90332), .B2(n108478), .ZN(
        n92560) );
  AOI22_X1 U78104 ( .A1(n90333), .A2(n71137), .B1(n90334), .B2(n108394), .ZN(
        n92559) );
  NAND2_X1 U78105 ( .A1(n92561), .A2(n92562), .ZN(n92554) );
  AOI22_X1 U78106 ( .A1(n90337), .A2(n108398), .B1(n90338), .B2(n71037), .ZN(
        n92562) );
  AOI22_X1 U78107 ( .A1(n90339), .A2(n108479), .B1(n90340), .B2(n108476), .ZN(
        n92561) );
  NAND2_X1 U78108 ( .A1(n92563), .A2(n92564), .ZN(n92553) );
  AOI22_X1 U78109 ( .A1(n90343), .A2(n108396), .B1(n90344), .B2(n108400), .ZN(
        n92564) );
  AOI22_X1 U78110 ( .A1(n90345), .A2(n108399), .B1(n90346), .B2(n71039), .ZN(
        n92563) );
  NOR4_X1 U78111 ( .A1(n92565), .A2(n92566), .A3(n92567), .A4(n92568), .ZN(
        n92551) );
  NAND2_X1 U78112 ( .A1(n92569), .A2(n92570), .ZN(n92568) );
  AOI22_X1 U78113 ( .A1(n90353), .A2(n108484), .B1(n90354), .B2(n108487), .ZN(
        n92570) );
  AOI22_X1 U78114 ( .A1(n90355), .A2(n108488), .B1(n90356), .B2(n108490), .ZN(
        n92569) );
  NAND2_X1 U78115 ( .A1(n92571), .A2(n92572), .ZN(n92567) );
  AOI22_X1 U78116 ( .A1(n90359), .A2(n108489), .B1(n90360), .B2(n108485), .ZN(
        n92572) );
  AOI22_X1 U78117 ( .A1(n90361), .A2(n108491), .B1(n90362), .B2(n108486), .ZN(
        n92571) );
  NAND2_X1 U78118 ( .A1(n92573), .A2(n92574), .ZN(n92566) );
  AOI22_X1 U78119 ( .A1(n90365), .A2(n71147), .B1(n90366), .B2(n71146), .ZN(
        n92574) );
  AOI22_X1 U78120 ( .A1(n90367), .A2(n71149), .B1(n90368), .B2(n108492), .ZN(
        n92573) );
  NAND2_X1 U78121 ( .A1(n92575), .A2(n92576), .ZN(n92565) );
  AOI22_X1 U78122 ( .A1(n90371), .A2(n108477), .B1(n90372), .B2(n108482), .ZN(
        n92576) );
  AOI22_X1 U78123 ( .A1(n90373), .A2(n71144), .B1(n90374), .B2(n108480), .ZN(
        n92575) );
  NAND2_X1 U78124 ( .A1(n92577), .A2(n92578), .ZN(n92549) );
  NOR4_X1 U78125 ( .A1(n92579), .A2(n92580), .A3(n92581), .A4(n92582), .ZN(
        n92578) );
  NAND2_X1 U78126 ( .A1(n92583), .A2(n92584), .ZN(n92582) );
  AOI22_X1 U78127 ( .A1(n90383), .A2(n108409), .B1(n90384), .B2(n108411), .ZN(
        n92584) );
  AOI22_X1 U78128 ( .A1(n90385), .A2(n71062), .B1(n90386), .B2(n108410), .ZN(
        n92583) );
  NAND2_X1 U78129 ( .A1(n92585), .A2(n92586), .ZN(n92581) );
  AOI22_X1 U78130 ( .A1(n90389), .A2(n71066), .B1(n90390), .B2(n71068), .ZN(
        n92586) );
  AOI22_X1 U78131 ( .A1(n90391), .A2(n108417), .B1(n90392), .B2(n108418), .ZN(
        n92585) );
  NAND2_X1 U78132 ( .A1(n92587), .A2(n92588), .ZN(n92580) );
  AOI22_X1 U78133 ( .A1(n90395), .A2(n108414), .B1(n90396), .B2(n108416), .ZN(
        n92588) );
  AOI22_X1 U78134 ( .A1(n90397), .A2(n108419), .B1(n90398), .B2(n108415), .ZN(
        n92587) );
  NAND2_X1 U78135 ( .A1(n92589), .A2(n92590), .ZN(n92579) );
  AOI22_X1 U78136 ( .A1(n90401), .A2(n108424), .B1(n90402), .B2(n71073), .ZN(
        n92590) );
  AOI22_X1 U78137 ( .A1(n90403), .A2(n108423), .B1(n90404), .B2(n71071), .ZN(
        n92589) );
  NOR4_X1 U78138 ( .A1(n92591), .A2(n92592), .A3(n92593), .A4(n92594), .ZN(
        n92577) );
  NAND2_X1 U78139 ( .A1(n92595), .A2(n92596), .ZN(n92594) );
  AOI22_X1 U78140 ( .A1(n90411), .A2(n108404), .B1(n90412), .B2(n108395), .ZN(
        n92596) );
  AOI22_X1 U78141 ( .A1(n90413), .A2(n108397), .B1(n90414), .B2(n71045), .ZN(
        n92595) );
  NAND2_X1 U78142 ( .A1(n92597), .A2(n92598), .ZN(n92593) );
  AOI22_X1 U78143 ( .A1(n90417), .A2(n108402), .B1(n90418), .B2(n108406), .ZN(
        n92598) );
  AOI22_X1 U78144 ( .A1(n90419), .A2(n108408), .B1(n90420), .B2(n108405), .ZN(
        n92597) );
  NAND2_X1 U78145 ( .A1(n92599), .A2(n92600), .ZN(n92592) );
  AOI22_X1 U78146 ( .A1(n90423), .A2(n71054), .B1(n90424), .B2(n108401), .ZN(
        n92600) );
  AOI22_X1 U78147 ( .A1(n90425), .A2(n108403), .B1(n90426), .B2(n108407), .ZN(
        n92599) );
  NAND2_X1 U78148 ( .A1(n92601), .A2(n92602), .ZN(n92591) );
  AOI22_X1 U78149 ( .A1(n90429), .A2(n108413), .B1(n90430), .B2(n71058), .ZN(
        n92602) );
  AOI22_X1 U78150 ( .A1(n90431), .A2(n71056), .B1(n90432), .B2(n108412), .ZN(
        n92601) );
  NAND2_X1 U78151 ( .A1(n92603), .A2(n92604), .ZN(n92548) );
  NOR4_X1 U78152 ( .A1(n92605), .A2(n92606), .A3(n92607), .A4(n92608), .ZN(
        n92604) );
  NAND2_X1 U78153 ( .A1(n92609), .A2(n92610), .ZN(n92608) );
  AOI22_X1 U78154 ( .A1(n90441), .A2(n71096), .B1(n90442), .B2(n108434), .ZN(
        n92610) );
  AOI22_X1 U78155 ( .A1(n90443), .A2(n108438), .B1(n90444), .B2(n108437), .ZN(
        n92609) );
  NAND2_X1 U78156 ( .A1(n92611), .A2(n92612), .ZN(n92607) );
  AOI22_X1 U78157 ( .A1(n90447), .A2(n108443), .B1(n90448), .B2(n108442), .ZN(
        n92612) );
  AOI22_X1 U78158 ( .A1(n90449), .A2(n108433), .B1(n90450), .B2(n108435), .ZN(
        n92611) );
  NAND2_X1 U78159 ( .A1(n92613), .A2(n92614), .ZN(n92606) );
  AOI22_X1 U78160 ( .A1(n90453), .A2(n108444), .B1(n90454), .B2(n108440), .ZN(
        n92614) );
  AOI22_X1 U78161 ( .A1(n90455), .A2(n71100), .B1(n90456), .B2(n71102), .ZN(
        n92613) );
  NAND2_X1 U78162 ( .A1(n92615), .A2(n92616), .ZN(n92605) );
  AOI22_X1 U78163 ( .A1(n90459), .A2(n108447), .B1(n90460), .B2(n71108), .ZN(
        n92616) );
  AOI22_X1 U78164 ( .A1(n90461), .A2(n108439), .B1(n90462), .B2(n108441), .ZN(
        n92615) );
  NOR4_X1 U78165 ( .A1(n92617), .A2(n92618), .A3(n92619), .A4(n92620), .ZN(
        n92603) );
  NAND2_X1 U78166 ( .A1(n92621), .A2(n92622), .ZN(n92620) );
  AOI22_X1 U78167 ( .A1(n90469), .A2(n108422), .B1(n90470), .B2(n108427), .ZN(
        n92622) );
  AOI22_X1 U78168 ( .A1(n90471), .A2(n108421), .B1(n90472), .B2(n71076), .ZN(
        n92621) );
  NAND2_X1 U78169 ( .A1(n92623), .A2(n92624), .ZN(n92619) );
  AOI22_X1 U78170 ( .A1(n90475), .A2(n71085), .B1(n90476), .B2(n108429), .ZN(
        n92624) );
  AOI22_X1 U78171 ( .A1(n90477), .A2(n108430), .B1(n90478), .B2(n108420), .ZN(
        n92623) );
  NAND2_X1 U78172 ( .A1(n92625), .A2(n92626), .ZN(n92618) );
  AOI22_X1 U78173 ( .A1(n90481), .A2(n108428), .B1(n90482), .B2(n108432), .ZN(
        n92626) );
  AOI22_X1 U78174 ( .A1(n90483), .A2(n108426), .B1(n90484), .B2(n108431), .ZN(
        n92625) );
  NAND2_X1 U78175 ( .A1(n92627), .A2(n92628), .ZN(n92617) );
  AOI22_X1 U78176 ( .A1(n90487), .A2(n71090), .B1(n90488), .B2(n108436), .ZN(
        n92628) );
  AOI22_X1 U78177 ( .A1(n90489), .A2(n71088), .B1(n90490), .B2(n108425), .ZN(
        n92627) );
  NAND2_X1 U78178 ( .A1(n92629), .A2(n92630), .ZN(n92547) );
  NOR4_X1 U78179 ( .A1(n92631), .A2(n92632), .A3(n92633), .A4(n92634), .ZN(
        n92630) );
  NAND2_X1 U78180 ( .A1(n92635), .A2(n92636), .ZN(n92634) );
  AOI22_X1 U78181 ( .A1(n90499), .A2(n108465), .B1(n90500), .B2(n108464), .ZN(
        n92636) );
  AOI22_X1 U78182 ( .A1(n90501), .A2(n71124), .B1(n90502), .B2(n108462), .ZN(
        n92635) );
  NAND2_X1 U78183 ( .A1(n92637), .A2(n92638), .ZN(n92633) );
  AOI22_X1 U78184 ( .A1(n90505), .A2(n108460), .B1(n90506), .B2(n108463), .ZN(
        n92638) );
  AOI22_X1 U78185 ( .A1(n105651), .A2(n71130), .B1(n90508), .B2(n108461), .ZN(
        n92637) );
  NAND2_X1 U78186 ( .A1(n92639), .A2(n92640), .ZN(n92632) );
  AOI22_X1 U78187 ( .A1(n105650), .A2(n108471), .B1(n105649), .B2(n71136), 
        .ZN(n92640) );
  AOI22_X1 U78188 ( .A1(n105648), .A2(n108469), .B1(n105647), .B2(n108470), 
        .ZN(n92639) );
  NAND2_X1 U78189 ( .A1(n92641), .A2(n92642), .ZN(n92631) );
  AOI22_X1 U78190 ( .A1(n90517), .A2(n108466), .B1(n105646), .B2(n108468), 
        .ZN(n92642) );
  AOI22_X1 U78191 ( .A1(n105645), .A2(n108472), .B1(n90520), .B2(n108467), 
        .ZN(n92641) );
  NOR4_X1 U78192 ( .A1(n92643), .A2(n92644), .A3(n92645), .A4(n92646), .ZN(
        n92629) );
  NAND2_X1 U78193 ( .A1(n92647), .A2(n92648), .ZN(n92646) );
  AOI22_X1 U78194 ( .A1(n90527), .A2(n108446), .B1(n90528), .B2(n108450), .ZN(
        n92648) );
  AOI22_X1 U78195 ( .A1(n90529), .A2(n108449), .B1(n90530), .B2(n71107), .ZN(
        n92647) );
  NAND2_X1 U78196 ( .A1(n92649), .A2(n92650), .ZN(n92645) );
  AOI22_X1 U78197 ( .A1(n90533), .A2(n108456), .B1(n90534), .B2(n108445), .ZN(
        n92650) );
  AOI22_X1 U78198 ( .A1(n90535), .A2(n108448), .B1(n90536), .B2(n108453), .ZN(
        n92649) );
  NAND2_X1 U78199 ( .A1(n92651), .A2(n92652), .ZN(n92644) );
  AOI22_X1 U78200 ( .A1(n90539), .A2(n108452), .B1(n90540), .B2(n108457), .ZN(
        n92652) );
  AOI22_X1 U78201 ( .A1(n90541), .A2(n108459), .B1(n90542), .B2(n108455), .ZN(
        n92651) );
  NAND2_X1 U78202 ( .A1(n92653), .A2(n92654), .ZN(n92643) );
  AOI22_X1 U78203 ( .A1(n90545), .A2(n71125), .B1(n90546), .B2(n108451), .ZN(
        n92654) );
  AOI22_X1 U78204 ( .A1(n90547), .A2(n108454), .B1(n90548), .B2(n108458), .ZN(
        n92653) );
  AOI21_X1 U78205 ( .B1(n90295), .B2(n88682), .A(n92656), .ZN(n92655) );
  OAI21_X1 U78206 ( .B1(n92657), .B2(n90298), .A(n92658), .ZN(n92656) );
  OAI21_X1 U78207 ( .B1(n92659), .B2(n92660), .A(n105658), .ZN(n92658) );
  OAI21_X1 U78208 ( .B1(n101876), .B2(n90303), .A(n92661), .ZN(n92660) );
  AOI22_X1 U78209 ( .A1(n105656), .A2(n107730), .B1(n105655), .B2(n70127), 
        .ZN(n92661) );
  NAND2_X1 U78210 ( .A1(n92662), .A2(n92663), .ZN(n92659) );
  AOI22_X1 U78211 ( .A1(n105654), .A2(n107735), .B1(n105653), .B2(n107732), 
        .ZN(n92663) );
  AOI22_X1 U78212 ( .A1(n90311), .A2(n70125), .B1(n105652), .B2(n107731), .ZN(
        n92662) );
  NOR4_X1 U78213 ( .A1(n92664), .A2(n92665), .A3(n92666), .A4(n92667), .ZN(
        n92657) );
  NAND2_X1 U78214 ( .A1(n92668), .A2(n92669), .ZN(n92667) );
  NOR4_X1 U78215 ( .A1(n92670), .A2(n92671), .A3(n92672), .A4(n92673), .ZN(
        n92669) );
  NAND2_X1 U78216 ( .A1(n92674), .A2(n92675), .ZN(n92673) );
  AOI22_X1 U78217 ( .A1(n90325), .A2(n107711), .B1(n90326), .B2(n107712), .ZN(
        n92675) );
  AOI22_X1 U78218 ( .A1(n90327), .A2(n107720), .B1(n90328), .B2(n107718), .ZN(
        n92674) );
  NAND2_X1 U78219 ( .A1(n92676), .A2(n92677), .ZN(n92672) );
  AOI22_X1 U78220 ( .A1(n90331), .A2(n69994), .B1(n90332), .B2(n107715), .ZN(
        n92677) );
  AOI22_X1 U78221 ( .A1(n90333), .A2(n70098), .B1(n90334), .B2(n107632), .ZN(
        n92676) );
  NAND2_X1 U78222 ( .A1(n92678), .A2(n92679), .ZN(n92671) );
  AOI22_X1 U78223 ( .A1(n90337), .A2(n107636), .B1(n90338), .B2(n69998), .ZN(
        n92679) );
  AOI22_X1 U78224 ( .A1(n90339), .A2(n107716), .B1(n90340), .B2(n107713), .ZN(
        n92678) );
  NAND2_X1 U78225 ( .A1(n92680), .A2(n92681), .ZN(n92670) );
  AOI22_X1 U78226 ( .A1(n90343), .A2(n107634), .B1(n90344), .B2(n107638), .ZN(
        n92681) );
  AOI22_X1 U78227 ( .A1(n90345), .A2(n107637), .B1(n90346), .B2(n70000), .ZN(
        n92680) );
  NOR4_X1 U78228 ( .A1(n92682), .A2(n92683), .A3(n92684), .A4(n92685), .ZN(
        n92668) );
  NAND2_X1 U78229 ( .A1(n92686), .A2(n92687), .ZN(n92685) );
  AOI22_X1 U78230 ( .A1(n90353), .A2(n107721), .B1(n90354), .B2(n107724), .ZN(
        n92687) );
  AOI22_X1 U78231 ( .A1(n90355), .A2(n107725), .B1(n90356), .B2(n107727), .ZN(
        n92686) );
  NAND2_X1 U78232 ( .A1(n92688), .A2(n92689), .ZN(n92684) );
  AOI22_X1 U78233 ( .A1(n90359), .A2(n107726), .B1(n90360), .B2(n107722), .ZN(
        n92689) );
  AOI22_X1 U78234 ( .A1(n90361), .A2(n107728), .B1(n90362), .B2(n107723), .ZN(
        n92688) );
  NAND2_X1 U78235 ( .A1(n92690), .A2(n92691), .ZN(n92683) );
  AOI22_X1 U78236 ( .A1(n90365), .A2(n70108), .B1(n90366), .B2(n70107), .ZN(
        n92691) );
  AOI22_X1 U78237 ( .A1(n90367), .A2(n70110), .B1(n90368), .B2(n107729), .ZN(
        n92690) );
  NAND2_X1 U78238 ( .A1(n92692), .A2(n92693), .ZN(n92682) );
  AOI22_X1 U78239 ( .A1(n90371), .A2(n107714), .B1(n90372), .B2(n107719), .ZN(
        n92693) );
  AOI22_X1 U78240 ( .A1(n90373), .A2(n70105), .B1(n90374), .B2(n107717), .ZN(
        n92692) );
  NAND2_X1 U78241 ( .A1(n92694), .A2(n92695), .ZN(n92666) );
  NOR4_X1 U78242 ( .A1(n92696), .A2(n92697), .A3(n92698), .A4(n92699), .ZN(
        n92695) );
  NAND2_X1 U78243 ( .A1(n92700), .A2(n92701), .ZN(n92699) );
  AOI22_X1 U78244 ( .A1(n90383), .A2(n107647), .B1(n90384), .B2(n107649), .ZN(
        n92701) );
  AOI22_X1 U78245 ( .A1(n90385), .A2(n70023), .B1(n90386), .B2(n107648), .ZN(
        n92700) );
  NAND2_X1 U78246 ( .A1(n92702), .A2(n92703), .ZN(n92698) );
  AOI22_X1 U78247 ( .A1(n90389), .A2(n70027), .B1(n90390), .B2(n70029), .ZN(
        n92703) );
  AOI22_X1 U78248 ( .A1(n90391), .A2(n107655), .B1(n90392), .B2(n107656), .ZN(
        n92702) );
  NAND2_X1 U78249 ( .A1(n92704), .A2(n92705), .ZN(n92697) );
  AOI22_X1 U78250 ( .A1(n90395), .A2(n107652), .B1(n90396), .B2(n107654), .ZN(
        n92705) );
  AOI22_X1 U78251 ( .A1(n90397), .A2(n107657), .B1(n90398), .B2(n107653), .ZN(
        n92704) );
  NAND2_X1 U78252 ( .A1(n92706), .A2(n92707), .ZN(n92696) );
  AOI22_X1 U78253 ( .A1(n90401), .A2(n107662), .B1(n90402), .B2(n70034), .ZN(
        n92707) );
  AOI22_X1 U78254 ( .A1(n90403), .A2(n107661), .B1(n90404), .B2(n70032), .ZN(
        n92706) );
  NOR4_X1 U78255 ( .A1(n92708), .A2(n92709), .A3(n92710), .A4(n92711), .ZN(
        n92694) );
  NAND2_X1 U78256 ( .A1(n92712), .A2(n92713), .ZN(n92711) );
  AOI22_X1 U78257 ( .A1(n90411), .A2(n107642), .B1(n90412), .B2(n107633), .ZN(
        n92713) );
  AOI22_X1 U78258 ( .A1(n90413), .A2(n107635), .B1(n90414), .B2(n70006), .ZN(
        n92712) );
  NAND2_X1 U78259 ( .A1(n92714), .A2(n92715), .ZN(n92710) );
  AOI22_X1 U78260 ( .A1(n90417), .A2(n107640), .B1(n90418), .B2(n107644), .ZN(
        n92715) );
  AOI22_X1 U78261 ( .A1(n90419), .A2(n107646), .B1(n90420), .B2(n107643), .ZN(
        n92714) );
  NAND2_X1 U78262 ( .A1(n92716), .A2(n92717), .ZN(n92709) );
  AOI22_X1 U78263 ( .A1(n90423), .A2(n70015), .B1(n90424), .B2(n107639), .ZN(
        n92717) );
  AOI22_X1 U78264 ( .A1(n90425), .A2(n107641), .B1(n90426), .B2(n107645), .ZN(
        n92716) );
  NAND2_X1 U78265 ( .A1(n92718), .A2(n92719), .ZN(n92708) );
  AOI22_X1 U78266 ( .A1(n90429), .A2(n107651), .B1(n90430), .B2(n70019), .ZN(
        n92719) );
  AOI22_X1 U78267 ( .A1(n90431), .A2(n70017), .B1(n90432), .B2(n107650), .ZN(
        n92718) );
  NAND2_X1 U78268 ( .A1(n92720), .A2(n92721), .ZN(n92665) );
  NOR4_X1 U78269 ( .A1(n92722), .A2(n92723), .A3(n92724), .A4(n92725), .ZN(
        n92721) );
  NAND2_X1 U78270 ( .A1(n92726), .A2(n92727), .ZN(n92725) );
  AOI22_X1 U78271 ( .A1(n90441), .A2(n70057), .B1(n90442), .B2(n107672), .ZN(
        n92727) );
  AOI22_X1 U78272 ( .A1(n90443), .A2(n107676), .B1(n90444), .B2(n107675), .ZN(
        n92726) );
  NAND2_X1 U78273 ( .A1(n92728), .A2(n92729), .ZN(n92724) );
  AOI22_X1 U78274 ( .A1(n90447), .A2(n107681), .B1(n90448), .B2(n107680), .ZN(
        n92729) );
  AOI22_X1 U78275 ( .A1(n90449), .A2(n107671), .B1(n90450), .B2(n107673), .ZN(
        n92728) );
  NAND2_X1 U78276 ( .A1(n92730), .A2(n92731), .ZN(n92723) );
  AOI22_X1 U78277 ( .A1(n90453), .A2(n107682), .B1(n90454), .B2(n107678), .ZN(
        n92731) );
  AOI22_X1 U78278 ( .A1(n90455), .A2(n70061), .B1(n90456), .B2(n70063), .ZN(
        n92730) );
  NAND2_X1 U78279 ( .A1(n92732), .A2(n92733), .ZN(n92722) );
  AOI22_X1 U78280 ( .A1(n90459), .A2(n107685), .B1(n90460), .B2(n70069), .ZN(
        n92733) );
  AOI22_X1 U78281 ( .A1(n90461), .A2(n107677), .B1(n90462), .B2(n107679), .ZN(
        n92732) );
  NOR4_X1 U78282 ( .A1(n92734), .A2(n92735), .A3(n92736), .A4(n92737), .ZN(
        n92720) );
  NAND2_X1 U78283 ( .A1(n92738), .A2(n92739), .ZN(n92737) );
  AOI22_X1 U78284 ( .A1(n90469), .A2(n107660), .B1(n90470), .B2(n107665), .ZN(
        n92739) );
  AOI22_X1 U78285 ( .A1(n90471), .A2(n107659), .B1(n90472), .B2(n70037), .ZN(
        n92738) );
  NAND2_X1 U78286 ( .A1(n92740), .A2(n92741), .ZN(n92736) );
  AOI22_X1 U78287 ( .A1(n90475), .A2(n70046), .B1(n90476), .B2(n107667), .ZN(
        n92741) );
  AOI22_X1 U78288 ( .A1(n90477), .A2(n107668), .B1(n90478), .B2(n107658), .ZN(
        n92740) );
  NAND2_X1 U78289 ( .A1(n92742), .A2(n92743), .ZN(n92735) );
  AOI22_X1 U78290 ( .A1(n90481), .A2(n107666), .B1(n90482), .B2(n107670), .ZN(
        n92743) );
  AOI22_X1 U78291 ( .A1(n90483), .A2(n107664), .B1(n90484), .B2(n107669), .ZN(
        n92742) );
  NAND2_X1 U78292 ( .A1(n92744), .A2(n92745), .ZN(n92734) );
  AOI22_X1 U78293 ( .A1(n90487), .A2(n70051), .B1(n90488), .B2(n107674), .ZN(
        n92745) );
  AOI22_X1 U78294 ( .A1(n90489), .A2(n70049), .B1(n90490), .B2(n107663), .ZN(
        n92744) );
  NAND2_X1 U78295 ( .A1(n92746), .A2(n92747), .ZN(n92664) );
  NOR4_X1 U78296 ( .A1(n92748), .A2(n92749), .A3(n92750), .A4(n92751), .ZN(
        n92747) );
  NAND2_X1 U78297 ( .A1(n92752), .A2(n92753), .ZN(n92751) );
  AOI22_X1 U78298 ( .A1(n90499), .A2(n107703), .B1(n90500), .B2(n107702), .ZN(
        n92753) );
  AOI22_X1 U78299 ( .A1(n90501), .A2(n70085), .B1(n90502), .B2(n107700), .ZN(
        n92752) );
  NAND2_X1 U78300 ( .A1(n92754), .A2(n92755), .ZN(n92750) );
  AOI22_X1 U78301 ( .A1(n90505), .A2(n107698), .B1(n90506), .B2(n107701), .ZN(
        n92755) );
  AOI22_X1 U78302 ( .A1(n105651), .A2(n70091), .B1(n90508), .B2(n107699), .ZN(
        n92754) );
  NAND2_X1 U78303 ( .A1(n92756), .A2(n92757), .ZN(n92749) );
  AOI22_X1 U78304 ( .A1(n105650), .A2(n107709), .B1(n105649), .B2(n70097), 
        .ZN(n92757) );
  AOI22_X1 U78305 ( .A1(n105648), .A2(n107707), .B1(n105647), .B2(n107708), 
        .ZN(n92756) );
  NAND2_X1 U78306 ( .A1(n92758), .A2(n92759), .ZN(n92748) );
  AOI22_X1 U78307 ( .A1(n90517), .A2(n107704), .B1(n105646), .B2(n107706), 
        .ZN(n92759) );
  AOI22_X1 U78308 ( .A1(n105645), .A2(n107710), .B1(n105644), .B2(n107705), 
        .ZN(n92758) );
  NOR4_X1 U78309 ( .A1(n92760), .A2(n92761), .A3(n92762), .A4(n92763), .ZN(
        n92746) );
  NAND2_X1 U78310 ( .A1(n92764), .A2(n92765), .ZN(n92763) );
  AOI22_X1 U78311 ( .A1(n90527), .A2(n107684), .B1(n90528), .B2(n107688), .ZN(
        n92765) );
  AOI22_X1 U78312 ( .A1(n90529), .A2(n107687), .B1(n90530), .B2(n70068), .ZN(
        n92764) );
  NAND2_X1 U78313 ( .A1(n92766), .A2(n92767), .ZN(n92762) );
  AOI22_X1 U78314 ( .A1(n90533), .A2(n107694), .B1(n90534), .B2(n107683), .ZN(
        n92767) );
  AOI22_X1 U78315 ( .A1(n90535), .A2(n107686), .B1(n90536), .B2(n107691), .ZN(
        n92766) );
  NAND2_X1 U78316 ( .A1(n92768), .A2(n92769), .ZN(n92761) );
  AOI22_X1 U78317 ( .A1(n90539), .A2(n107690), .B1(n90540), .B2(n107695), .ZN(
        n92769) );
  AOI22_X1 U78318 ( .A1(n90541), .A2(n107697), .B1(n90542), .B2(n107693), .ZN(
        n92768) );
  NAND2_X1 U78319 ( .A1(n92770), .A2(n92771), .ZN(n92760) );
  AOI22_X1 U78320 ( .A1(n90545), .A2(n70086), .B1(n90546), .B2(n107689), .ZN(
        n92771) );
  AOI22_X1 U78321 ( .A1(n90547), .A2(n107692), .B1(n90548), .B2(n107696), .ZN(
        n92770) );
  AOI21_X1 U78322 ( .B1(n90295), .B2(n88800), .A(n92773), .ZN(n92772) );
  OAI21_X1 U78323 ( .B1(n92774), .B2(n90298), .A(n92775), .ZN(n92773) );
  OAI21_X1 U78324 ( .B1(n92776), .B2(n92777), .A(n105658), .ZN(n92775) );
  OAI21_X1 U78325 ( .B1(n101858), .B2(n105657), .A(n92778), .ZN(n92777) );
  AOI22_X1 U78326 ( .A1(n105656), .A2(n109645), .B1(n105655), .B2(n72656), 
        .ZN(n92778) );
  NAND2_X1 U78327 ( .A1(n92779), .A2(n92780), .ZN(n92776) );
  AOI22_X1 U78328 ( .A1(n105654), .A2(n109650), .B1(n90310), .B2(n109647), 
        .ZN(n92780) );
  AOI22_X1 U78329 ( .A1(n90311), .A2(n72654), .B1(n105652), .B2(n109646), .ZN(
        n92779) );
  NOR4_X1 U78330 ( .A1(n92781), .A2(n92782), .A3(n92783), .A4(n92784), .ZN(
        n92774) );
  NAND2_X1 U78331 ( .A1(n92785), .A2(n92786), .ZN(n92784) );
  NOR4_X1 U78332 ( .A1(n92787), .A2(n92788), .A3(n92789), .A4(n92790), .ZN(
        n92786) );
  NAND2_X1 U78333 ( .A1(n92791), .A2(n92792), .ZN(n92790) );
  AOI22_X1 U78334 ( .A1(n90325), .A2(n109626), .B1(n90326), .B2(n109627), .ZN(
        n92792) );
  AOI22_X1 U78335 ( .A1(n90327), .A2(n109635), .B1(n90328), .B2(n109633), .ZN(
        n92791) );
  NAND2_X1 U78336 ( .A1(n92793), .A2(n92794), .ZN(n92789) );
  AOI22_X1 U78337 ( .A1(n90331), .A2(n72523), .B1(n90332), .B2(n109630), .ZN(
        n92794) );
  AOI22_X1 U78338 ( .A1(n90333), .A2(n72627), .B1(n90334), .B2(n109550), .ZN(
        n92793) );
  NAND2_X1 U78339 ( .A1(n92795), .A2(n92796), .ZN(n92788) );
  AOI22_X1 U78340 ( .A1(n90337), .A2(n109554), .B1(n90338), .B2(n72527), .ZN(
        n92796) );
  AOI22_X1 U78341 ( .A1(n90339), .A2(n109631), .B1(n90340), .B2(n109628), .ZN(
        n92795) );
  NAND2_X1 U78342 ( .A1(n92797), .A2(n92798), .ZN(n92787) );
  AOI22_X1 U78343 ( .A1(n90343), .A2(n109552), .B1(n90344), .B2(n109556), .ZN(
        n92798) );
  AOI22_X1 U78344 ( .A1(n90345), .A2(n109555), .B1(n90346), .B2(n72529), .ZN(
        n92797) );
  NOR4_X1 U78345 ( .A1(n92799), .A2(n92800), .A3(n92801), .A4(n92802), .ZN(
        n92785) );
  NAND2_X1 U78346 ( .A1(n92803), .A2(n92804), .ZN(n92802) );
  AOI22_X1 U78347 ( .A1(n90353), .A2(n109636), .B1(n90354), .B2(n109639), .ZN(
        n92804) );
  AOI22_X1 U78348 ( .A1(n90355), .A2(n109640), .B1(n90356), .B2(n109642), .ZN(
        n92803) );
  NAND2_X1 U78349 ( .A1(n92805), .A2(n92806), .ZN(n92801) );
  AOI22_X1 U78350 ( .A1(n90359), .A2(n109641), .B1(n90360), .B2(n109637), .ZN(
        n92806) );
  AOI22_X1 U78351 ( .A1(n90361), .A2(n109643), .B1(n90362), .B2(n109638), .ZN(
        n92805) );
  NAND2_X1 U78352 ( .A1(n92807), .A2(n92808), .ZN(n92800) );
  AOI22_X1 U78353 ( .A1(n90365), .A2(n72637), .B1(n90366), .B2(n72636), .ZN(
        n92808) );
  AOI22_X1 U78354 ( .A1(n90367), .A2(n72639), .B1(n90368), .B2(n109644), .ZN(
        n92807) );
  NAND2_X1 U78355 ( .A1(n92809), .A2(n92810), .ZN(n92799) );
  AOI22_X1 U78356 ( .A1(n90371), .A2(n109629), .B1(n90372), .B2(n109634), .ZN(
        n92810) );
  AOI22_X1 U78357 ( .A1(n90373), .A2(n72634), .B1(n90374), .B2(n109632), .ZN(
        n92809) );
  NAND2_X1 U78358 ( .A1(n92811), .A2(n92812), .ZN(n92783) );
  NOR4_X1 U78359 ( .A1(n92813), .A2(n92814), .A3(n92815), .A4(n92816), .ZN(
        n92812) );
  NAND2_X1 U78360 ( .A1(n92817), .A2(n92818), .ZN(n92816) );
  AOI22_X1 U78361 ( .A1(n90383), .A2(n109565), .B1(n90384), .B2(n109567), .ZN(
        n92818) );
  AOI22_X1 U78362 ( .A1(n90385), .A2(n72552), .B1(n90386), .B2(n109566), .ZN(
        n92817) );
  NAND2_X1 U78363 ( .A1(n92819), .A2(n92820), .ZN(n92815) );
  AOI22_X1 U78364 ( .A1(n90389), .A2(n72556), .B1(n90390), .B2(n72558), .ZN(
        n92820) );
  AOI22_X1 U78365 ( .A1(n90391), .A2(n109573), .B1(n90392), .B2(n109574), .ZN(
        n92819) );
  NAND2_X1 U78366 ( .A1(n92821), .A2(n92822), .ZN(n92814) );
  AOI22_X1 U78367 ( .A1(n90395), .A2(n109570), .B1(n90396), .B2(n109572), .ZN(
        n92822) );
  AOI22_X1 U78368 ( .A1(n90397), .A2(n109575), .B1(n90398), .B2(n109571), .ZN(
        n92821) );
  NAND2_X1 U78369 ( .A1(n92823), .A2(n92824), .ZN(n92813) );
  AOI22_X1 U78370 ( .A1(n90401), .A2(n109580), .B1(n90402), .B2(n72563), .ZN(
        n92824) );
  AOI22_X1 U78371 ( .A1(n90403), .A2(n109579), .B1(n90404), .B2(n72561), .ZN(
        n92823) );
  NOR4_X1 U78372 ( .A1(n92825), .A2(n92826), .A3(n92827), .A4(n92828), .ZN(
        n92811) );
  NAND2_X1 U78373 ( .A1(n92829), .A2(n92830), .ZN(n92828) );
  AOI22_X1 U78374 ( .A1(n90411), .A2(n109560), .B1(n90412), .B2(n109551), .ZN(
        n92830) );
  AOI22_X1 U78375 ( .A1(n90413), .A2(n109553), .B1(n90414), .B2(n72535), .ZN(
        n92829) );
  NAND2_X1 U78376 ( .A1(n92831), .A2(n92832), .ZN(n92827) );
  AOI22_X1 U78377 ( .A1(n90417), .A2(n109558), .B1(n90418), .B2(n109562), .ZN(
        n92832) );
  AOI22_X1 U78378 ( .A1(n90419), .A2(n109564), .B1(n90420), .B2(n109561), .ZN(
        n92831) );
  NAND2_X1 U78379 ( .A1(n92833), .A2(n92834), .ZN(n92826) );
  AOI22_X1 U78380 ( .A1(n90423), .A2(n72544), .B1(n90424), .B2(n109557), .ZN(
        n92834) );
  AOI22_X1 U78381 ( .A1(n90425), .A2(n109559), .B1(n90426), .B2(n109563), .ZN(
        n92833) );
  NAND2_X1 U78382 ( .A1(n92835), .A2(n92836), .ZN(n92825) );
  AOI22_X1 U78383 ( .A1(n90429), .A2(n109569), .B1(n90430), .B2(n72548), .ZN(
        n92836) );
  AOI22_X1 U78384 ( .A1(n90431), .A2(n72546), .B1(n90432), .B2(n109568), .ZN(
        n92835) );
  NAND2_X1 U78385 ( .A1(n92837), .A2(n92838), .ZN(n92782) );
  NOR4_X1 U78386 ( .A1(n92839), .A2(n92840), .A3(n92841), .A4(n92842), .ZN(
        n92838) );
  NAND2_X1 U78387 ( .A1(n92843), .A2(n92844), .ZN(n92842) );
  AOI22_X1 U78388 ( .A1(n90441), .A2(n72586), .B1(n90442), .B2(n109590), .ZN(
        n92844) );
  AOI22_X1 U78389 ( .A1(n90443), .A2(n109594), .B1(n90444), .B2(n109593), .ZN(
        n92843) );
  NAND2_X1 U78390 ( .A1(n92845), .A2(n92846), .ZN(n92841) );
  AOI22_X1 U78391 ( .A1(n90447), .A2(n109599), .B1(n90448), .B2(n109598), .ZN(
        n92846) );
  AOI22_X1 U78392 ( .A1(n90449), .A2(n109589), .B1(n90450), .B2(n109591), .ZN(
        n92845) );
  NAND2_X1 U78393 ( .A1(n92847), .A2(n92848), .ZN(n92840) );
  AOI22_X1 U78394 ( .A1(n90453), .A2(n109600), .B1(n90454), .B2(n109596), .ZN(
        n92848) );
  AOI22_X1 U78395 ( .A1(n90455), .A2(n72590), .B1(n90456), .B2(n72592), .ZN(
        n92847) );
  NAND2_X1 U78396 ( .A1(n92849), .A2(n92850), .ZN(n92839) );
  AOI22_X1 U78397 ( .A1(n90459), .A2(n109603), .B1(n90460), .B2(n72598), .ZN(
        n92850) );
  AOI22_X1 U78398 ( .A1(n90461), .A2(n109595), .B1(n90462), .B2(n109597), .ZN(
        n92849) );
  NOR4_X1 U78399 ( .A1(n92851), .A2(n92852), .A3(n92853), .A4(n92854), .ZN(
        n92837) );
  NAND2_X1 U78400 ( .A1(n92855), .A2(n92856), .ZN(n92854) );
  AOI22_X1 U78401 ( .A1(n90469), .A2(n109578), .B1(n90470), .B2(n109583), .ZN(
        n92856) );
  AOI22_X1 U78402 ( .A1(n90471), .A2(n109577), .B1(n90472), .B2(n72566), .ZN(
        n92855) );
  NAND2_X1 U78403 ( .A1(n92857), .A2(n92858), .ZN(n92853) );
  AOI22_X1 U78404 ( .A1(n90475), .A2(n72575), .B1(n90476), .B2(n109585), .ZN(
        n92858) );
  AOI22_X1 U78405 ( .A1(n90477), .A2(n109586), .B1(n90478), .B2(n109576), .ZN(
        n92857) );
  NAND2_X1 U78406 ( .A1(n92859), .A2(n92860), .ZN(n92852) );
  AOI22_X1 U78407 ( .A1(n90481), .A2(n109584), .B1(n90482), .B2(n109588), .ZN(
        n92860) );
  AOI22_X1 U78408 ( .A1(n90483), .A2(n109582), .B1(n90484), .B2(n109587), .ZN(
        n92859) );
  NAND2_X1 U78409 ( .A1(n92861), .A2(n92862), .ZN(n92851) );
  AOI22_X1 U78410 ( .A1(n90487), .A2(n72580), .B1(n90488), .B2(n109592), .ZN(
        n92862) );
  AOI22_X1 U78411 ( .A1(n90489), .A2(n72578), .B1(n90490), .B2(n109581), .ZN(
        n92861) );
  NAND2_X1 U78412 ( .A1(n92863), .A2(n92864), .ZN(n92781) );
  NOR4_X1 U78413 ( .A1(n92865), .A2(n92866), .A3(n92867), .A4(n92868), .ZN(
        n92864) );
  NAND2_X1 U78414 ( .A1(n92869), .A2(n92870), .ZN(n92868) );
  AOI22_X1 U78415 ( .A1(n90499), .A2(n109618), .B1(n90500), .B2(n109617), .ZN(
        n92870) );
  AOI22_X1 U78416 ( .A1(n90501), .A2(n72614), .B1(n90502), .B2(n109615), .ZN(
        n92869) );
  NAND2_X1 U78417 ( .A1(n92871), .A2(n92872), .ZN(n92867) );
  AOI22_X1 U78418 ( .A1(n90505), .A2(n109613), .B1(n90506), .B2(n109616), .ZN(
        n92872) );
  AOI22_X1 U78419 ( .A1(n105651), .A2(n72620), .B1(n90508), .B2(n109614), .ZN(
        n92871) );
  NAND2_X1 U78420 ( .A1(n92873), .A2(n92874), .ZN(n92866) );
  AOI22_X1 U78421 ( .A1(n90511), .A2(n109624), .B1(n105649), .B2(n72626), .ZN(
        n92874) );
  AOI22_X1 U78422 ( .A1(n105648), .A2(n109622), .B1(n105647), .B2(n109623), 
        .ZN(n92873) );
  NAND2_X1 U78423 ( .A1(n92875), .A2(n92876), .ZN(n92865) );
  AOI22_X1 U78424 ( .A1(n90517), .A2(n109619), .B1(n105646), .B2(n109621), 
        .ZN(n92876) );
  AOI22_X1 U78425 ( .A1(n105645), .A2(n109625), .B1(n90520), .B2(n109620), 
        .ZN(n92875) );
  NOR4_X1 U78426 ( .A1(n92877), .A2(n92878), .A3(n92879), .A4(n92880), .ZN(
        n92863) );
  NAND2_X1 U78427 ( .A1(n92881), .A2(n92882), .ZN(n92880) );
  AOI22_X1 U78428 ( .A1(n90527), .A2(n109602), .B1(n90528), .B2(n72600), .ZN(
        n92882) );
  AOI22_X1 U78429 ( .A1(n90529), .A2(n109605), .B1(n90530), .B2(n72597), .ZN(
        n92881) );
  NAND2_X1 U78430 ( .A1(n92883), .A2(n92884), .ZN(n92879) );
  AOI22_X1 U78431 ( .A1(n90533), .A2(n109610), .B1(n90534), .B2(n109601), .ZN(
        n92884) );
  AOI22_X1 U78432 ( .A1(n90535), .A2(n109604), .B1(n90536), .B2(n72603), .ZN(
        n92883) );
  NAND2_X1 U78433 ( .A1(n92885), .A2(n92886), .ZN(n92878) );
  AOI22_X1 U78434 ( .A1(n90539), .A2(n109607), .B1(n90540), .B2(n72607), .ZN(
        n92886) );
  AOI22_X1 U78435 ( .A1(n90541), .A2(n109612), .B1(n90542), .B2(n109609), .ZN(
        n92885) );
  NAND2_X1 U78436 ( .A1(n92887), .A2(n92888), .ZN(n92877) );
  AOI22_X1 U78437 ( .A1(n90545), .A2(n72615), .B1(n90546), .B2(n109606), .ZN(
        n92888) );
  AOI22_X1 U78438 ( .A1(n90547), .A2(n109608), .B1(n90548), .B2(n109611), .ZN(
        n92887) );
  AOI21_X1 U78439 ( .B1(n90295), .B2(n88918), .A(n92890), .ZN(n92889) );
  OAI21_X1 U78440 ( .B1(n92891), .B2(n90298), .A(n92892), .ZN(n92890) );
  OAI21_X1 U78441 ( .B1(n92893), .B2(n92894), .A(n105658), .ZN(n92892) );
  OAI21_X1 U78442 ( .B1(n101842), .B2(n105657), .A(n92895), .ZN(n92894) );
  AOI22_X1 U78443 ( .A1(n105656), .A2(n108607), .B1(n105655), .B2(n71315), 
        .ZN(n92895) );
  NAND2_X1 U78444 ( .A1(n92896), .A2(n92897), .ZN(n92893) );
  AOI22_X1 U78445 ( .A1(n105654), .A2(n108612), .B1(n90310), .B2(n108609), 
        .ZN(n92897) );
  AOI22_X1 U78446 ( .A1(n90311), .A2(n71313), .B1(n105652), .B2(n108608), .ZN(
        n92896) );
  NOR4_X1 U78447 ( .A1(n92898), .A2(n92899), .A3(n92900), .A4(n92901), .ZN(
        n92891) );
  NAND2_X1 U78448 ( .A1(n92902), .A2(n92903), .ZN(n92901) );
  NOR4_X1 U78449 ( .A1(n92904), .A2(n92905), .A3(n92906), .A4(n92907), .ZN(
        n92903) );
  NAND2_X1 U78450 ( .A1(n92908), .A2(n92909), .ZN(n92907) );
  AOI22_X1 U78451 ( .A1(n90325), .A2(n108588), .B1(n90326), .B2(n108589), .ZN(
        n92909) );
  AOI22_X1 U78452 ( .A1(n90327), .A2(n108597), .B1(n90328), .B2(n108595), .ZN(
        n92908) );
  NAND2_X1 U78453 ( .A1(n92910), .A2(n92911), .ZN(n92906) );
  AOI22_X1 U78454 ( .A1(n90331), .A2(n71182), .B1(n90332), .B2(n108592), .ZN(
        n92911) );
  AOI22_X1 U78455 ( .A1(n90333), .A2(n71286), .B1(n90334), .B2(n108511), .ZN(
        n92910) );
  NAND2_X1 U78456 ( .A1(n92912), .A2(n92913), .ZN(n92905) );
  AOI22_X1 U78457 ( .A1(n90337), .A2(n108515), .B1(n90338), .B2(n71186), .ZN(
        n92913) );
  AOI22_X1 U78458 ( .A1(n90339), .A2(n108593), .B1(n90340), .B2(n108590), .ZN(
        n92912) );
  NAND2_X1 U78459 ( .A1(n92914), .A2(n92915), .ZN(n92904) );
  AOI22_X1 U78460 ( .A1(n90343), .A2(n108513), .B1(n90344), .B2(n108517), .ZN(
        n92915) );
  AOI22_X1 U78461 ( .A1(n90345), .A2(n108516), .B1(n90346), .B2(n71188), .ZN(
        n92914) );
  NOR4_X1 U78462 ( .A1(n92916), .A2(n92917), .A3(n92918), .A4(n92919), .ZN(
        n92902) );
  NAND2_X1 U78463 ( .A1(n92920), .A2(n92921), .ZN(n92919) );
  AOI22_X1 U78464 ( .A1(n90353), .A2(n108598), .B1(n90354), .B2(n108601), .ZN(
        n92921) );
  AOI22_X1 U78465 ( .A1(n90355), .A2(n108602), .B1(n90356), .B2(n108604), .ZN(
        n92920) );
  NAND2_X1 U78466 ( .A1(n92922), .A2(n92923), .ZN(n92918) );
  AOI22_X1 U78467 ( .A1(n90359), .A2(n108603), .B1(n90360), .B2(n108599), .ZN(
        n92923) );
  AOI22_X1 U78468 ( .A1(n90361), .A2(n108605), .B1(n90362), .B2(n108600), .ZN(
        n92922) );
  NAND2_X1 U78469 ( .A1(n92924), .A2(n92925), .ZN(n92917) );
  AOI22_X1 U78470 ( .A1(n90365), .A2(n71296), .B1(n90366), .B2(n71295), .ZN(
        n92925) );
  AOI22_X1 U78471 ( .A1(n90367), .A2(n71298), .B1(n90368), .B2(n108606), .ZN(
        n92924) );
  NAND2_X1 U78472 ( .A1(n92926), .A2(n92927), .ZN(n92916) );
  AOI22_X1 U78473 ( .A1(n90371), .A2(n108591), .B1(n90372), .B2(n108596), .ZN(
        n92927) );
  AOI22_X1 U78474 ( .A1(n90373), .A2(n71293), .B1(n90374), .B2(n108594), .ZN(
        n92926) );
  NAND2_X1 U78475 ( .A1(n92928), .A2(n92929), .ZN(n92900) );
  NOR4_X1 U78476 ( .A1(n92930), .A2(n92931), .A3(n92932), .A4(n92933), .ZN(
        n92929) );
  NAND2_X1 U78477 ( .A1(n92934), .A2(n92935), .ZN(n92933) );
  AOI22_X1 U78478 ( .A1(n90383), .A2(n108526), .B1(n90384), .B2(n108528), .ZN(
        n92935) );
  AOI22_X1 U78479 ( .A1(n90385), .A2(n71211), .B1(n90386), .B2(n108527), .ZN(
        n92934) );
  NAND2_X1 U78480 ( .A1(n92936), .A2(n92937), .ZN(n92932) );
  AOI22_X1 U78481 ( .A1(n90389), .A2(n71215), .B1(n90390), .B2(n71217), .ZN(
        n92937) );
  AOI22_X1 U78482 ( .A1(n90391), .A2(n108534), .B1(n90392), .B2(n108535), .ZN(
        n92936) );
  NAND2_X1 U78483 ( .A1(n92938), .A2(n92939), .ZN(n92931) );
  AOI22_X1 U78484 ( .A1(n90395), .A2(n108531), .B1(n90396), .B2(n108533), .ZN(
        n92939) );
  AOI22_X1 U78485 ( .A1(n90397), .A2(n108536), .B1(n90398), .B2(n108532), .ZN(
        n92938) );
  NAND2_X1 U78486 ( .A1(n92940), .A2(n92941), .ZN(n92930) );
  AOI22_X1 U78487 ( .A1(n90401), .A2(n108541), .B1(n90402), .B2(n71222), .ZN(
        n92941) );
  AOI22_X1 U78488 ( .A1(n90403), .A2(n108540), .B1(n90404), .B2(n71220), .ZN(
        n92940) );
  NOR4_X1 U78489 ( .A1(n92942), .A2(n92943), .A3(n92944), .A4(n92945), .ZN(
        n92928) );
  NAND2_X1 U78490 ( .A1(n92946), .A2(n92947), .ZN(n92945) );
  AOI22_X1 U78491 ( .A1(n90411), .A2(n108521), .B1(n90412), .B2(n108512), .ZN(
        n92947) );
  AOI22_X1 U78492 ( .A1(n90413), .A2(n108514), .B1(n90414), .B2(n71194), .ZN(
        n92946) );
  NAND2_X1 U78493 ( .A1(n92948), .A2(n92949), .ZN(n92944) );
  AOI22_X1 U78494 ( .A1(n90417), .A2(n108519), .B1(n90418), .B2(n108523), .ZN(
        n92949) );
  AOI22_X1 U78495 ( .A1(n90419), .A2(n108525), .B1(n90420), .B2(n108522), .ZN(
        n92948) );
  NAND2_X1 U78496 ( .A1(n92950), .A2(n92951), .ZN(n92943) );
  AOI22_X1 U78497 ( .A1(n90423), .A2(n71203), .B1(n90424), .B2(n108518), .ZN(
        n92951) );
  AOI22_X1 U78498 ( .A1(n90425), .A2(n108520), .B1(n90426), .B2(n108524), .ZN(
        n92950) );
  NAND2_X1 U78499 ( .A1(n92952), .A2(n92953), .ZN(n92942) );
  AOI22_X1 U78500 ( .A1(n90429), .A2(n108530), .B1(n90430), .B2(n71207), .ZN(
        n92953) );
  AOI22_X1 U78501 ( .A1(n90431), .A2(n71205), .B1(n90432), .B2(n108529), .ZN(
        n92952) );
  NAND2_X1 U78502 ( .A1(n92954), .A2(n92955), .ZN(n92899) );
  NOR4_X1 U78503 ( .A1(n92956), .A2(n92957), .A3(n92958), .A4(n92959), .ZN(
        n92955) );
  NAND2_X1 U78504 ( .A1(n92960), .A2(n92961), .ZN(n92959) );
  AOI22_X1 U78505 ( .A1(n90441), .A2(n71245), .B1(n90442), .B2(n108551), .ZN(
        n92961) );
  AOI22_X1 U78506 ( .A1(n90443), .A2(n108555), .B1(n90444), .B2(n108554), .ZN(
        n92960) );
  NAND2_X1 U78507 ( .A1(n92962), .A2(n92963), .ZN(n92958) );
  AOI22_X1 U78508 ( .A1(n90447), .A2(n108560), .B1(n90448), .B2(n108559), .ZN(
        n92963) );
  AOI22_X1 U78509 ( .A1(n90449), .A2(n108550), .B1(n90450), .B2(n108552), .ZN(
        n92962) );
  NAND2_X1 U78510 ( .A1(n92964), .A2(n92965), .ZN(n92957) );
  AOI22_X1 U78511 ( .A1(n90453), .A2(n108561), .B1(n90454), .B2(n108557), .ZN(
        n92965) );
  AOI22_X1 U78512 ( .A1(n90455), .A2(n71249), .B1(n90456), .B2(n71251), .ZN(
        n92964) );
  NAND2_X1 U78513 ( .A1(n92966), .A2(n92967), .ZN(n92956) );
  AOI22_X1 U78514 ( .A1(n90459), .A2(n108564), .B1(n90460), .B2(n71257), .ZN(
        n92967) );
  AOI22_X1 U78515 ( .A1(n90461), .A2(n108556), .B1(n90462), .B2(n108558), .ZN(
        n92966) );
  NOR4_X1 U78516 ( .A1(n92968), .A2(n92969), .A3(n92970), .A4(n92971), .ZN(
        n92954) );
  NAND2_X1 U78517 ( .A1(n92972), .A2(n92973), .ZN(n92971) );
  AOI22_X1 U78518 ( .A1(n90469), .A2(n108539), .B1(n90470), .B2(n108544), .ZN(
        n92973) );
  AOI22_X1 U78519 ( .A1(n90471), .A2(n108538), .B1(n90472), .B2(n71225), .ZN(
        n92972) );
  NAND2_X1 U78520 ( .A1(n92974), .A2(n92975), .ZN(n92970) );
  AOI22_X1 U78521 ( .A1(n90475), .A2(n71234), .B1(n90476), .B2(n108546), .ZN(
        n92975) );
  AOI22_X1 U78522 ( .A1(n90477), .A2(n108547), .B1(n90478), .B2(n108537), .ZN(
        n92974) );
  NAND2_X1 U78523 ( .A1(n92976), .A2(n92977), .ZN(n92969) );
  AOI22_X1 U78524 ( .A1(n90481), .A2(n108545), .B1(n90482), .B2(n108549), .ZN(
        n92977) );
  AOI22_X1 U78525 ( .A1(n90483), .A2(n108543), .B1(n90484), .B2(n108548), .ZN(
        n92976) );
  NAND2_X1 U78526 ( .A1(n92978), .A2(n92979), .ZN(n92968) );
  AOI22_X1 U78527 ( .A1(n90487), .A2(n71239), .B1(n90488), .B2(n108553), .ZN(
        n92979) );
  AOI22_X1 U78528 ( .A1(n90489), .A2(n71237), .B1(n90490), .B2(n108542), .ZN(
        n92978) );
  NAND2_X1 U78529 ( .A1(n92980), .A2(n92981), .ZN(n92898) );
  NOR4_X1 U78530 ( .A1(n92982), .A2(n92983), .A3(n92984), .A4(n92985), .ZN(
        n92981) );
  NAND2_X1 U78531 ( .A1(n92986), .A2(n92987), .ZN(n92985) );
  AOI22_X1 U78532 ( .A1(n90499), .A2(n108580), .B1(n90500), .B2(n108579), .ZN(
        n92987) );
  AOI22_X1 U78533 ( .A1(n90501), .A2(n71273), .B1(n90502), .B2(n108577), .ZN(
        n92986) );
  NAND2_X1 U78534 ( .A1(n92988), .A2(n92989), .ZN(n92984) );
  AOI22_X1 U78535 ( .A1(n90505), .A2(n108575), .B1(n90506), .B2(n108578), .ZN(
        n92989) );
  AOI22_X1 U78536 ( .A1(n105651), .A2(n71279), .B1(n90508), .B2(n108576), .ZN(
        n92988) );
  NAND2_X1 U78537 ( .A1(n92990), .A2(n92991), .ZN(n92983) );
  AOI22_X1 U78538 ( .A1(n90511), .A2(n108586), .B1(n105649), .B2(n71285), .ZN(
        n92991) );
  AOI22_X1 U78539 ( .A1(n105648), .A2(n108584), .B1(n105647), .B2(n108585), 
        .ZN(n92990) );
  NAND2_X1 U78540 ( .A1(n92992), .A2(n92993), .ZN(n92982) );
  AOI22_X1 U78541 ( .A1(n90517), .A2(n108581), .B1(n105646), .B2(n108583), 
        .ZN(n92993) );
  AOI22_X1 U78542 ( .A1(n105645), .A2(n108587), .B1(n90520), .B2(n108582), 
        .ZN(n92992) );
  NOR4_X1 U78543 ( .A1(n92994), .A2(n92995), .A3(n92996), .A4(n92997), .ZN(
        n92980) );
  NAND2_X1 U78544 ( .A1(n92998), .A2(n92999), .ZN(n92997) );
  AOI22_X1 U78545 ( .A1(n90527), .A2(n108563), .B1(n90528), .B2(n108567), .ZN(
        n92999) );
  AOI22_X1 U78546 ( .A1(n90529), .A2(n108566), .B1(n90530), .B2(n71256), .ZN(
        n92998) );
  NAND2_X1 U78547 ( .A1(n93000), .A2(n93001), .ZN(n92996) );
  AOI22_X1 U78548 ( .A1(n90533), .A2(n108572), .B1(n90534), .B2(n108562), .ZN(
        n93001) );
  AOI22_X1 U78549 ( .A1(n90535), .A2(n108565), .B1(n90536), .B2(n71262), .ZN(
        n93000) );
  NAND2_X1 U78550 ( .A1(n93002), .A2(n93003), .ZN(n92995) );
  AOI22_X1 U78551 ( .A1(n90539), .A2(n108569), .B1(n90540), .B2(n71266), .ZN(
        n93003) );
  AOI22_X1 U78552 ( .A1(n90541), .A2(n108574), .B1(n90542), .B2(n108571), .ZN(
        n93002) );
  NAND2_X1 U78553 ( .A1(n93004), .A2(n93005), .ZN(n92994) );
  AOI22_X1 U78554 ( .A1(n90545), .A2(n71274), .B1(n90546), .B2(n108568), .ZN(
        n93005) );
  AOI22_X1 U78555 ( .A1(n90547), .A2(n108570), .B1(n90548), .B2(n108573), .ZN(
        n93004) );
  AOI21_X1 U78556 ( .B1(n90295), .B2(n81794), .A(n93007), .ZN(n93006) );
  OAI21_X1 U78557 ( .B1(n93008), .B2(n90298), .A(n93009), .ZN(n93007) );
  OAI21_X1 U78558 ( .B1(n93010), .B2(n93011), .A(n105658), .ZN(n93009) );
  OAI21_X1 U78559 ( .B1(n101824), .B2(n105657), .A(n93012), .ZN(n93011) );
  AOI22_X1 U78560 ( .A1(n105656), .A2(n109752), .B1(n105655), .B2(n72798), 
        .ZN(n93012) );
  NAND2_X1 U78561 ( .A1(n93013), .A2(n93014), .ZN(n93010) );
  AOI22_X1 U78562 ( .A1(n105654), .A2(n109757), .B1(n90310), .B2(n109754), 
        .ZN(n93014) );
  AOI22_X1 U78563 ( .A1(n90311), .A2(n72796), .B1(n105652), .B2(n109753), .ZN(
        n93013) );
  NOR4_X1 U78564 ( .A1(n93015), .A2(n93016), .A3(n93017), .A4(n93018), .ZN(
        n93008) );
  NAND2_X1 U78565 ( .A1(n93019), .A2(n93020), .ZN(n93018) );
  NOR4_X1 U78566 ( .A1(n93021), .A2(n93022), .A3(n93023), .A4(n93024), .ZN(
        n93020) );
  NAND2_X1 U78567 ( .A1(n93025), .A2(n93026), .ZN(n93024) );
  AOI22_X1 U78568 ( .A1(n90325), .A2(n109733), .B1(n90326), .B2(n109734), .ZN(
        n93026) );
  AOI22_X1 U78569 ( .A1(n90327), .A2(n109742), .B1(n90328), .B2(n109740), .ZN(
        n93025) );
  NAND2_X1 U78570 ( .A1(n93027), .A2(n93028), .ZN(n93023) );
  AOI22_X1 U78571 ( .A1(n90331), .A2(n72665), .B1(n90332), .B2(n109737), .ZN(
        n93028) );
  AOI22_X1 U78572 ( .A1(n90333), .A2(n72769), .B1(n90334), .B2(n109655), .ZN(
        n93027) );
  NAND2_X1 U78573 ( .A1(n93029), .A2(n93030), .ZN(n93022) );
  AOI22_X1 U78574 ( .A1(n90337), .A2(n109659), .B1(n90338), .B2(n72669), .ZN(
        n93030) );
  AOI22_X1 U78575 ( .A1(n90339), .A2(n109738), .B1(n90340), .B2(n109735), .ZN(
        n93029) );
  NAND2_X1 U78576 ( .A1(n93031), .A2(n93032), .ZN(n93021) );
  AOI22_X1 U78577 ( .A1(n90343), .A2(n109657), .B1(n90344), .B2(n109661), .ZN(
        n93032) );
  AOI22_X1 U78578 ( .A1(n90345), .A2(n109660), .B1(n90346), .B2(n72671), .ZN(
        n93031) );
  NOR4_X1 U78579 ( .A1(n93033), .A2(n93034), .A3(n93035), .A4(n93036), .ZN(
        n93019) );
  NAND2_X1 U78580 ( .A1(n93037), .A2(n93038), .ZN(n93036) );
  AOI22_X1 U78581 ( .A1(n90353), .A2(n109743), .B1(n90354), .B2(n109746), .ZN(
        n93038) );
  AOI22_X1 U78582 ( .A1(n90355), .A2(n109747), .B1(n90356), .B2(n109749), .ZN(
        n93037) );
  NAND2_X1 U78583 ( .A1(n93039), .A2(n93040), .ZN(n93035) );
  AOI22_X1 U78584 ( .A1(n90359), .A2(n109748), .B1(n90360), .B2(n109744), .ZN(
        n93040) );
  AOI22_X1 U78585 ( .A1(n90361), .A2(n109750), .B1(n90362), .B2(n109745), .ZN(
        n93039) );
  NAND2_X1 U78586 ( .A1(n93041), .A2(n93042), .ZN(n93034) );
  AOI22_X1 U78587 ( .A1(n90365), .A2(n72779), .B1(n90366), .B2(n72778), .ZN(
        n93042) );
  AOI22_X1 U78588 ( .A1(n90367), .A2(n72781), .B1(n90368), .B2(n109751), .ZN(
        n93041) );
  NAND2_X1 U78589 ( .A1(n93043), .A2(n93044), .ZN(n93033) );
  AOI22_X1 U78590 ( .A1(n90371), .A2(n109736), .B1(n90372), .B2(n109741), .ZN(
        n93044) );
  AOI22_X1 U78591 ( .A1(n90373), .A2(n72776), .B1(n90374), .B2(n109739), .ZN(
        n93043) );
  NAND2_X1 U78592 ( .A1(n93045), .A2(n93046), .ZN(n93017) );
  NOR4_X1 U78593 ( .A1(n93047), .A2(n93048), .A3(n93049), .A4(n93050), .ZN(
        n93046) );
  NAND2_X1 U78594 ( .A1(n93051), .A2(n93052), .ZN(n93050) );
  AOI22_X1 U78595 ( .A1(n90383), .A2(n109670), .B1(n90384), .B2(n109672), .ZN(
        n93052) );
  AOI22_X1 U78596 ( .A1(n90385), .A2(n72694), .B1(n90386), .B2(n109671), .ZN(
        n93051) );
  NAND2_X1 U78597 ( .A1(n93053), .A2(n93054), .ZN(n93049) );
  AOI22_X1 U78598 ( .A1(n90389), .A2(n72698), .B1(n90390), .B2(n72700), .ZN(
        n93054) );
  AOI22_X1 U78599 ( .A1(n90391), .A2(n109678), .B1(n90392), .B2(n109679), .ZN(
        n93053) );
  NAND2_X1 U78600 ( .A1(n93055), .A2(n93056), .ZN(n93048) );
  AOI22_X1 U78601 ( .A1(n90395), .A2(n109675), .B1(n90396), .B2(n109677), .ZN(
        n93056) );
  AOI22_X1 U78602 ( .A1(n90397), .A2(n109680), .B1(n90398), .B2(n109676), .ZN(
        n93055) );
  NAND2_X1 U78603 ( .A1(n93057), .A2(n93058), .ZN(n93047) );
  AOI22_X1 U78604 ( .A1(n90401), .A2(n109685), .B1(n90402), .B2(n72705), .ZN(
        n93058) );
  AOI22_X1 U78605 ( .A1(n90403), .A2(n109684), .B1(n90404), .B2(n72703), .ZN(
        n93057) );
  NOR4_X1 U78606 ( .A1(n93059), .A2(n93060), .A3(n93061), .A4(n93062), .ZN(
        n93045) );
  NAND2_X1 U78607 ( .A1(n93063), .A2(n93064), .ZN(n93062) );
  AOI22_X1 U78608 ( .A1(n90411), .A2(n109665), .B1(n90412), .B2(n109656), .ZN(
        n93064) );
  AOI22_X1 U78609 ( .A1(n90413), .A2(n109658), .B1(n90414), .B2(n72677), .ZN(
        n93063) );
  NAND2_X1 U78610 ( .A1(n93065), .A2(n93066), .ZN(n93061) );
  AOI22_X1 U78611 ( .A1(n90417), .A2(n109663), .B1(n90418), .B2(n109667), .ZN(
        n93066) );
  AOI22_X1 U78612 ( .A1(n90419), .A2(n109669), .B1(n90420), .B2(n109666), .ZN(
        n93065) );
  NAND2_X1 U78613 ( .A1(n93067), .A2(n93068), .ZN(n93060) );
  AOI22_X1 U78614 ( .A1(n90423), .A2(n72686), .B1(n90424), .B2(n109662), .ZN(
        n93068) );
  AOI22_X1 U78615 ( .A1(n90425), .A2(n109664), .B1(n90426), .B2(n109668), .ZN(
        n93067) );
  NAND2_X1 U78616 ( .A1(n93069), .A2(n93070), .ZN(n93059) );
  AOI22_X1 U78617 ( .A1(n90429), .A2(n109674), .B1(n90430), .B2(n72690), .ZN(
        n93070) );
  AOI22_X1 U78618 ( .A1(n90431), .A2(n72688), .B1(n90432), .B2(n109673), .ZN(
        n93069) );
  NAND2_X1 U78619 ( .A1(n93071), .A2(n93072), .ZN(n93016) );
  NOR4_X1 U78620 ( .A1(n93073), .A2(n93074), .A3(n93075), .A4(n93076), .ZN(
        n93072) );
  NAND2_X1 U78621 ( .A1(n93077), .A2(n93078), .ZN(n93076) );
  AOI22_X1 U78622 ( .A1(n90441), .A2(n72728), .B1(n90442), .B2(n109695), .ZN(
        n93078) );
  AOI22_X1 U78623 ( .A1(n90443), .A2(n109699), .B1(n90444), .B2(n109698), .ZN(
        n93077) );
  NAND2_X1 U78624 ( .A1(n93079), .A2(n93080), .ZN(n93075) );
  AOI22_X1 U78625 ( .A1(n90447), .A2(n109704), .B1(n90448), .B2(n109703), .ZN(
        n93080) );
  AOI22_X1 U78626 ( .A1(n90449), .A2(n109694), .B1(n90450), .B2(n109696), .ZN(
        n93079) );
  NAND2_X1 U78627 ( .A1(n93081), .A2(n93082), .ZN(n93074) );
  AOI22_X1 U78628 ( .A1(n90453), .A2(n109705), .B1(n90454), .B2(n109701), .ZN(
        n93082) );
  AOI22_X1 U78629 ( .A1(n90455), .A2(n72732), .B1(n90456), .B2(n72734), .ZN(
        n93081) );
  NAND2_X1 U78630 ( .A1(n93083), .A2(n93084), .ZN(n93073) );
  AOI22_X1 U78631 ( .A1(n90459), .A2(n109708), .B1(n90460), .B2(n72740), .ZN(
        n93084) );
  AOI22_X1 U78632 ( .A1(n90461), .A2(n109700), .B1(n90462), .B2(n109702), .ZN(
        n93083) );
  NOR4_X1 U78633 ( .A1(n93085), .A2(n93086), .A3(n93087), .A4(n93088), .ZN(
        n93071) );
  NAND2_X1 U78634 ( .A1(n93089), .A2(n93090), .ZN(n93088) );
  AOI22_X1 U78635 ( .A1(n90469), .A2(n109683), .B1(n90470), .B2(n109688), .ZN(
        n93090) );
  AOI22_X1 U78636 ( .A1(n90471), .A2(n109682), .B1(n90472), .B2(n72708), .ZN(
        n93089) );
  NAND2_X1 U78637 ( .A1(n93091), .A2(n93092), .ZN(n93087) );
  AOI22_X1 U78638 ( .A1(n90475), .A2(n72717), .B1(n90476), .B2(n109690), .ZN(
        n93092) );
  AOI22_X1 U78639 ( .A1(n90477), .A2(n109691), .B1(n90478), .B2(n109681), .ZN(
        n93091) );
  NAND2_X1 U78640 ( .A1(n93093), .A2(n93094), .ZN(n93086) );
  AOI22_X1 U78641 ( .A1(n90481), .A2(n109689), .B1(n90482), .B2(n109693), .ZN(
        n93094) );
  AOI22_X1 U78642 ( .A1(n90483), .A2(n109687), .B1(n90484), .B2(n109692), .ZN(
        n93093) );
  NAND2_X1 U78643 ( .A1(n93095), .A2(n93096), .ZN(n93085) );
  AOI22_X1 U78644 ( .A1(n90487), .A2(n72722), .B1(n90488), .B2(n109697), .ZN(
        n93096) );
  AOI22_X1 U78645 ( .A1(n90489), .A2(n72720), .B1(n90490), .B2(n109686), .ZN(
        n93095) );
  NAND2_X1 U78646 ( .A1(n93097), .A2(n93098), .ZN(n93015) );
  NOR4_X1 U78647 ( .A1(n93099), .A2(n93100), .A3(n93101), .A4(n93102), .ZN(
        n93098) );
  NAND2_X1 U78648 ( .A1(n93103), .A2(n93104), .ZN(n93102) );
  AOI22_X1 U78649 ( .A1(n90499), .A2(n109725), .B1(n90500), .B2(n109724), .ZN(
        n93104) );
  AOI22_X1 U78650 ( .A1(n90501), .A2(n72756), .B1(n90502), .B2(n109722), .ZN(
        n93103) );
  NAND2_X1 U78651 ( .A1(n93105), .A2(n93106), .ZN(n93101) );
  AOI22_X1 U78652 ( .A1(n90505), .A2(n109720), .B1(n90506), .B2(n109723), .ZN(
        n93106) );
  AOI22_X1 U78653 ( .A1(n105651), .A2(n72762), .B1(n90508), .B2(n109721), .ZN(
        n93105) );
  NAND2_X1 U78654 ( .A1(n93107), .A2(n93108), .ZN(n93100) );
  AOI22_X1 U78655 ( .A1(n90511), .A2(n109731), .B1(n105649), .B2(n72768), .ZN(
        n93108) );
  AOI22_X1 U78656 ( .A1(n105648), .A2(n109729), .B1(n105647), .B2(n109730), 
        .ZN(n93107) );
  NAND2_X1 U78657 ( .A1(n93109), .A2(n93110), .ZN(n93099) );
  AOI22_X1 U78658 ( .A1(n90517), .A2(n109726), .B1(n105646), .B2(n109728), 
        .ZN(n93110) );
  AOI22_X1 U78659 ( .A1(n105645), .A2(n109732), .B1(n105644), .B2(n109727), 
        .ZN(n93109) );
  NOR4_X1 U78660 ( .A1(n93111), .A2(n93112), .A3(n93113), .A4(n93114), .ZN(
        n93097) );
  NAND2_X1 U78661 ( .A1(n93115), .A2(n93116), .ZN(n93114) );
  AOI22_X1 U78662 ( .A1(n90527), .A2(n109707), .B1(n90528), .B2(n109711), .ZN(
        n93116) );
  AOI22_X1 U78663 ( .A1(n90529), .A2(n109710), .B1(n90530), .B2(n72739), .ZN(
        n93115) );
  NAND2_X1 U78664 ( .A1(n93117), .A2(n93118), .ZN(n93113) );
  AOI22_X1 U78665 ( .A1(n90533), .A2(n109716), .B1(n90534), .B2(n109706), .ZN(
        n93118) );
  AOI22_X1 U78666 ( .A1(n90535), .A2(n109709), .B1(n90536), .B2(n72745), .ZN(
        n93117) );
  NAND2_X1 U78667 ( .A1(n93119), .A2(n93120), .ZN(n93112) );
  AOI22_X1 U78668 ( .A1(n90539), .A2(n109713), .B1(n90540), .B2(n109717), .ZN(
        n93120) );
  AOI22_X1 U78669 ( .A1(n90541), .A2(n109719), .B1(n90542), .B2(n109715), .ZN(
        n93119) );
  NAND2_X1 U78670 ( .A1(n93121), .A2(n93122), .ZN(n93111) );
  AOI22_X1 U78671 ( .A1(n90545), .A2(n72757), .B1(n90546), .B2(n109712), .ZN(
        n93122) );
  AOI22_X1 U78672 ( .A1(n90547), .A2(n109714), .B1(n90548), .B2(n109718), .ZN(
        n93121) );
  AOI21_X1 U78673 ( .B1(n90295), .B2(n89153), .A(n93124), .ZN(n93123) );
  OAI21_X1 U78674 ( .B1(n93125), .B2(n90298), .A(n93126), .ZN(n93124) );
  OAI21_X1 U78675 ( .B1(n93127), .B2(n93128), .A(n105658), .ZN(n93126) );
  OAI21_X1 U78676 ( .B1(n101806), .B2(n105657), .A(n93129), .ZN(n93128) );
  AOI22_X1 U78677 ( .A1(n105656), .A2(n109537), .B1(n105655), .B2(n72508), 
        .ZN(n93129) );
  NAND2_X1 U78678 ( .A1(n93130), .A2(n93131), .ZN(n93127) );
  AOI22_X1 U78679 ( .A1(n105654), .A2(n109542), .B1(n90310), .B2(n109539), 
        .ZN(n93131) );
  AOI22_X1 U78680 ( .A1(n90311), .A2(n72506), .B1(n105652), .B2(n109538), .ZN(
        n93130) );
  NOR4_X1 U78681 ( .A1(n93132), .A2(n93133), .A3(n93134), .A4(n93135), .ZN(
        n93125) );
  NAND2_X1 U78682 ( .A1(n93136), .A2(n93137), .ZN(n93135) );
  NOR4_X1 U78683 ( .A1(n93138), .A2(n93139), .A3(n93140), .A4(n93141), .ZN(
        n93137) );
  NAND2_X1 U78684 ( .A1(n93142), .A2(n93143), .ZN(n93141) );
  AOI22_X1 U78685 ( .A1(n90325), .A2(n109518), .B1(n90326), .B2(n109519), .ZN(
        n93143) );
  AOI22_X1 U78686 ( .A1(n90327), .A2(n109527), .B1(n90328), .B2(n109525), .ZN(
        n93142) );
  NAND2_X1 U78687 ( .A1(n93144), .A2(n93145), .ZN(n93140) );
  AOI22_X1 U78688 ( .A1(n90331), .A2(n72375), .B1(n90332), .B2(n109522), .ZN(
        n93145) );
  AOI22_X1 U78689 ( .A1(n90333), .A2(n72479), .B1(n90334), .B2(n109439), .ZN(
        n93144) );
  NAND2_X1 U78690 ( .A1(n93146), .A2(n93147), .ZN(n93139) );
  AOI22_X1 U78691 ( .A1(n90337), .A2(n109443), .B1(n90338), .B2(n72379), .ZN(
        n93147) );
  AOI22_X1 U78692 ( .A1(n90339), .A2(n109523), .B1(n90340), .B2(n109520), .ZN(
        n93146) );
  NAND2_X1 U78693 ( .A1(n93148), .A2(n93149), .ZN(n93138) );
  AOI22_X1 U78694 ( .A1(n90343), .A2(n109441), .B1(n90344), .B2(n109445), .ZN(
        n93149) );
  AOI22_X1 U78695 ( .A1(n90345), .A2(n109444), .B1(n90346), .B2(n72381), .ZN(
        n93148) );
  NOR4_X1 U78696 ( .A1(n93150), .A2(n93151), .A3(n93152), .A4(n93153), .ZN(
        n93136) );
  NAND2_X1 U78697 ( .A1(n93154), .A2(n93155), .ZN(n93153) );
  AOI22_X1 U78698 ( .A1(n90353), .A2(n109528), .B1(n90354), .B2(n109531), .ZN(
        n93155) );
  AOI22_X1 U78699 ( .A1(n90355), .A2(n109532), .B1(n90356), .B2(n109534), .ZN(
        n93154) );
  NAND2_X1 U78700 ( .A1(n93156), .A2(n93157), .ZN(n93152) );
  AOI22_X1 U78701 ( .A1(n90359), .A2(n109533), .B1(n90360), .B2(n109529), .ZN(
        n93157) );
  AOI22_X1 U78702 ( .A1(n90361), .A2(n109535), .B1(n90362), .B2(n109530), .ZN(
        n93156) );
  NAND2_X1 U78703 ( .A1(n93158), .A2(n93159), .ZN(n93151) );
  AOI22_X1 U78704 ( .A1(n90365), .A2(n72489), .B1(n90366), .B2(n72488), .ZN(
        n93159) );
  AOI22_X1 U78705 ( .A1(n90367), .A2(n72491), .B1(n90368), .B2(n109536), .ZN(
        n93158) );
  NAND2_X1 U78706 ( .A1(n93160), .A2(n93161), .ZN(n93150) );
  AOI22_X1 U78707 ( .A1(n90371), .A2(n109521), .B1(n90372), .B2(n109526), .ZN(
        n93161) );
  AOI22_X1 U78708 ( .A1(n90373), .A2(n72486), .B1(n90374), .B2(n109524), .ZN(
        n93160) );
  NAND2_X1 U78709 ( .A1(n93162), .A2(n93163), .ZN(n93134) );
  NOR4_X1 U78710 ( .A1(n93164), .A2(n93165), .A3(n93166), .A4(n93167), .ZN(
        n93163) );
  NAND2_X1 U78711 ( .A1(n93168), .A2(n93169), .ZN(n93167) );
  AOI22_X1 U78712 ( .A1(n90383), .A2(n109454), .B1(n90384), .B2(n109456), .ZN(
        n93169) );
  AOI22_X1 U78713 ( .A1(n90385), .A2(n72404), .B1(n90386), .B2(n109455), .ZN(
        n93168) );
  NAND2_X1 U78714 ( .A1(n93170), .A2(n93171), .ZN(n93166) );
  AOI22_X1 U78715 ( .A1(n90389), .A2(n72408), .B1(n90390), .B2(n72410), .ZN(
        n93171) );
  AOI22_X1 U78716 ( .A1(n90391), .A2(n109462), .B1(n90392), .B2(n109463), .ZN(
        n93170) );
  NAND2_X1 U78717 ( .A1(n93172), .A2(n93173), .ZN(n93165) );
  AOI22_X1 U78718 ( .A1(n90395), .A2(n109459), .B1(n90396), .B2(n109461), .ZN(
        n93173) );
  AOI22_X1 U78719 ( .A1(n90397), .A2(n109464), .B1(n90398), .B2(n109460), .ZN(
        n93172) );
  NAND2_X1 U78720 ( .A1(n93174), .A2(n93175), .ZN(n93164) );
  AOI22_X1 U78721 ( .A1(n90401), .A2(n109469), .B1(n90402), .B2(n72415), .ZN(
        n93175) );
  AOI22_X1 U78722 ( .A1(n90403), .A2(n109468), .B1(n90404), .B2(n72413), .ZN(
        n93174) );
  NOR4_X1 U78723 ( .A1(n93176), .A2(n93177), .A3(n93178), .A4(n93179), .ZN(
        n93162) );
  NAND2_X1 U78724 ( .A1(n93180), .A2(n93181), .ZN(n93179) );
  AOI22_X1 U78725 ( .A1(n90411), .A2(n109449), .B1(n90412), .B2(n109440), .ZN(
        n93181) );
  AOI22_X1 U78726 ( .A1(n90413), .A2(n109442), .B1(n90414), .B2(n72387), .ZN(
        n93180) );
  NAND2_X1 U78727 ( .A1(n93182), .A2(n93183), .ZN(n93178) );
  AOI22_X1 U78728 ( .A1(n90417), .A2(n109447), .B1(n90418), .B2(n109451), .ZN(
        n93183) );
  AOI22_X1 U78729 ( .A1(n90419), .A2(n109453), .B1(n90420), .B2(n109450), .ZN(
        n93182) );
  NAND2_X1 U78730 ( .A1(n93184), .A2(n93185), .ZN(n93177) );
  AOI22_X1 U78731 ( .A1(n90423), .A2(n72396), .B1(n90424), .B2(n109446), .ZN(
        n93185) );
  AOI22_X1 U78732 ( .A1(n90425), .A2(n109448), .B1(n90426), .B2(n109452), .ZN(
        n93184) );
  NAND2_X1 U78733 ( .A1(n93186), .A2(n93187), .ZN(n93176) );
  AOI22_X1 U78734 ( .A1(n90429), .A2(n109458), .B1(n90430), .B2(n72400), .ZN(
        n93187) );
  AOI22_X1 U78735 ( .A1(n90431), .A2(n72398), .B1(n90432), .B2(n109457), .ZN(
        n93186) );
  NAND2_X1 U78736 ( .A1(n93188), .A2(n93189), .ZN(n93133) );
  NOR4_X1 U78737 ( .A1(n93190), .A2(n93191), .A3(n93192), .A4(n93193), .ZN(
        n93189) );
  NAND2_X1 U78738 ( .A1(n93194), .A2(n93195), .ZN(n93193) );
  AOI22_X1 U78739 ( .A1(n90441), .A2(n72438), .B1(n90442), .B2(n109479), .ZN(
        n93195) );
  AOI22_X1 U78740 ( .A1(n90443), .A2(n109483), .B1(n90444), .B2(n109482), .ZN(
        n93194) );
  NAND2_X1 U78741 ( .A1(n93196), .A2(n93197), .ZN(n93192) );
  AOI22_X1 U78742 ( .A1(n90447), .A2(n109488), .B1(n90448), .B2(n109487), .ZN(
        n93197) );
  AOI22_X1 U78743 ( .A1(n90449), .A2(n109478), .B1(n90450), .B2(n109480), .ZN(
        n93196) );
  NAND2_X1 U78744 ( .A1(n93198), .A2(n93199), .ZN(n93191) );
  AOI22_X1 U78745 ( .A1(n90453), .A2(n109489), .B1(n90454), .B2(n109485), .ZN(
        n93199) );
  AOI22_X1 U78746 ( .A1(n90455), .A2(n72442), .B1(n90456), .B2(n72444), .ZN(
        n93198) );
  NAND2_X1 U78747 ( .A1(n93200), .A2(n93201), .ZN(n93190) );
  AOI22_X1 U78748 ( .A1(n90459), .A2(n109492), .B1(n90460), .B2(n72450), .ZN(
        n93201) );
  AOI22_X1 U78749 ( .A1(n90461), .A2(n109484), .B1(n90462), .B2(n109486), .ZN(
        n93200) );
  NOR4_X1 U78750 ( .A1(n93202), .A2(n93203), .A3(n93204), .A4(n93205), .ZN(
        n93188) );
  NAND2_X1 U78751 ( .A1(n93206), .A2(n93207), .ZN(n93205) );
  AOI22_X1 U78752 ( .A1(n90469), .A2(n109467), .B1(n90470), .B2(n109472), .ZN(
        n93207) );
  AOI22_X1 U78753 ( .A1(n90471), .A2(n109466), .B1(n90472), .B2(n72418), .ZN(
        n93206) );
  NAND2_X1 U78754 ( .A1(n93208), .A2(n93209), .ZN(n93204) );
  AOI22_X1 U78755 ( .A1(n90475), .A2(n72427), .B1(n90476), .B2(n109474), .ZN(
        n93209) );
  AOI22_X1 U78756 ( .A1(n90477), .A2(n109475), .B1(n90478), .B2(n109465), .ZN(
        n93208) );
  NAND2_X1 U78757 ( .A1(n93210), .A2(n93211), .ZN(n93203) );
  AOI22_X1 U78758 ( .A1(n90481), .A2(n109473), .B1(n90482), .B2(n109477), .ZN(
        n93211) );
  AOI22_X1 U78759 ( .A1(n90483), .A2(n109471), .B1(n90484), .B2(n109476), .ZN(
        n93210) );
  NAND2_X1 U78760 ( .A1(n93212), .A2(n93213), .ZN(n93202) );
  AOI22_X1 U78761 ( .A1(n90487), .A2(n72432), .B1(n90488), .B2(n109481), .ZN(
        n93213) );
  AOI22_X1 U78762 ( .A1(n90489), .A2(n72430), .B1(n90490), .B2(n109470), .ZN(
        n93212) );
  NAND2_X1 U78763 ( .A1(n93214), .A2(n93215), .ZN(n93132) );
  NOR4_X1 U78764 ( .A1(n93216), .A2(n93217), .A3(n93218), .A4(n93219), .ZN(
        n93215) );
  NAND2_X1 U78765 ( .A1(n93220), .A2(n93221), .ZN(n93219) );
  AOI22_X1 U78766 ( .A1(n90499), .A2(n109510), .B1(n90500), .B2(n109509), .ZN(
        n93221) );
  AOI22_X1 U78767 ( .A1(n90501), .A2(n72466), .B1(n90502), .B2(n109507), .ZN(
        n93220) );
  NAND2_X1 U78768 ( .A1(n93222), .A2(n93223), .ZN(n93218) );
  AOI22_X1 U78769 ( .A1(n90505), .A2(n109505), .B1(n90506), .B2(n109508), .ZN(
        n93223) );
  AOI22_X1 U78770 ( .A1(n105651), .A2(n72472), .B1(n90508), .B2(n109506), .ZN(
        n93222) );
  NAND2_X1 U78771 ( .A1(n93224), .A2(n93225), .ZN(n93217) );
  AOI22_X1 U78772 ( .A1(n90511), .A2(n109516), .B1(n105649), .B2(n72478), .ZN(
        n93225) );
  AOI22_X1 U78773 ( .A1(n105648), .A2(n109514), .B1(n105647), .B2(n109515), 
        .ZN(n93224) );
  NAND2_X1 U78774 ( .A1(n93226), .A2(n93227), .ZN(n93216) );
  AOI22_X1 U78775 ( .A1(n90517), .A2(n109511), .B1(n105646), .B2(n109513), 
        .ZN(n93227) );
  AOI22_X1 U78776 ( .A1(n105645), .A2(n109517), .B1(n90520), .B2(n109512), 
        .ZN(n93226) );
  NOR4_X1 U78777 ( .A1(n93228), .A2(n93229), .A3(n93230), .A4(n93231), .ZN(
        n93214) );
  NAND2_X1 U78778 ( .A1(n93232), .A2(n93233), .ZN(n93231) );
  AOI22_X1 U78779 ( .A1(n90527), .A2(n109491), .B1(n90528), .B2(n109495), .ZN(
        n93233) );
  AOI22_X1 U78780 ( .A1(n90529), .A2(n109494), .B1(n90530), .B2(n72449), .ZN(
        n93232) );
  NAND2_X1 U78781 ( .A1(n93234), .A2(n93235), .ZN(n93230) );
  AOI22_X1 U78782 ( .A1(n90533), .A2(n109501), .B1(n90534), .B2(n109490), .ZN(
        n93235) );
  AOI22_X1 U78783 ( .A1(n90535), .A2(n109493), .B1(n90536), .B2(n109498), .ZN(
        n93234) );
  NAND2_X1 U78784 ( .A1(n93236), .A2(n93237), .ZN(n93229) );
  AOI22_X1 U78785 ( .A1(n90539), .A2(n109497), .B1(n90540), .B2(n109502), .ZN(
        n93237) );
  AOI22_X1 U78786 ( .A1(n90541), .A2(n109504), .B1(n90542), .B2(n109500), .ZN(
        n93236) );
  NAND2_X1 U78787 ( .A1(n93238), .A2(n93239), .ZN(n93228) );
  AOI22_X1 U78788 ( .A1(n90545), .A2(n72467), .B1(n90546), .B2(n109496), .ZN(
        n93239) );
  AOI22_X1 U78789 ( .A1(n90547), .A2(n109499), .B1(n90548), .B2(n109503), .ZN(
        n93238) );
  AOI21_X1 U78790 ( .B1(n90295), .B2(n89271), .A(n93241), .ZN(n93240) );
  OAI21_X1 U78791 ( .B1(n93242), .B2(n90298), .A(n93243), .ZN(n93241) );
  OAI21_X1 U78792 ( .B1(n93244), .B2(n93245), .A(n105658), .ZN(n93243) );
  OAI21_X1 U78793 ( .B1(n101790), .B2(n105657), .A(n93246), .ZN(n93245) );
  AOI22_X1 U78794 ( .A1(n105656), .A2(n109075), .B1(n105655), .B2(n71908), 
        .ZN(n93246) );
  NAND2_X1 U78795 ( .A1(n93247), .A2(n93248), .ZN(n93244) );
  AOI22_X1 U78796 ( .A1(n105654), .A2(n109080), .B1(n90310), .B2(n109077), 
        .ZN(n93248) );
  AOI22_X1 U78797 ( .A1(n90311), .A2(n71906), .B1(n105652), .B2(n109076), .ZN(
        n93247) );
  NOR4_X1 U78798 ( .A1(n93249), .A2(n93250), .A3(n93251), .A4(n93252), .ZN(
        n93242) );
  NAND2_X1 U78799 ( .A1(n93253), .A2(n93254), .ZN(n93252) );
  NOR4_X1 U78800 ( .A1(n93255), .A2(n93256), .A3(n93257), .A4(n93258), .ZN(
        n93254) );
  NAND2_X1 U78801 ( .A1(n93259), .A2(n93260), .ZN(n93258) );
  AOI22_X1 U78802 ( .A1(n90325), .A2(n109056), .B1(n90326), .B2(n109057), .ZN(
        n93260) );
  AOI22_X1 U78803 ( .A1(n90327), .A2(n109065), .B1(n90328), .B2(n109063), .ZN(
        n93259) );
  NAND2_X1 U78804 ( .A1(n93261), .A2(n93262), .ZN(n93257) );
  AOI22_X1 U78805 ( .A1(n90331), .A2(n71775), .B1(n90332), .B2(n109060), .ZN(
        n93262) );
  AOI22_X1 U78806 ( .A1(n90333), .A2(n71879), .B1(n90334), .B2(n108976), .ZN(
        n93261) );
  NAND2_X1 U78807 ( .A1(n93263), .A2(n93264), .ZN(n93256) );
  AOI22_X1 U78808 ( .A1(n90337), .A2(n108980), .B1(n90338), .B2(n71779), .ZN(
        n93264) );
  AOI22_X1 U78809 ( .A1(n90339), .A2(n109061), .B1(n90340), .B2(n109058), .ZN(
        n93263) );
  NAND2_X1 U78810 ( .A1(n93265), .A2(n93266), .ZN(n93255) );
  AOI22_X1 U78811 ( .A1(n90343), .A2(n108978), .B1(n90344), .B2(n108982), .ZN(
        n93266) );
  AOI22_X1 U78812 ( .A1(n90345), .A2(n108981), .B1(n90346), .B2(n71781), .ZN(
        n93265) );
  NOR4_X1 U78813 ( .A1(n93267), .A2(n93268), .A3(n93269), .A4(n93270), .ZN(
        n93253) );
  NAND2_X1 U78814 ( .A1(n93271), .A2(n93272), .ZN(n93270) );
  AOI22_X1 U78815 ( .A1(n90353), .A2(n109066), .B1(n90354), .B2(n109069), .ZN(
        n93272) );
  AOI22_X1 U78816 ( .A1(n90355), .A2(n109070), .B1(n90356), .B2(n109072), .ZN(
        n93271) );
  NAND2_X1 U78817 ( .A1(n93273), .A2(n93274), .ZN(n93269) );
  AOI22_X1 U78818 ( .A1(n90359), .A2(n109071), .B1(n90360), .B2(n109067), .ZN(
        n93274) );
  AOI22_X1 U78819 ( .A1(n90361), .A2(n109073), .B1(n90362), .B2(n109068), .ZN(
        n93273) );
  NAND2_X1 U78820 ( .A1(n93275), .A2(n93276), .ZN(n93268) );
  AOI22_X1 U78821 ( .A1(n90365), .A2(n71889), .B1(n90366), .B2(n71888), .ZN(
        n93276) );
  AOI22_X1 U78822 ( .A1(n90367), .A2(n71891), .B1(n90368), .B2(n109074), .ZN(
        n93275) );
  NAND2_X1 U78823 ( .A1(n93277), .A2(n93278), .ZN(n93267) );
  AOI22_X1 U78824 ( .A1(n90371), .A2(n109059), .B1(n90372), .B2(n109064), .ZN(
        n93278) );
  AOI22_X1 U78825 ( .A1(n90373), .A2(n71886), .B1(n90374), .B2(n109062), .ZN(
        n93277) );
  NAND2_X1 U78826 ( .A1(n93279), .A2(n93280), .ZN(n93251) );
  NOR4_X1 U78827 ( .A1(n93281), .A2(n93282), .A3(n93283), .A4(n93284), .ZN(
        n93280) );
  NAND2_X1 U78828 ( .A1(n93285), .A2(n93286), .ZN(n93284) );
  AOI22_X1 U78829 ( .A1(n90383), .A2(n108991), .B1(n90384), .B2(n108993), .ZN(
        n93286) );
  AOI22_X1 U78830 ( .A1(n90385), .A2(n71804), .B1(n90386), .B2(n108992), .ZN(
        n93285) );
  NAND2_X1 U78831 ( .A1(n93287), .A2(n93288), .ZN(n93283) );
  AOI22_X1 U78832 ( .A1(n90389), .A2(n71808), .B1(n90390), .B2(n71810), .ZN(
        n93288) );
  AOI22_X1 U78833 ( .A1(n90391), .A2(n108999), .B1(n90392), .B2(n109000), .ZN(
        n93287) );
  NAND2_X1 U78834 ( .A1(n93289), .A2(n93290), .ZN(n93282) );
  AOI22_X1 U78835 ( .A1(n90395), .A2(n108996), .B1(n90396), .B2(n108998), .ZN(
        n93290) );
  AOI22_X1 U78836 ( .A1(n90397), .A2(n109001), .B1(n90398), .B2(n108997), .ZN(
        n93289) );
  NAND2_X1 U78837 ( .A1(n93291), .A2(n93292), .ZN(n93281) );
  AOI22_X1 U78838 ( .A1(n90401), .A2(n109006), .B1(n90402), .B2(n71815), .ZN(
        n93292) );
  AOI22_X1 U78839 ( .A1(n90403), .A2(n109005), .B1(n90404), .B2(n71813), .ZN(
        n93291) );
  NOR4_X1 U78840 ( .A1(n93293), .A2(n93294), .A3(n93295), .A4(n93296), .ZN(
        n93279) );
  NAND2_X1 U78841 ( .A1(n93297), .A2(n93298), .ZN(n93296) );
  AOI22_X1 U78842 ( .A1(n90411), .A2(n108986), .B1(n90412), .B2(n108977), .ZN(
        n93298) );
  AOI22_X1 U78843 ( .A1(n90413), .A2(n108979), .B1(n90414), .B2(n71787), .ZN(
        n93297) );
  NAND2_X1 U78844 ( .A1(n93299), .A2(n93300), .ZN(n93295) );
  AOI22_X1 U78845 ( .A1(n90417), .A2(n108984), .B1(n90418), .B2(n108988), .ZN(
        n93300) );
  AOI22_X1 U78846 ( .A1(n90419), .A2(n108990), .B1(n90420), .B2(n108987), .ZN(
        n93299) );
  NAND2_X1 U78847 ( .A1(n93301), .A2(n93302), .ZN(n93294) );
  AOI22_X1 U78848 ( .A1(n90423), .A2(n71796), .B1(n90424), .B2(n108983), .ZN(
        n93302) );
  AOI22_X1 U78849 ( .A1(n90425), .A2(n108985), .B1(n90426), .B2(n108989), .ZN(
        n93301) );
  NAND2_X1 U78850 ( .A1(n93303), .A2(n93304), .ZN(n93293) );
  AOI22_X1 U78851 ( .A1(n90429), .A2(n108995), .B1(n90430), .B2(n71800), .ZN(
        n93304) );
  AOI22_X1 U78852 ( .A1(n90431), .A2(n71798), .B1(n90432), .B2(n108994), .ZN(
        n93303) );
  NAND2_X1 U78853 ( .A1(n93305), .A2(n93306), .ZN(n93250) );
  NOR4_X1 U78854 ( .A1(n93307), .A2(n93308), .A3(n93309), .A4(n93310), .ZN(
        n93306) );
  NAND2_X1 U78855 ( .A1(n93311), .A2(n93312), .ZN(n93310) );
  AOI22_X1 U78856 ( .A1(n90441), .A2(n71838), .B1(n90442), .B2(n109016), .ZN(
        n93312) );
  AOI22_X1 U78857 ( .A1(n90443), .A2(n109020), .B1(n90444), .B2(n109019), .ZN(
        n93311) );
  NAND2_X1 U78858 ( .A1(n93313), .A2(n93314), .ZN(n93309) );
  AOI22_X1 U78859 ( .A1(n90447), .A2(n109025), .B1(n90448), .B2(n109024), .ZN(
        n93314) );
  AOI22_X1 U78860 ( .A1(n90449), .A2(n109015), .B1(n90450), .B2(n109017), .ZN(
        n93313) );
  NAND2_X1 U78861 ( .A1(n93315), .A2(n93316), .ZN(n93308) );
  AOI22_X1 U78862 ( .A1(n90453), .A2(n109026), .B1(n90454), .B2(n109022), .ZN(
        n93316) );
  AOI22_X1 U78863 ( .A1(n90455), .A2(n71842), .B1(n90456), .B2(n71844), .ZN(
        n93315) );
  NAND2_X1 U78864 ( .A1(n93317), .A2(n93318), .ZN(n93307) );
  AOI22_X1 U78865 ( .A1(n90459), .A2(n109029), .B1(n90460), .B2(n71850), .ZN(
        n93318) );
  AOI22_X1 U78866 ( .A1(n90461), .A2(n109021), .B1(n90462), .B2(n109023), .ZN(
        n93317) );
  NOR4_X1 U78867 ( .A1(n93319), .A2(n93320), .A3(n93321), .A4(n93322), .ZN(
        n93305) );
  NAND2_X1 U78868 ( .A1(n93323), .A2(n93324), .ZN(n93322) );
  AOI22_X1 U78869 ( .A1(n90469), .A2(n109004), .B1(n90470), .B2(n109009), .ZN(
        n93324) );
  AOI22_X1 U78870 ( .A1(n90471), .A2(n109003), .B1(n90472), .B2(n71818), .ZN(
        n93323) );
  NAND2_X1 U78871 ( .A1(n93325), .A2(n93326), .ZN(n93321) );
  AOI22_X1 U78872 ( .A1(n90475), .A2(n71827), .B1(n90476), .B2(n109011), .ZN(
        n93326) );
  AOI22_X1 U78873 ( .A1(n90477), .A2(n109012), .B1(n90478), .B2(n109002), .ZN(
        n93325) );
  NAND2_X1 U78874 ( .A1(n93327), .A2(n93328), .ZN(n93320) );
  AOI22_X1 U78875 ( .A1(n90481), .A2(n109010), .B1(n90482), .B2(n109014), .ZN(
        n93328) );
  AOI22_X1 U78876 ( .A1(n90483), .A2(n109008), .B1(n90484), .B2(n109013), .ZN(
        n93327) );
  NAND2_X1 U78877 ( .A1(n93329), .A2(n93330), .ZN(n93319) );
  AOI22_X1 U78878 ( .A1(n90487), .A2(n71832), .B1(n90488), .B2(n109018), .ZN(
        n93330) );
  AOI22_X1 U78879 ( .A1(n90489), .A2(n71830), .B1(n90490), .B2(n109007), .ZN(
        n93329) );
  NAND2_X1 U78880 ( .A1(n93331), .A2(n93332), .ZN(n93249) );
  NOR4_X1 U78881 ( .A1(n93333), .A2(n93334), .A3(n93335), .A4(n93336), .ZN(
        n93332) );
  NAND2_X1 U78882 ( .A1(n93337), .A2(n93338), .ZN(n93336) );
  AOI22_X1 U78883 ( .A1(n90499), .A2(n109047), .B1(n90500), .B2(n109046), .ZN(
        n93338) );
  AOI22_X1 U78884 ( .A1(n90501), .A2(n71866), .B1(n90502), .B2(n109044), .ZN(
        n93337) );
  NAND2_X1 U78885 ( .A1(n93339), .A2(n93340), .ZN(n93335) );
  AOI22_X1 U78886 ( .A1(n90505), .A2(n109042), .B1(n90506), .B2(n109045), .ZN(
        n93340) );
  AOI22_X1 U78887 ( .A1(n105651), .A2(n71872), .B1(n90508), .B2(n109043), .ZN(
        n93339) );
  NAND2_X1 U78888 ( .A1(n93341), .A2(n93342), .ZN(n93334) );
  AOI22_X1 U78889 ( .A1(n90511), .A2(n109053), .B1(n105649), .B2(n71878), .ZN(
        n93342) );
  AOI22_X1 U78890 ( .A1(n105648), .A2(n109051), .B1(n105647), .B2(n109052), 
        .ZN(n93341) );
  NAND2_X1 U78891 ( .A1(n93343), .A2(n93344), .ZN(n93333) );
  AOI22_X1 U78892 ( .A1(n90517), .A2(n109048), .B1(n105646), .B2(n109050), 
        .ZN(n93344) );
  AOI22_X1 U78893 ( .A1(n105645), .A2(n109054), .B1(n105644), .B2(n109049), 
        .ZN(n93343) );
  NOR4_X1 U78894 ( .A1(n93345), .A2(n93346), .A3(n93347), .A4(n93348), .ZN(
        n93331) );
  NAND2_X1 U78895 ( .A1(n93349), .A2(n93350), .ZN(n93348) );
  AOI22_X1 U78896 ( .A1(n90527), .A2(n109028), .B1(n90528), .B2(n109032), .ZN(
        n93350) );
  AOI22_X1 U78897 ( .A1(n90529), .A2(n109031), .B1(n90530), .B2(n71849), .ZN(
        n93349) );
  NAND2_X1 U78898 ( .A1(n93351), .A2(n93352), .ZN(n93347) );
  AOI22_X1 U78899 ( .A1(n90533), .A2(n109038), .B1(n90534), .B2(n109027), .ZN(
        n93352) );
  AOI22_X1 U78900 ( .A1(n90535), .A2(n109030), .B1(n90536), .B2(n109035), .ZN(
        n93351) );
  NAND2_X1 U78901 ( .A1(n93353), .A2(n93354), .ZN(n93346) );
  AOI22_X1 U78902 ( .A1(n90539), .A2(n109034), .B1(n90540), .B2(n109039), .ZN(
        n93354) );
  AOI22_X1 U78903 ( .A1(n90541), .A2(n109041), .B1(n90542), .B2(n109037), .ZN(
        n93353) );
  NAND2_X1 U78904 ( .A1(n93355), .A2(n93356), .ZN(n93345) );
  AOI22_X1 U78905 ( .A1(n90545), .A2(n71867), .B1(n90546), .B2(n109033), .ZN(
        n93356) );
  AOI22_X1 U78906 ( .A1(n90547), .A2(n109036), .B1(n90548), .B2(n109040), .ZN(
        n93355) );
  AOI21_X1 U78907 ( .B1(n90295), .B2(n81792), .A(n93358), .ZN(n93357) );
  OAI21_X1 U78908 ( .B1(n93359), .B2(n90298), .A(n93360), .ZN(n93358) );
  OAI21_X1 U78909 ( .B1(n93361), .B2(n93362), .A(n105658), .ZN(n93360) );
  OAI21_X1 U78910 ( .B1(n101772), .B2(n105657), .A(n93363), .ZN(n93362) );
  AOI22_X1 U78911 ( .A1(n105656), .A2(n109422), .B1(n105655), .B2(n72357), 
        .ZN(n93363) );
  NAND2_X1 U78912 ( .A1(n93364), .A2(n93365), .ZN(n93361) );
  AOI22_X1 U78913 ( .A1(n105654), .A2(n109427), .B1(n90310), .B2(n109424), 
        .ZN(n93365) );
  AOI22_X1 U78914 ( .A1(n90311), .A2(n72355), .B1(n105652), .B2(n109423), .ZN(
        n93364) );
  NOR4_X1 U78915 ( .A1(n93366), .A2(n93367), .A3(n93368), .A4(n93369), .ZN(
        n93359) );
  NAND2_X1 U78916 ( .A1(n93370), .A2(n93371), .ZN(n93369) );
  NOR4_X1 U78917 ( .A1(n93372), .A2(n93373), .A3(n93374), .A4(n93375), .ZN(
        n93371) );
  NAND2_X1 U78918 ( .A1(n93376), .A2(n93377), .ZN(n93375) );
  AOI22_X1 U78919 ( .A1(n90325), .A2(n109403), .B1(n90326), .B2(n109404), .ZN(
        n93377) );
  AOI22_X1 U78920 ( .A1(n90327), .A2(n109412), .B1(n90328), .B2(n109410), .ZN(
        n93376) );
  NAND2_X1 U78921 ( .A1(n93378), .A2(n93379), .ZN(n93374) );
  AOI22_X1 U78922 ( .A1(n90331), .A2(n72224), .B1(n90332), .B2(n109407), .ZN(
        n93379) );
  AOI22_X1 U78923 ( .A1(n90333), .A2(n72328), .B1(n90334), .B2(n109324), .ZN(
        n93378) );
  NAND2_X1 U78924 ( .A1(n93380), .A2(n93381), .ZN(n93373) );
  AOI22_X1 U78925 ( .A1(n90337), .A2(n109328), .B1(n90338), .B2(n72228), .ZN(
        n93381) );
  AOI22_X1 U78926 ( .A1(n90339), .A2(n109408), .B1(n90340), .B2(n109405), .ZN(
        n93380) );
  NAND2_X1 U78927 ( .A1(n93382), .A2(n93383), .ZN(n93372) );
  AOI22_X1 U78928 ( .A1(n90343), .A2(n109326), .B1(n90344), .B2(n109330), .ZN(
        n93383) );
  AOI22_X1 U78929 ( .A1(n90345), .A2(n109329), .B1(n90346), .B2(n72230), .ZN(
        n93382) );
  NOR4_X1 U78930 ( .A1(n93384), .A2(n93385), .A3(n93386), .A4(n93387), .ZN(
        n93370) );
  NAND2_X1 U78931 ( .A1(n93388), .A2(n93389), .ZN(n93387) );
  AOI22_X1 U78932 ( .A1(n90353), .A2(n109413), .B1(n90354), .B2(n109416), .ZN(
        n93389) );
  AOI22_X1 U78933 ( .A1(n90355), .A2(n109417), .B1(n90356), .B2(n109419), .ZN(
        n93388) );
  NAND2_X1 U78934 ( .A1(n93390), .A2(n93391), .ZN(n93386) );
  AOI22_X1 U78935 ( .A1(n90359), .A2(n109418), .B1(n90360), .B2(n109414), .ZN(
        n93391) );
  AOI22_X1 U78936 ( .A1(n90361), .A2(n109420), .B1(n90362), .B2(n109415), .ZN(
        n93390) );
  NAND2_X1 U78937 ( .A1(n93392), .A2(n93393), .ZN(n93385) );
  AOI22_X1 U78938 ( .A1(n90365), .A2(n72338), .B1(n90366), .B2(n72337), .ZN(
        n93393) );
  AOI22_X1 U78939 ( .A1(n90367), .A2(n72340), .B1(n90368), .B2(n109421), .ZN(
        n93392) );
  NAND2_X1 U78940 ( .A1(n93394), .A2(n93395), .ZN(n93384) );
  AOI22_X1 U78941 ( .A1(n90371), .A2(n109406), .B1(n90372), .B2(n109411), .ZN(
        n93395) );
  AOI22_X1 U78942 ( .A1(n90373), .A2(n72335), .B1(n90374), .B2(n109409), .ZN(
        n93394) );
  NAND2_X1 U78943 ( .A1(n93396), .A2(n93397), .ZN(n93368) );
  NOR4_X1 U78944 ( .A1(n93398), .A2(n93399), .A3(n93400), .A4(n93401), .ZN(
        n93397) );
  NAND2_X1 U78945 ( .A1(n93402), .A2(n93403), .ZN(n93401) );
  AOI22_X1 U78946 ( .A1(n90383), .A2(n109339), .B1(n90384), .B2(n109341), .ZN(
        n93403) );
  AOI22_X1 U78947 ( .A1(n90385), .A2(n72253), .B1(n90386), .B2(n109340), .ZN(
        n93402) );
  NAND2_X1 U78948 ( .A1(n93404), .A2(n93405), .ZN(n93400) );
  AOI22_X1 U78949 ( .A1(n90389), .A2(n72257), .B1(n90390), .B2(n72259), .ZN(
        n93405) );
  AOI22_X1 U78950 ( .A1(n90391), .A2(n109347), .B1(n90392), .B2(n109348), .ZN(
        n93404) );
  NAND2_X1 U78951 ( .A1(n93406), .A2(n93407), .ZN(n93399) );
  AOI22_X1 U78952 ( .A1(n90395), .A2(n109344), .B1(n90396), .B2(n109346), .ZN(
        n93407) );
  AOI22_X1 U78953 ( .A1(n90397), .A2(n109349), .B1(n90398), .B2(n109345), .ZN(
        n93406) );
  NAND2_X1 U78954 ( .A1(n93408), .A2(n93409), .ZN(n93398) );
  AOI22_X1 U78955 ( .A1(n90401), .A2(n109354), .B1(n90402), .B2(n72264), .ZN(
        n93409) );
  AOI22_X1 U78956 ( .A1(n90403), .A2(n109353), .B1(n90404), .B2(n72262), .ZN(
        n93408) );
  NOR4_X1 U78957 ( .A1(n93410), .A2(n93411), .A3(n93412), .A4(n93413), .ZN(
        n93396) );
  NAND2_X1 U78958 ( .A1(n93414), .A2(n93415), .ZN(n93413) );
  AOI22_X1 U78959 ( .A1(n90411), .A2(n109334), .B1(n90412), .B2(n109325), .ZN(
        n93415) );
  AOI22_X1 U78960 ( .A1(n90413), .A2(n109327), .B1(n90414), .B2(n72236), .ZN(
        n93414) );
  NAND2_X1 U78961 ( .A1(n93416), .A2(n93417), .ZN(n93412) );
  AOI22_X1 U78962 ( .A1(n90417), .A2(n109332), .B1(n90418), .B2(n109336), .ZN(
        n93417) );
  AOI22_X1 U78963 ( .A1(n90419), .A2(n109338), .B1(n90420), .B2(n109335), .ZN(
        n93416) );
  NAND2_X1 U78964 ( .A1(n93418), .A2(n93419), .ZN(n93411) );
  AOI22_X1 U78965 ( .A1(n90423), .A2(n72245), .B1(n90424), .B2(n109331), .ZN(
        n93419) );
  AOI22_X1 U78966 ( .A1(n90425), .A2(n109333), .B1(n90426), .B2(n109337), .ZN(
        n93418) );
  NAND2_X1 U78967 ( .A1(n93420), .A2(n93421), .ZN(n93410) );
  AOI22_X1 U78968 ( .A1(n90429), .A2(n109343), .B1(n90430), .B2(n72249), .ZN(
        n93421) );
  AOI22_X1 U78969 ( .A1(n90431), .A2(n72247), .B1(n90432), .B2(n109342), .ZN(
        n93420) );
  NAND2_X1 U78970 ( .A1(n93422), .A2(n93423), .ZN(n93367) );
  NOR4_X1 U78971 ( .A1(n93424), .A2(n93425), .A3(n93426), .A4(n93427), .ZN(
        n93423) );
  NAND2_X1 U78972 ( .A1(n93428), .A2(n93429), .ZN(n93427) );
  AOI22_X1 U78973 ( .A1(n90441), .A2(n72287), .B1(n90442), .B2(n109364), .ZN(
        n93429) );
  AOI22_X1 U78974 ( .A1(n90443), .A2(n109368), .B1(n90444), .B2(n109367), .ZN(
        n93428) );
  NAND2_X1 U78975 ( .A1(n93430), .A2(n93431), .ZN(n93426) );
  AOI22_X1 U78976 ( .A1(n90447), .A2(n109373), .B1(n90448), .B2(n109372), .ZN(
        n93431) );
  AOI22_X1 U78977 ( .A1(n90449), .A2(n109363), .B1(n90450), .B2(n109365), .ZN(
        n93430) );
  NAND2_X1 U78978 ( .A1(n93432), .A2(n93433), .ZN(n93425) );
  AOI22_X1 U78979 ( .A1(n90453), .A2(n109374), .B1(n90454), .B2(n109370), .ZN(
        n93433) );
  AOI22_X1 U78980 ( .A1(n90455), .A2(n72291), .B1(n90456), .B2(n72293), .ZN(
        n93432) );
  NAND2_X1 U78981 ( .A1(n93434), .A2(n93435), .ZN(n93424) );
  AOI22_X1 U78982 ( .A1(n90459), .A2(n109377), .B1(n90460), .B2(n72299), .ZN(
        n93435) );
  AOI22_X1 U78983 ( .A1(n90461), .A2(n109369), .B1(n90462), .B2(n109371), .ZN(
        n93434) );
  NOR4_X1 U78984 ( .A1(n93436), .A2(n93437), .A3(n93438), .A4(n93439), .ZN(
        n93422) );
  NAND2_X1 U78985 ( .A1(n93440), .A2(n93441), .ZN(n93439) );
  AOI22_X1 U78986 ( .A1(n90469), .A2(n109352), .B1(n90470), .B2(n109357), .ZN(
        n93441) );
  AOI22_X1 U78987 ( .A1(n90471), .A2(n109351), .B1(n90472), .B2(n72267), .ZN(
        n93440) );
  NAND2_X1 U78988 ( .A1(n93442), .A2(n93443), .ZN(n93438) );
  AOI22_X1 U78989 ( .A1(n90475), .A2(n72276), .B1(n90476), .B2(n109359), .ZN(
        n93443) );
  AOI22_X1 U78990 ( .A1(n90477), .A2(n109360), .B1(n90478), .B2(n109350), .ZN(
        n93442) );
  NAND2_X1 U78991 ( .A1(n93444), .A2(n93445), .ZN(n93437) );
  AOI22_X1 U78992 ( .A1(n90481), .A2(n109358), .B1(n90482), .B2(n109362), .ZN(
        n93445) );
  AOI22_X1 U78993 ( .A1(n90483), .A2(n109356), .B1(n90484), .B2(n109361), .ZN(
        n93444) );
  NAND2_X1 U78994 ( .A1(n93446), .A2(n93447), .ZN(n93436) );
  AOI22_X1 U78995 ( .A1(n90487), .A2(n72281), .B1(n90488), .B2(n109366), .ZN(
        n93447) );
  AOI22_X1 U78996 ( .A1(n90489), .A2(n72279), .B1(n90490), .B2(n109355), .ZN(
        n93446) );
  NAND2_X1 U78997 ( .A1(n93448), .A2(n93449), .ZN(n93366) );
  NOR4_X1 U78998 ( .A1(n93450), .A2(n93451), .A3(n93452), .A4(n93453), .ZN(
        n93449) );
  NAND2_X1 U78999 ( .A1(n93454), .A2(n93455), .ZN(n93453) );
  AOI22_X1 U79000 ( .A1(n90499), .A2(n109395), .B1(n90500), .B2(n109394), .ZN(
        n93455) );
  AOI22_X1 U79001 ( .A1(n90501), .A2(n72315), .B1(n90502), .B2(n109392), .ZN(
        n93454) );
  NAND2_X1 U79002 ( .A1(n93456), .A2(n93457), .ZN(n93452) );
  AOI22_X1 U79003 ( .A1(n90505), .A2(n109390), .B1(n90506), .B2(n109393), .ZN(
        n93457) );
  AOI22_X1 U79004 ( .A1(n105651), .A2(n72321), .B1(n90508), .B2(n109391), .ZN(
        n93456) );
  NAND2_X1 U79005 ( .A1(n93458), .A2(n93459), .ZN(n93451) );
  AOI22_X1 U79006 ( .A1(n90511), .A2(n109401), .B1(n105649), .B2(n72327), .ZN(
        n93459) );
  AOI22_X1 U79007 ( .A1(n105648), .A2(n109399), .B1(n105647), .B2(n109400), 
        .ZN(n93458) );
  NAND2_X1 U79008 ( .A1(n93460), .A2(n93461), .ZN(n93450) );
  AOI22_X1 U79009 ( .A1(n90517), .A2(n109396), .B1(n105646), .B2(n109398), 
        .ZN(n93461) );
  AOI22_X1 U79010 ( .A1(n105645), .A2(n109402), .B1(n105644), .B2(n109397), 
        .ZN(n93460) );
  NOR4_X1 U79011 ( .A1(n93462), .A2(n93463), .A3(n93464), .A4(n93465), .ZN(
        n93448) );
  NAND2_X1 U79012 ( .A1(n93466), .A2(n93467), .ZN(n93465) );
  AOI22_X1 U79013 ( .A1(n90527), .A2(n109376), .B1(n90528), .B2(n109380), .ZN(
        n93467) );
  AOI22_X1 U79014 ( .A1(n90529), .A2(n109379), .B1(n90530), .B2(n72298), .ZN(
        n93466) );
  NAND2_X1 U79015 ( .A1(n93468), .A2(n93469), .ZN(n93464) );
  AOI22_X1 U79016 ( .A1(n90533), .A2(n109386), .B1(n90534), .B2(n109375), .ZN(
        n93469) );
  AOI22_X1 U79017 ( .A1(n90535), .A2(n109378), .B1(n90536), .B2(n109383), .ZN(
        n93468) );
  NAND2_X1 U79018 ( .A1(n93470), .A2(n93471), .ZN(n93463) );
  AOI22_X1 U79019 ( .A1(n90539), .A2(n109382), .B1(n90540), .B2(n109387), .ZN(
        n93471) );
  AOI22_X1 U79020 ( .A1(n90541), .A2(n109389), .B1(n90542), .B2(n109385), .ZN(
        n93470) );
  NAND2_X1 U79021 ( .A1(n93472), .A2(n93473), .ZN(n93462) );
  AOI22_X1 U79022 ( .A1(n90545), .A2(n72316), .B1(n90546), .B2(n109381), .ZN(
        n93473) );
  AOI22_X1 U79023 ( .A1(n90547), .A2(n109384), .B1(n90548), .B2(n109388), .ZN(
        n93472) );
  AOI21_X1 U79024 ( .B1(n90295), .B2(n89506), .A(n93475), .ZN(n93474) );
  OAI21_X1 U79025 ( .B1(n93476), .B2(n90298), .A(n93477), .ZN(n93475) );
  OAI21_X1 U79026 ( .B1(n93478), .B2(n93479), .A(n105658), .ZN(n93477) );
  OAI21_X1 U79027 ( .B1(n101756), .B2(n105657), .A(n93480), .ZN(n93479) );
  AOI22_X1 U79028 ( .A1(n105656), .A2(n109303), .B1(n105655), .B2(n72206), 
        .ZN(n93480) );
  NAND2_X1 U79029 ( .A1(n93481), .A2(n93482), .ZN(n93478) );
  AOI22_X1 U79030 ( .A1(n105654), .A2(n109308), .B1(n90310), .B2(n109305), 
        .ZN(n93482) );
  AOI22_X1 U79031 ( .A1(n90311), .A2(n72204), .B1(n105652), .B2(n109304), .ZN(
        n93481) );
  NOR4_X1 U79032 ( .A1(n93483), .A2(n93484), .A3(n93485), .A4(n93486), .ZN(
        n93476) );
  NAND2_X1 U79033 ( .A1(n93487), .A2(n93488), .ZN(n93486) );
  NOR4_X1 U79034 ( .A1(n93489), .A2(n93490), .A3(n93491), .A4(n93492), .ZN(
        n93488) );
  NAND2_X1 U79035 ( .A1(n93493), .A2(n93494), .ZN(n93492) );
  AOI22_X1 U79036 ( .A1(n90325), .A2(n109284), .B1(n90326), .B2(n109285), .ZN(
        n93494) );
  AOI22_X1 U79037 ( .A1(n90327), .A2(n109293), .B1(n90328), .B2(n109291), .ZN(
        n93493) );
  NAND2_X1 U79038 ( .A1(n93495), .A2(n93496), .ZN(n93491) );
  AOI22_X1 U79039 ( .A1(n90331), .A2(n72073), .B1(n90332), .B2(n109288), .ZN(
        n93496) );
  AOI22_X1 U79040 ( .A1(n90333), .A2(n72177), .B1(n90334), .B2(n109206), .ZN(
        n93495) );
  NAND2_X1 U79041 ( .A1(n93497), .A2(n93498), .ZN(n93490) );
  AOI22_X1 U79042 ( .A1(n90337), .A2(n109210), .B1(n90338), .B2(n72077), .ZN(
        n93498) );
  AOI22_X1 U79043 ( .A1(n90339), .A2(n109289), .B1(n90340), .B2(n109286), .ZN(
        n93497) );
  NAND2_X1 U79044 ( .A1(n93499), .A2(n93500), .ZN(n93489) );
  AOI22_X1 U79045 ( .A1(n90343), .A2(n109208), .B1(n90344), .B2(n109212), .ZN(
        n93500) );
  AOI22_X1 U79046 ( .A1(n90345), .A2(n109211), .B1(n90346), .B2(n72079), .ZN(
        n93499) );
  NOR4_X1 U79047 ( .A1(n93501), .A2(n93502), .A3(n93503), .A4(n93504), .ZN(
        n93487) );
  NAND2_X1 U79048 ( .A1(n93505), .A2(n93506), .ZN(n93504) );
  AOI22_X1 U79049 ( .A1(n90353), .A2(n109294), .B1(n90354), .B2(n109297), .ZN(
        n93506) );
  AOI22_X1 U79050 ( .A1(n90355), .A2(n109298), .B1(n90356), .B2(n109300), .ZN(
        n93505) );
  NAND2_X1 U79051 ( .A1(n93507), .A2(n93508), .ZN(n93503) );
  AOI22_X1 U79052 ( .A1(n90359), .A2(n109299), .B1(n90360), .B2(n109295), .ZN(
        n93508) );
  AOI22_X1 U79053 ( .A1(n90361), .A2(n109301), .B1(n90362), .B2(n109296), .ZN(
        n93507) );
  NAND2_X1 U79054 ( .A1(n93509), .A2(n93510), .ZN(n93502) );
  AOI22_X1 U79055 ( .A1(n90365), .A2(n72187), .B1(n90366), .B2(n72186), .ZN(
        n93510) );
  AOI22_X1 U79056 ( .A1(n90367), .A2(n72189), .B1(n90368), .B2(n109302), .ZN(
        n93509) );
  NAND2_X1 U79057 ( .A1(n93511), .A2(n93512), .ZN(n93501) );
  AOI22_X1 U79058 ( .A1(n90371), .A2(n109287), .B1(n90372), .B2(n109292), .ZN(
        n93512) );
  AOI22_X1 U79059 ( .A1(n90373), .A2(n72184), .B1(n90374), .B2(n109290), .ZN(
        n93511) );
  NAND2_X1 U79060 ( .A1(n93513), .A2(n93514), .ZN(n93485) );
  NOR4_X1 U79061 ( .A1(n93515), .A2(n93516), .A3(n93517), .A4(n93518), .ZN(
        n93514) );
  NAND2_X1 U79062 ( .A1(n93519), .A2(n93520), .ZN(n93518) );
  AOI22_X1 U79063 ( .A1(n90383), .A2(n109221), .B1(n90384), .B2(n109223), .ZN(
        n93520) );
  AOI22_X1 U79064 ( .A1(n90385), .A2(n72102), .B1(n90386), .B2(n109222), .ZN(
        n93519) );
  NAND2_X1 U79065 ( .A1(n93521), .A2(n93522), .ZN(n93517) );
  AOI22_X1 U79066 ( .A1(n90389), .A2(n72106), .B1(n90390), .B2(n72108), .ZN(
        n93522) );
  AOI22_X1 U79067 ( .A1(n90391), .A2(n109229), .B1(n90392), .B2(n109230), .ZN(
        n93521) );
  NAND2_X1 U79068 ( .A1(n93523), .A2(n93524), .ZN(n93516) );
  AOI22_X1 U79069 ( .A1(n90395), .A2(n109226), .B1(n90396), .B2(n109228), .ZN(
        n93524) );
  AOI22_X1 U79070 ( .A1(n90397), .A2(n109231), .B1(n90398), .B2(n109227), .ZN(
        n93523) );
  NAND2_X1 U79071 ( .A1(n93525), .A2(n93526), .ZN(n93515) );
  AOI22_X1 U79072 ( .A1(n90401), .A2(n109236), .B1(n90402), .B2(n72113), .ZN(
        n93526) );
  AOI22_X1 U79073 ( .A1(n90403), .A2(n109235), .B1(n90404), .B2(n72111), .ZN(
        n93525) );
  NOR4_X1 U79074 ( .A1(n93527), .A2(n93528), .A3(n93529), .A4(n93530), .ZN(
        n93513) );
  NAND2_X1 U79075 ( .A1(n93531), .A2(n93532), .ZN(n93530) );
  AOI22_X1 U79076 ( .A1(n90411), .A2(n109216), .B1(n90412), .B2(n109207), .ZN(
        n93532) );
  AOI22_X1 U79077 ( .A1(n90413), .A2(n109209), .B1(n90414), .B2(n72085), .ZN(
        n93531) );
  NAND2_X1 U79078 ( .A1(n93533), .A2(n93534), .ZN(n93529) );
  AOI22_X1 U79079 ( .A1(n90417), .A2(n109214), .B1(n90418), .B2(n109218), .ZN(
        n93534) );
  AOI22_X1 U79080 ( .A1(n90419), .A2(n109220), .B1(n90420), .B2(n109217), .ZN(
        n93533) );
  NAND2_X1 U79081 ( .A1(n93535), .A2(n93536), .ZN(n93528) );
  AOI22_X1 U79082 ( .A1(n90423), .A2(n72094), .B1(n90424), .B2(n109213), .ZN(
        n93536) );
  AOI22_X1 U79083 ( .A1(n90425), .A2(n109215), .B1(n90426), .B2(n109219), .ZN(
        n93535) );
  NAND2_X1 U79084 ( .A1(n93537), .A2(n93538), .ZN(n93527) );
  AOI22_X1 U79085 ( .A1(n90429), .A2(n109225), .B1(n90430), .B2(n72098), .ZN(
        n93538) );
  AOI22_X1 U79086 ( .A1(n90431), .A2(n72096), .B1(n90432), .B2(n109224), .ZN(
        n93537) );
  NAND2_X1 U79087 ( .A1(n93539), .A2(n93540), .ZN(n93484) );
  NOR4_X1 U79088 ( .A1(n93541), .A2(n93542), .A3(n93543), .A4(n93544), .ZN(
        n93540) );
  NAND2_X1 U79089 ( .A1(n93545), .A2(n93546), .ZN(n93544) );
  AOI22_X1 U79090 ( .A1(n90441), .A2(n72136), .B1(n90442), .B2(n109246), .ZN(
        n93546) );
  AOI22_X1 U79091 ( .A1(n90443), .A2(n109250), .B1(n90444), .B2(n109249), .ZN(
        n93545) );
  NAND2_X1 U79092 ( .A1(n93547), .A2(n93548), .ZN(n93543) );
  AOI22_X1 U79093 ( .A1(n90447), .A2(n109255), .B1(n90448), .B2(n109254), .ZN(
        n93548) );
  AOI22_X1 U79094 ( .A1(n90449), .A2(n109245), .B1(n90450), .B2(n109247), .ZN(
        n93547) );
  NAND2_X1 U79095 ( .A1(n93549), .A2(n93550), .ZN(n93542) );
  AOI22_X1 U79096 ( .A1(n90453), .A2(n109256), .B1(n90454), .B2(n109252), .ZN(
        n93550) );
  AOI22_X1 U79097 ( .A1(n90455), .A2(n72140), .B1(n90456), .B2(n72142), .ZN(
        n93549) );
  NAND2_X1 U79098 ( .A1(n93551), .A2(n93552), .ZN(n93541) );
  AOI22_X1 U79099 ( .A1(n90459), .A2(n109259), .B1(n90460), .B2(n72148), .ZN(
        n93552) );
  AOI22_X1 U79100 ( .A1(n90461), .A2(n109251), .B1(n90462), .B2(n109253), .ZN(
        n93551) );
  NOR4_X1 U79101 ( .A1(n93553), .A2(n93554), .A3(n93555), .A4(n93556), .ZN(
        n93539) );
  NAND2_X1 U79102 ( .A1(n93557), .A2(n93558), .ZN(n93556) );
  AOI22_X1 U79103 ( .A1(n90469), .A2(n109234), .B1(n90470), .B2(n109239), .ZN(
        n93558) );
  AOI22_X1 U79104 ( .A1(n90471), .A2(n109233), .B1(n90472), .B2(n72116), .ZN(
        n93557) );
  NAND2_X1 U79105 ( .A1(n93559), .A2(n93560), .ZN(n93555) );
  AOI22_X1 U79106 ( .A1(n90475), .A2(n72125), .B1(n90476), .B2(n109241), .ZN(
        n93560) );
  AOI22_X1 U79107 ( .A1(n90477), .A2(n109242), .B1(n90478), .B2(n109232), .ZN(
        n93559) );
  NAND2_X1 U79108 ( .A1(n93561), .A2(n93562), .ZN(n93554) );
  AOI22_X1 U79109 ( .A1(n90481), .A2(n109240), .B1(n90482), .B2(n109244), .ZN(
        n93562) );
  AOI22_X1 U79110 ( .A1(n90483), .A2(n109238), .B1(n90484), .B2(n109243), .ZN(
        n93561) );
  NAND2_X1 U79111 ( .A1(n93563), .A2(n93564), .ZN(n93553) );
  AOI22_X1 U79112 ( .A1(n90487), .A2(n72130), .B1(n90488), .B2(n109248), .ZN(
        n93564) );
  AOI22_X1 U79113 ( .A1(n90489), .A2(n72128), .B1(n90490), .B2(n109237), .ZN(
        n93563) );
  NAND2_X1 U79114 ( .A1(n93565), .A2(n93566), .ZN(n93483) );
  NOR4_X1 U79115 ( .A1(n93567), .A2(n93568), .A3(n93569), .A4(n93570), .ZN(
        n93566) );
  NAND2_X1 U79116 ( .A1(n93571), .A2(n93572), .ZN(n93570) );
  AOI22_X1 U79117 ( .A1(n90499), .A2(n109277), .B1(n90500), .B2(n109276), .ZN(
        n93572) );
  AOI22_X1 U79118 ( .A1(n90501), .A2(n72164), .B1(n90502), .B2(n109274), .ZN(
        n93571) );
  NAND2_X1 U79119 ( .A1(n93573), .A2(n93574), .ZN(n93569) );
  AOI22_X1 U79120 ( .A1(n90505), .A2(n109272), .B1(n90506), .B2(n109275), .ZN(
        n93574) );
  AOI22_X1 U79121 ( .A1(n105651), .A2(n72170), .B1(n90508), .B2(n109273), .ZN(
        n93573) );
  NAND2_X1 U79122 ( .A1(n93575), .A2(n93576), .ZN(n93568) );
  AOI22_X1 U79123 ( .A1(n90511), .A2(n109282), .B1(n105649), .B2(n72176), .ZN(
        n93576) );
  AOI22_X1 U79124 ( .A1(n105648), .A2(n109280), .B1(n105647), .B2(n109281), 
        .ZN(n93575) );
  NAND2_X1 U79125 ( .A1(n93577), .A2(n93578), .ZN(n93567) );
  AOI22_X1 U79126 ( .A1(n90517), .A2(n109278), .B1(n105646), .B2(n72171), .ZN(
        n93578) );
  AOI22_X1 U79127 ( .A1(n105645), .A2(n109283), .B1(n105644), .B2(n109279), 
        .ZN(n93577) );
  NOR4_X1 U79128 ( .A1(n93579), .A2(n93580), .A3(n93581), .A4(n93582), .ZN(
        n93565) );
  NAND2_X1 U79129 ( .A1(n93583), .A2(n93584), .ZN(n93582) );
  AOI22_X1 U79130 ( .A1(n90527), .A2(n109258), .B1(n90528), .B2(n109262), .ZN(
        n93584) );
  AOI22_X1 U79131 ( .A1(n90529), .A2(n109261), .B1(n90530), .B2(n72147), .ZN(
        n93583) );
  NAND2_X1 U79132 ( .A1(n93585), .A2(n93586), .ZN(n93581) );
  AOI22_X1 U79133 ( .A1(n90533), .A2(n109268), .B1(n90534), .B2(n109257), .ZN(
        n93586) );
  AOI22_X1 U79134 ( .A1(n90535), .A2(n109260), .B1(n90536), .B2(n109265), .ZN(
        n93585) );
  NAND2_X1 U79135 ( .A1(n93587), .A2(n93588), .ZN(n93580) );
  AOI22_X1 U79136 ( .A1(n90539), .A2(n109264), .B1(n90540), .B2(n109269), .ZN(
        n93588) );
  AOI22_X1 U79137 ( .A1(n90541), .A2(n109271), .B1(n90542), .B2(n109267), .ZN(
        n93587) );
  NAND2_X1 U79138 ( .A1(n93589), .A2(n93590), .ZN(n93579) );
  AOI22_X1 U79139 ( .A1(n90545), .A2(n72165), .B1(n90546), .B2(n109263), .ZN(
        n93590) );
  AOI22_X1 U79140 ( .A1(n90547), .A2(n109266), .B1(n90548), .B2(n109270), .ZN(
        n93589) );
  AOI21_X1 U79141 ( .B1(n90295), .B2(n89624), .A(n93592), .ZN(n93591) );
  OAI21_X1 U79142 ( .B1(n93593), .B2(n105659), .A(n93594), .ZN(n93592) );
  OAI21_X1 U79143 ( .B1(n93595), .B2(n93596), .A(n105658), .ZN(n93594) );
  OAI21_X1 U79144 ( .B1(n101738), .B2(n105657), .A(n93597), .ZN(n93596) );
  AOI22_X1 U79145 ( .A1(n105656), .A2(n109195), .B1(n105655), .B2(n72062), 
        .ZN(n93597) );
  NAND2_X1 U79146 ( .A1(n93598), .A2(n93599), .ZN(n93595) );
  AOI22_X1 U79147 ( .A1(n105654), .A2(n109200), .B1(n90310), .B2(n109197), 
        .ZN(n93599) );
  AOI22_X1 U79148 ( .A1(n90311), .A2(n72060), .B1(n105652), .B2(n109196), .ZN(
        n93598) );
  NOR4_X1 U79149 ( .A1(n93600), .A2(n93601), .A3(n93602), .A4(n93603), .ZN(
        n93593) );
  NAND2_X1 U79150 ( .A1(n93604), .A2(n93605), .ZN(n93603) );
  NOR4_X1 U79151 ( .A1(n93606), .A2(n93607), .A3(n93608), .A4(n93609), .ZN(
        n93605) );
  NAND2_X1 U79152 ( .A1(n93610), .A2(n93611), .ZN(n93609) );
  AOI22_X1 U79153 ( .A1(n90325), .A2(n109176), .B1(n90326), .B2(n109177), .ZN(
        n93611) );
  AOI22_X1 U79154 ( .A1(n90327), .A2(n109185), .B1(n90328), .B2(n109183), .ZN(
        n93610) );
  NAND2_X1 U79155 ( .A1(n93612), .A2(n93613), .ZN(n93608) );
  AOI22_X1 U79156 ( .A1(n90331), .A2(n71929), .B1(n90332), .B2(n109180), .ZN(
        n93613) );
  AOI22_X1 U79157 ( .A1(n90333), .A2(n72033), .B1(n90334), .B2(n109098), .ZN(
        n93612) );
  NAND2_X1 U79158 ( .A1(n93614), .A2(n93615), .ZN(n93607) );
  AOI22_X1 U79159 ( .A1(n90337), .A2(n109102), .B1(n90338), .B2(n71933), .ZN(
        n93615) );
  AOI22_X1 U79160 ( .A1(n90339), .A2(n109181), .B1(n90340), .B2(n109178), .ZN(
        n93614) );
  NAND2_X1 U79161 ( .A1(n93616), .A2(n93617), .ZN(n93606) );
  AOI22_X1 U79162 ( .A1(n90343), .A2(n109100), .B1(n90344), .B2(n109104), .ZN(
        n93617) );
  AOI22_X1 U79163 ( .A1(n90345), .A2(n109103), .B1(n90346), .B2(n71935), .ZN(
        n93616) );
  NOR4_X1 U79164 ( .A1(n93618), .A2(n93619), .A3(n93620), .A4(n93621), .ZN(
        n93604) );
  NAND2_X1 U79165 ( .A1(n93622), .A2(n93623), .ZN(n93621) );
  AOI22_X1 U79166 ( .A1(n90353), .A2(n109186), .B1(n90354), .B2(n109189), .ZN(
        n93623) );
  AOI22_X1 U79167 ( .A1(n90355), .A2(n109190), .B1(n90356), .B2(n109192), .ZN(
        n93622) );
  NAND2_X1 U79168 ( .A1(n93624), .A2(n93625), .ZN(n93620) );
  AOI22_X1 U79169 ( .A1(n90359), .A2(n109191), .B1(n90360), .B2(n109187), .ZN(
        n93625) );
  AOI22_X1 U79170 ( .A1(n90361), .A2(n109193), .B1(n90362), .B2(n109188), .ZN(
        n93624) );
  NAND2_X1 U79171 ( .A1(n93626), .A2(n93627), .ZN(n93619) );
  AOI22_X1 U79172 ( .A1(n90365), .A2(n72043), .B1(n90366), .B2(n72042), .ZN(
        n93627) );
  AOI22_X1 U79173 ( .A1(n90367), .A2(n72045), .B1(n90368), .B2(n109194), .ZN(
        n93626) );
  NAND2_X1 U79174 ( .A1(n93628), .A2(n93629), .ZN(n93618) );
  AOI22_X1 U79175 ( .A1(n90371), .A2(n109179), .B1(n90372), .B2(n109184), .ZN(
        n93629) );
  AOI22_X1 U79176 ( .A1(n90373), .A2(n72040), .B1(n90374), .B2(n109182), .ZN(
        n93628) );
  NAND2_X1 U79177 ( .A1(n93630), .A2(n93631), .ZN(n93602) );
  NOR4_X1 U79178 ( .A1(n93632), .A2(n93633), .A3(n93634), .A4(n93635), .ZN(
        n93631) );
  NAND2_X1 U79179 ( .A1(n93636), .A2(n93637), .ZN(n93635) );
  AOI22_X1 U79180 ( .A1(n90383), .A2(n109113), .B1(n90384), .B2(n109115), .ZN(
        n93637) );
  AOI22_X1 U79181 ( .A1(n90385), .A2(n71958), .B1(n90386), .B2(n109114), .ZN(
        n93636) );
  NAND2_X1 U79182 ( .A1(n93638), .A2(n93639), .ZN(n93634) );
  AOI22_X1 U79183 ( .A1(n90389), .A2(n71962), .B1(n90390), .B2(n71964), .ZN(
        n93639) );
  AOI22_X1 U79184 ( .A1(n90391), .A2(n109121), .B1(n90392), .B2(n109122), .ZN(
        n93638) );
  NAND2_X1 U79185 ( .A1(n93640), .A2(n93641), .ZN(n93633) );
  AOI22_X1 U79186 ( .A1(n90395), .A2(n109118), .B1(n90396), .B2(n109120), .ZN(
        n93641) );
  AOI22_X1 U79187 ( .A1(n90397), .A2(n109123), .B1(n90398), .B2(n109119), .ZN(
        n93640) );
  NAND2_X1 U79188 ( .A1(n93642), .A2(n93643), .ZN(n93632) );
  AOI22_X1 U79189 ( .A1(n90401), .A2(n109128), .B1(n90402), .B2(n71969), .ZN(
        n93643) );
  AOI22_X1 U79190 ( .A1(n90403), .A2(n109127), .B1(n90404), .B2(n71967), .ZN(
        n93642) );
  NOR4_X1 U79191 ( .A1(n93644), .A2(n93645), .A3(n93646), .A4(n93647), .ZN(
        n93630) );
  NAND2_X1 U79192 ( .A1(n93648), .A2(n93649), .ZN(n93647) );
  AOI22_X1 U79193 ( .A1(n90411), .A2(n109108), .B1(n90412), .B2(n109099), .ZN(
        n93649) );
  AOI22_X1 U79194 ( .A1(n90413), .A2(n109101), .B1(n90414), .B2(n71941), .ZN(
        n93648) );
  NAND2_X1 U79195 ( .A1(n93650), .A2(n93651), .ZN(n93646) );
  AOI22_X1 U79196 ( .A1(n90417), .A2(n109106), .B1(n90418), .B2(n109110), .ZN(
        n93651) );
  AOI22_X1 U79197 ( .A1(n90419), .A2(n109112), .B1(n90420), .B2(n109109), .ZN(
        n93650) );
  NAND2_X1 U79198 ( .A1(n93652), .A2(n93653), .ZN(n93645) );
  AOI22_X1 U79199 ( .A1(n90423), .A2(n71950), .B1(n90424), .B2(n109105), .ZN(
        n93653) );
  AOI22_X1 U79200 ( .A1(n90425), .A2(n109107), .B1(n90426), .B2(n109111), .ZN(
        n93652) );
  NAND2_X1 U79201 ( .A1(n93654), .A2(n93655), .ZN(n93644) );
  AOI22_X1 U79202 ( .A1(n90429), .A2(n109117), .B1(n90430), .B2(n71954), .ZN(
        n93655) );
  AOI22_X1 U79203 ( .A1(n90431), .A2(n71952), .B1(n90432), .B2(n109116), .ZN(
        n93654) );
  NAND2_X1 U79204 ( .A1(n93656), .A2(n93657), .ZN(n93601) );
  NOR4_X1 U79205 ( .A1(n93658), .A2(n93659), .A3(n93660), .A4(n93661), .ZN(
        n93657) );
  NAND2_X1 U79206 ( .A1(n93662), .A2(n93663), .ZN(n93661) );
  AOI22_X1 U79207 ( .A1(n90441), .A2(n71992), .B1(n90442), .B2(n109138), .ZN(
        n93663) );
  AOI22_X1 U79208 ( .A1(n90443), .A2(n109142), .B1(n90444), .B2(n109141), .ZN(
        n93662) );
  NAND2_X1 U79209 ( .A1(n93664), .A2(n93665), .ZN(n93660) );
  AOI22_X1 U79210 ( .A1(n90447), .A2(n109147), .B1(n90448), .B2(n109146), .ZN(
        n93665) );
  AOI22_X1 U79211 ( .A1(n90449), .A2(n109137), .B1(n90450), .B2(n109139), .ZN(
        n93664) );
  NAND2_X1 U79212 ( .A1(n93666), .A2(n93667), .ZN(n93659) );
  AOI22_X1 U79213 ( .A1(n90453), .A2(n71997), .B1(n90454), .B2(n109144), .ZN(
        n93667) );
  AOI22_X1 U79214 ( .A1(n90455), .A2(n71996), .B1(n90456), .B2(n71998), .ZN(
        n93666) );
  NAND2_X1 U79215 ( .A1(n93668), .A2(n93669), .ZN(n93658) );
  AOI22_X1 U79216 ( .A1(n90459), .A2(n109150), .B1(n90460), .B2(n72004), .ZN(
        n93669) );
  AOI22_X1 U79217 ( .A1(n90461), .A2(n109143), .B1(n90462), .B2(n109145), .ZN(
        n93668) );
  NOR4_X1 U79218 ( .A1(n93670), .A2(n93671), .A3(n93672), .A4(n93673), .ZN(
        n93656) );
  NAND2_X1 U79219 ( .A1(n93674), .A2(n93675), .ZN(n93673) );
  AOI22_X1 U79220 ( .A1(n90469), .A2(n109126), .B1(n90470), .B2(n109131), .ZN(
        n93675) );
  AOI22_X1 U79221 ( .A1(n90471), .A2(n109125), .B1(n90472), .B2(n71972), .ZN(
        n93674) );
  NAND2_X1 U79222 ( .A1(n93676), .A2(n93677), .ZN(n93672) );
  AOI22_X1 U79223 ( .A1(n90475), .A2(n71981), .B1(n90476), .B2(n109133), .ZN(
        n93677) );
  AOI22_X1 U79224 ( .A1(n90477), .A2(n109134), .B1(n90478), .B2(n109124), .ZN(
        n93676) );
  NAND2_X1 U79225 ( .A1(n93678), .A2(n93679), .ZN(n93671) );
  AOI22_X1 U79226 ( .A1(n90481), .A2(n109132), .B1(n90482), .B2(n109136), .ZN(
        n93679) );
  AOI22_X1 U79227 ( .A1(n90483), .A2(n109130), .B1(n90484), .B2(n109135), .ZN(
        n93678) );
  NAND2_X1 U79228 ( .A1(n93680), .A2(n93681), .ZN(n93670) );
  AOI22_X1 U79229 ( .A1(n90487), .A2(n71986), .B1(n90488), .B2(n109140), .ZN(
        n93681) );
  AOI22_X1 U79230 ( .A1(n90489), .A2(n71984), .B1(n90490), .B2(n109129), .ZN(
        n93680) );
  NAND2_X1 U79231 ( .A1(n93682), .A2(n93683), .ZN(n93600) );
  NOR4_X1 U79232 ( .A1(n93684), .A2(n93685), .A3(n93686), .A4(n93687), .ZN(
        n93683) );
  NAND2_X1 U79233 ( .A1(n93688), .A2(n93689), .ZN(n93687) );
  AOI22_X1 U79234 ( .A1(n90499), .A2(n109168), .B1(n90500), .B2(n109167), .ZN(
        n93689) );
  AOI22_X1 U79235 ( .A1(n90501), .A2(n72020), .B1(n90502), .B2(n109165), .ZN(
        n93688) );
  NAND2_X1 U79236 ( .A1(n93690), .A2(n93691), .ZN(n93686) );
  AOI22_X1 U79237 ( .A1(n90505), .A2(n109163), .B1(n90506), .B2(n109166), .ZN(
        n93691) );
  AOI22_X1 U79238 ( .A1(n105651), .A2(n72026), .B1(n90508), .B2(n109164), .ZN(
        n93690) );
  NAND2_X1 U79239 ( .A1(n93692), .A2(n93693), .ZN(n93685) );
  AOI22_X1 U79240 ( .A1(n90511), .A2(n109174), .B1(n105649), .B2(n72032), .ZN(
        n93693) );
  AOI22_X1 U79241 ( .A1(n105648), .A2(n109172), .B1(n105647), .B2(n109173), 
        .ZN(n93692) );
  NAND2_X1 U79242 ( .A1(n93694), .A2(n93695), .ZN(n93684) );
  AOI22_X1 U79243 ( .A1(n90517), .A2(n109169), .B1(n105646), .B2(n109171), 
        .ZN(n93695) );
  AOI22_X1 U79244 ( .A1(n105645), .A2(n109175), .B1(n105644), .B2(n109170), 
        .ZN(n93694) );
  NOR4_X1 U79245 ( .A1(n93696), .A2(n93697), .A3(n93698), .A4(n93699), .ZN(
        n93682) );
  NAND2_X1 U79246 ( .A1(n93700), .A2(n93701), .ZN(n93699) );
  AOI22_X1 U79247 ( .A1(n90527), .A2(n109149), .B1(n90528), .B2(n109153), .ZN(
        n93701) );
  AOI22_X1 U79248 ( .A1(n90529), .A2(n109152), .B1(n90530), .B2(n72003), .ZN(
        n93700) );
  NAND2_X1 U79249 ( .A1(n93702), .A2(n93703), .ZN(n93698) );
  AOI22_X1 U79250 ( .A1(n90533), .A2(n109159), .B1(n90534), .B2(n109148), .ZN(
        n93703) );
  AOI22_X1 U79251 ( .A1(n90535), .A2(n109151), .B1(n90536), .B2(n109156), .ZN(
        n93702) );
  NAND2_X1 U79252 ( .A1(n93704), .A2(n93705), .ZN(n93697) );
  AOI22_X1 U79253 ( .A1(n90539), .A2(n109155), .B1(n90540), .B2(n109160), .ZN(
        n93705) );
  AOI22_X1 U79254 ( .A1(n90541), .A2(n109162), .B1(n90542), .B2(n109158), .ZN(
        n93704) );
  NAND2_X1 U79255 ( .A1(n93706), .A2(n93707), .ZN(n93696) );
  AOI22_X1 U79256 ( .A1(n90545), .A2(n72021), .B1(n90546), .B2(n109154), .ZN(
        n93707) );
  AOI22_X1 U79257 ( .A1(n90547), .A2(n109157), .B1(n90548), .B2(n109161), .ZN(
        n93706) );
  AOI21_X1 U79258 ( .B1(n90295), .B2(n89742), .A(n93709), .ZN(n93708) );
  OAI21_X1 U79259 ( .B1(n93710), .B2(n90298), .A(n93711), .ZN(n93709) );
  OAI21_X1 U79260 ( .B1(n93712), .B2(n93713), .A(n105658), .ZN(n93711) );
  OAI21_X1 U79261 ( .B1(n101720), .B2(n105657), .A(n93714), .ZN(n93713) );
  AOI22_X1 U79262 ( .A1(n105656), .A2(n108730), .B1(n105655), .B2(n71464), 
        .ZN(n93714) );
  NAND2_X1 U79263 ( .A1(n93715), .A2(n93716), .ZN(n93712) );
  AOI22_X1 U79264 ( .A1(n105654), .A2(n108735), .B1(n90310), .B2(n108732), 
        .ZN(n93716) );
  AOI22_X1 U79265 ( .A1(n90311), .A2(n71462), .B1(n105652), .B2(n108731), .ZN(
        n93715) );
  NOR4_X1 U79266 ( .A1(n93717), .A2(n93718), .A3(n93719), .A4(n93720), .ZN(
        n93710) );
  NAND2_X1 U79267 ( .A1(n93721), .A2(n93722), .ZN(n93720) );
  NOR4_X1 U79268 ( .A1(n93723), .A2(n93724), .A3(n93725), .A4(n93726), .ZN(
        n93722) );
  NAND2_X1 U79269 ( .A1(n93727), .A2(n93728), .ZN(n93726) );
  AOI22_X1 U79270 ( .A1(n90325), .A2(n108711), .B1(n90326), .B2(n108712), .ZN(
        n93728) );
  AOI22_X1 U79271 ( .A1(n90327), .A2(n108720), .B1(n90328), .B2(n108718), .ZN(
        n93727) );
  NAND2_X1 U79272 ( .A1(n93729), .A2(n93730), .ZN(n93725) );
  AOI22_X1 U79273 ( .A1(n90331), .A2(n71331), .B1(n90332), .B2(n108715), .ZN(
        n93730) );
  AOI22_X1 U79274 ( .A1(n90333), .A2(n71435), .B1(n90334), .B2(n108633), .ZN(
        n93729) );
  NAND2_X1 U79275 ( .A1(n93731), .A2(n93732), .ZN(n93724) );
  AOI22_X1 U79276 ( .A1(n90337), .A2(n108637), .B1(n90338), .B2(n71335), .ZN(
        n93732) );
  AOI22_X1 U79277 ( .A1(n90339), .A2(n108716), .B1(n90340), .B2(n108713), .ZN(
        n93731) );
  NAND2_X1 U79278 ( .A1(n93733), .A2(n93734), .ZN(n93723) );
  AOI22_X1 U79279 ( .A1(n90343), .A2(n108635), .B1(n90344), .B2(n108639), .ZN(
        n93734) );
  AOI22_X1 U79280 ( .A1(n90345), .A2(n108638), .B1(n90346), .B2(n71337), .ZN(
        n93733) );
  NOR4_X1 U79281 ( .A1(n93735), .A2(n93736), .A3(n93737), .A4(n93738), .ZN(
        n93721) );
  NAND2_X1 U79282 ( .A1(n93739), .A2(n93740), .ZN(n93738) );
  AOI22_X1 U79283 ( .A1(n90353), .A2(n108721), .B1(n90354), .B2(n108724), .ZN(
        n93740) );
  AOI22_X1 U79284 ( .A1(n90355), .A2(n108725), .B1(n90356), .B2(n108727), .ZN(
        n93739) );
  NAND2_X1 U79285 ( .A1(n93741), .A2(n93742), .ZN(n93737) );
  AOI22_X1 U79286 ( .A1(n90359), .A2(n108726), .B1(n90360), .B2(n108722), .ZN(
        n93742) );
  AOI22_X1 U79287 ( .A1(n90361), .A2(n108728), .B1(n90362), .B2(n108723), .ZN(
        n93741) );
  NAND2_X1 U79288 ( .A1(n93743), .A2(n93744), .ZN(n93736) );
  AOI22_X1 U79289 ( .A1(n90365), .A2(n71445), .B1(n90366), .B2(n71444), .ZN(
        n93744) );
  AOI22_X1 U79290 ( .A1(n90367), .A2(n71447), .B1(n90368), .B2(n108729), .ZN(
        n93743) );
  NAND2_X1 U79291 ( .A1(n93745), .A2(n93746), .ZN(n93735) );
  AOI22_X1 U79292 ( .A1(n90371), .A2(n108714), .B1(n90372), .B2(n108719), .ZN(
        n93746) );
  AOI22_X1 U79293 ( .A1(n90373), .A2(n71442), .B1(n90374), .B2(n108717), .ZN(
        n93745) );
  NAND2_X1 U79294 ( .A1(n93747), .A2(n93748), .ZN(n93719) );
  NOR4_X1 U79295 ( .A1(n93749), .A2(n93750), .A3(n93751), .A4(n93752), .ZN(
        n93748) );
  NAND2_X1 U79296 ( .A1(n93753), .A2(n93754), .ZN(n93752) );
  AOI22_X1 U79297 ( .A1(n90383), .A2(n108648), .B1(n90384), .B2(n108650), .ZN(
        n93754) );
  AOI22_X1 U79298 ( .A1(n90385), .A2(n71360), .B1(n90386), .B2(n108649), .ZN(
        n93753) );
  NAND2_X1 U79299 ( .A1(n93755), .A2(n93756), .ZN(n93751) );
  AOI22_X1 U79300 ( .A1(n90389), .A2(n71364), .B1(n90390), .B2(n71366), .ZN(
        n93756) );
  AOI22_X1 U79301 ( .A1(n90391), .A2(n108656), .B1(n90392), .B2(n108657), .ZN(
        n93755) );
  NAND2_X1 U79302 ( .A1(n93757), .A2(n93758), .ZN(n93750) );
  AOI22_X1 U79303 ( .A1(n90395), .A2(n108653), .B1(n90396), .B2(n108655), .ZN(
        n93758) );
  AOI22_X1 U79304 ( .A1(n90397), .A2(n108658), .B1(n90398), .B2(n108654), .ZN(
        n93757) );
  NAND2_X1 U79305 ( .A1(n93759), .A2(n93760), .ZN(n93749) );
  AOI22_X1 U79306 ( .A1(n90401), .A2(n108663), .B1(n90402), .B2(n71371), .ZN(
        n93760) );
  AOI22_X1 U79307 ( .A1(n90403), .A2(n108662), .B1(n90404), .B2(n71369), .ZN(
        n93759) );
  NOR4_X1 U79308 ( .A1(n93761), .A2(n93762), .A3(n93763), .A4(n93764), .ZN(
        n93747) );
  NAND2_X1 U79309 ( .A1(n93765), .A2(n93766), .ZN(n93764) );
  AOI22_X1 U79310 ( .A1(n90411), .A2(n108643), .B1(n90412), .B2(n108634), .ZN(
        n93766) );
  AOI22_X1 U79311 ( .A1(n90413), .A2(n108636), .B1(n90414), .B2(n71343), .ZN(
        n93765) );
  NAND2_X1 U79312 ( .A1(n93767), .A2(n93768), .ZN(n93763) );
  AOI22_X1 U79313 ( .A1(n90417), .A2(n108641), .B1(n90418), .B2(n108645), .ZN(
        n93768) );
  AOI22_X1 U79314 ( .A1(n90419), .A2(n108647), .B1(n90420), .B2(n108644), .ZN(
        n93767) );
  NAND2_X1 U79315 ( .A1(n93769), .A2(n93770), .ZN(n93762) );
  AOI22_X1 U79316 ( .A1(n90423), .A2(n71352), .B1(n90424), .B2(n108640), .ZN(
        n93770) );
  AOI22_X1 U79317 ( .A1(n90425), .A2(n108642), .B1(n90426), .B2(n108646), .ZN(
        n93769) );
  NAND2_X1 U79318 ( .A1(n93771), .A2(n93772), .ZN(n93761) );
  AOI22_X1 U79319 ( .A1(n90429), .A2(n108652), .B1(n90430), .B2(n71356), .ZN(
        n93772) );
  AOI22_X1 U79320 ( .A1(n90431), .A2(n71354), .B1(n90432), .B2(n108651), .ZN(
        n93771) );
  NAND2_X1 U79321 ( .A1(n93773), .A2(n93774), .ZN(n93718) );
  NOR4_X1 U79322 ( .A1(n93775), .A2(n93776), .A3(n93777), .A4(n93778), .ZN(
        n93774) );
  NAND2_X1 U79323 ( .A1(n93779), .A2(n93780), .ZN(n93778) );
  AOI22_X1 U79324 ( .A1(n90441), .A2(n71394), .B1(n90442), .B2(n108673), .ZN(
        n93780) );
  AOI22_X1 U79325 ( .A1(n90443), .A2(n108677), .B1(n90444), .B2(n108676), .ZN(
        n93779) );
  NAND2_X1 U79326 ( .A1(n93781), .A2(n93782), .ZN(n93777) );
  AOI22_X1 U79327 ( .A1(n90447), .A2(n108682), .B1(n90448), .B2(n108681), .ZN(
        n93782) );
  AOI22_X1 U79328 ( .A1(n90449), .A2(n108672), .B1(n90450), .B2(n108674), .ZN(
        n93781) );
  NAND2_X1 U79329 ( .A1(n93783), .A2(n93784), .ZN(n93776) );
  AOI22_X1 U79330 ( .A1(n90453), .A2(n108683), .B1(n90454), .B2(n108679), .ZN(
        n93784) );
  AOI22_X1 U79331 ( .A1(n90455), .A2(n71398), .B1(n90456), .B2(n71400), .ZN(
        n93783) );
  NAND2_X1 U79332 ( .A1(n93785), .A2(n93786), .ZN(n93775) );
  AOI22_X1 U79333 ( .A1(n90459), .A2(n108686), .B1(n90460), .B2(n71406), .ZN(
        n93786) );
  AOI22_X1 U79334 ( .A1(n90461), .A2(n108678), .B1(n90462), .B2(n108680), .ZN(
        n93785) );
  NOR4_X1 U79335 ( .A1(n93787), .A2(n93788), .A3(n93789), .A4(n93790), .ZN(
        n93773) );
  NAND2_X1 U79336 ( .A1(n93791), .A2(n93792), .ZN(n93790) );
  AOI22_X1 U79337 ( .A1(n90469), .A2(n108661), .B1(n90470), .B2(n108666), .ZN(
        n93792) );
  AOI22_X1 U79338 ( .A1(n90471), .A2(n108660), .B1(n90472), .B2(n71374), .ZN(
        n93791) );
  NAND2_X1 U79339 ( .A1(n93793), .A2(n93794), .ZN(n93789) );
  AOI22_X1 U79340 ( .A1(n90475), .A2(n71383), .B1(n90476), .B2(n108668), .ZN(
        n93794) );
  AOI22_X1 U79341 ( .A1(n90477), .A2(n108669), .B1(n90478), .B2(n108659), .ZN(
        n93793) );
  NAND2_X1 U79342 ( .A1(n93795), .A2(n93796), .ZN(n93788) );
  AOI22_X1 U79343 ( .A1(n90481), .A2(n108667), .B1(n90482), .B2(n108671), .ZN(
        n93796) );
  AOI22_X1 U79344 ( .A1(n90483), .A2(n108665), .B1(n90484), .B2(n108670), .ZN(
        n93795) );
  NAND2_X1 U79345 ( .A1(n93797), .A2(n93798), .ZN(n93787) );
  AOI22_X1 U79346 ( .A1(n90487), .A2(n71388), .B1(n90488), .B2(n108675), .ZN(
        n93798) );
  AOI22_X1 U79347 ( .A1(n90489), .A2(n71386), .B1(n90490), .B2(n108664), .ZN(
        n93797) );
  NAND2_X1 U79348 ( .A1(n93799), .A2(n93800), .ZN(n93717) );
  NOR4_X1 U79349 ( .A1(n93801), .A2(n93802), .A3(n93803), .A4(n93804), .ZN(
        n93800) );
  NAND2_X1 U79350 ( .A1(n93805), .A2(n93806), .ZN(n93804) );
  AOI22_X1 U79351 ( .A1(n90499), .A2(n108704), .B1(n90500), .B2(n108703), .ZN(
        n93806) );
  AOI22_X1 U79352 ( .A1(n90501), .A2(n71422), .B1(n90502), .B2(n108701), .ZN(
        n93805) );
  NAND2_X1 U79353 ( .A1(n93807), .A2(n93808), .ZN(n93803) );
  AOI22_X1 U79354 ( .A1(n90505), .A2(n108699), .B1(n90506), .B2(n108702), .ZN(
        n93808) );
  AOI22_X1 U79355 ( .A1(n105651), .A2(n71428), .B1(n90508), .B2(n108700), .ZN(
        n93807) );
  NAND2_X1 U79356 ( .A1(n93809), .A2(n93810), .ZN(n93802) );
  AOI22_X1 U79357 ( .A1(n90511), .A2(n108709), .B1(n105649), .B2(n71434), .ZN(
        n93810) );
  AOI22_X1 U79358 ( .A1(n105648), .A2(n108707), .B1(n105647), .B2(n108708), 
        .ZN(n93809) );
  NAND2_X1 U79359 ( .A1(n93811), .A2(n93812), .ZN(n93801) );
  AOI22_X1 U79360 ( .A1(n90517), .A2(n108705), .B1(n105646), .B2(n71429), .ZN(
        n93812) );
  AOI22_X1 U79361 ( .A1(n105645), .A2(n108710), .B1(n105644), .B2(n108706), 
        .ZN(n93811) );
  NOR4_X1 U79362 ( .A1(n93813), .A2(n93814), .A3(n93815), .A4(n93816), .ZN(
        n93799) );
  NAND2_X1 U79363 ( .A1(n93817), .A2(n93818), .ZN(n93816) );
  AOI22_X1 U79364 ( .A1(n90527), .A2(n108685), .B1(n90528), .B2(n108689), .ZN(
        n93818) );
  AOI22_X1 U79365 ( .A1(n90529), .A2(n108688), .B1(n90530), .B2(n71405), .ZN(
        n93817) );
  NAND2_X1 U79366 ( .A1(n93819), .A2(n93820), .ZN(n93815) );
  AOI22_X1 U79367 ( .A1(n90533), .A2(n108695), .B1(n90534), .B2(n108684), .ZN(
        n93820) );
  AOI22_X1 U79368 ( .A1(n90535), .A2(n108687), .B1(n90536), .B2(n108692), .ZN(
        n93819) );
  NAND2_X1 U79369 ( .A1(n93821), .A2(n93822), .ZN(n93814) );
  AOI22_X1 U79370 ( .A1(n90539), .A2(n108691), .B1(n90540), .B2(n108696), .ZN(
        n93822) );
  AOI22_X1 U79371 ( .A1(n90541), .A2(n108698), .B1(n90542), .B2(n108694), .ZN(
        n93821) );
  NAND2_X1 U79372 ( .A1(n93823), .A2(n93824), .ZN(n93813) );
  AOI22_X1 U79373 ( .A1(n90545), .A2(n71423), .B1(n90546), .B2(n108690), .ZN(
        n93824) );
  AOI22_X1 U79374 ( .A1(n90547), .A2(n108693), .B1(n90548), .B2(n108697), .ZN(
        n93823) );
  AOI21_X1 U79375 ( .B1(n90295), .B2(n81790), .A(n93826), .ZN(n93825) );
  OAI21_X1 U79376 ( .B1(n93827), .B2(n105659), .A(n93828), .ZN(n93826) );
  OAI21_X1 U79377 ( .B1(n93829), .B2(n93830), .A(n105658), .ZN(n93828) );
  OAI21_X1 U79378 ( .B1(n101702), .B2(n105657), .A(n93831), .ZN(n93830) );
  AOI22_X1 U79379 ( .A1(n105656), .A2(n108958), .B1(n105655), .B2(n71759), 
        .ZN(n93831) );
  NAND2_X1 U79380 ( .A1(n93832), .A2(n93833), .ZN(n93829) );
  AOI22_X1 U79381 ( .A1(n105654), .A2(n108963), .B1(n90310), .B2(n108960), 
        .ZN(n93833) );
  AOI22_X1 U79382 ( .A1(n90311), .A2(n71757), .B1(n105652), .B2(n108959), .ZN(
        n93832) );
  NOR4_X1 U79383 ( .A1(n93834), .A2(n93835), .A3(n93836), .A4(n93837), .ZN(
        n93827) );
  NAND2_X1 U79384 ( .A1(n93838), .A2(n93839), .ZN(n93837) );
  NOR4_X1 U79385 ( .A1(n93840), .A2(n93841), .A3(n93842), .A4(n93843), .ZN(
        n93839) );
  NAND2_X1 U79386 ( .A1(n93844), .A2(n93845), .ZN(n93843) );
  AOI22_X1 U79387 ( .A1(n90325), .A2(n108939), .B1(n90326), .B2(n108940), .ZN(
        n93845) );
  AOI22_X1 U79388 ( .A1(n90327), .A2(n108948), .B1(n90328), .B2(n108946), .ZN(
        n93844) );
  NAND2_X1 U79389 ( .A1(n93846), .A2(n93847), .ZN(n93842) );
  AOI22_X1 U79390 ( .A1(n90331), .A2(n71626), .B1(n90332), .B2(n108943), .ZN(
        n93847) );
  AOI22_X1 U79391 ( .A1(n90333), .A2(n71730), .B1(n90334), .B2(n108860), .ZN(
        n93846) );
  NAND2_X1 U79392 ( .A1(n93848), .A2(n93849), .ZN(n93841) );
  AOI22_X1 U79393 ( .A1(n90337), .A2(n108864), .B1(n90338), .B2(n71630), .ZN(
        n93849) );
  AOI22_X1 U79394 ( .A1(n90339), .A2(n108944), .B1(n90340), .B2(n108941), .ZN(
        n93848) );
  NAND2_X1 U79395 ( .A1(n93850), .A2(n93851), .ZN(n93840) );
  AOI22_X1 U79396 ( .A1(n90343), .A2(n108862), .B1(n90344), .B2(n108866), .ZN(
        n93851) );
  AOI22_X1 U79397 ( .A1(n90345), .A2(n108865), .B1(n90346), .B2(n71632), .ZN(
        n93850) );
  NOR4_X1 U79398 ( .A1(n93852), .A2(n93853), .A3(n93854), .A4(n93855), .ZN(
        n93838) );
  NAND2_X1 U79399 ( .A1(n93856), .A2(n93857), .ZN(n93855) );
  AOI22_X1 U79400 ( .A1(n90353), .A2(n108949), .B1(n90354), .B2(n108952), .ZN(
        n93857) );
  AOI22_X1 U79401 ( .A1(n90355), .A2(n108953), .B1(n90356), .B2(n108955), .ZN(
        n93856) );
  NAND2_X1 U79402 ( .A1(n93858), .A2(n93859), .ZN(n93854) );
  AOI22_X1 U79403 ( .A1(n90359), .A2(n108954), .B1(n90360), .B2(n108950), .ZN(
        n93859) );
  AOI22_X1 U79404 ( .A1(n90361), .A2(n108956), .B1(n90362), .B2(n108951), .ZN(
        n93858) );
  NAND2_X1 U79405 ( .A1(n93860), .A2(n93861), .ZN(n93853) );
  AOI22_X1 U79406 ( .A1(n90365), .A2(n71740), .B1(n90366), .B2(n71739), .ZN(
        n93861) );
  AOI22_X1 U79407 ( .A1(n90367), .A2(n71742), .B1(n90368), .B2(n108957), .ZN(
        n93860) );
  NAND2_X1 U79408 ( .A1(n93862), .A2(n93863), .ZN(n93852) );
  AOI22_X1 U79409 ( .A1(n90371), .A2(n108942), .B1(n90372), .B2(n108947), .ZN(
        n93863) );
  AOI22_X1 U79410 ( .A1(n90373), .A2(n71737), .B1(n90374), .B2(n108945), .ZN(
        n93862) );
  NAND2_X1 U79411 ( .A1(n93864), .A2(n93865), .ZN(n93836) );
  NOR4_X1 U79412 ( .A1(n93866), .A2(n93867), .A3(n93868), .A4(n93869), .ZN(
        n93865) );
  NAND2_X1 U79413 ( .A1(n93870), .A2(n93871), .ZN(n93869) );
  AOI22_X1 U79414 ( .A1(n90383), .A2(n108875), .B1(n90384), .B2(n108877), .ZN(
        n93871) );
  AOI22_X1 U79415 ( .A1(n90385), .A2(n71655), .B1(n90386), .B2(n108876), .ZN(
        n93870) );
  NAND2_X1 U79416 ( .A1(n93872), .A2(n93873), .ZN(n93868) );
  AOI22_X1 U79417 ( .A1(n90389), .A2(n71659), .B1(n90390), .B2(n71661), .ZN(
        n93873) );
  AOI22_X1 U79418 ( .A1(n90391), .A2(n108883), .B1(n90392), .B2(n108884), .ZN(
        n93872) );
  NAND2_X1 U79419 ( .A1(n93874), .A2(n93875), .ZN(n93867) );
  AOI22_X1 U79420 ( .A1(n90395), .A2(n108880), .B1(n90396), .B2(n108882), .ZN(
        n93875) );
  AOI22_X1 U79421 ( .A1(n90397), .A2(n108885), .B1(n90398), .B2(n108881), .ZN(
        n93874) );
  NAND2_X1 U79422 ( .A1(n93876), .A2(n93877), .ZN(n93866) );
  AOI22_X1 U79423 ( .A1(n90401), .A2(n108890), .B1(n90402), .B2(n71666), .ZN(
        n93877) );
  AOI22_X1 U79424 ( .A1(n90403), .A2(n108889), .B1(n90404), .B2(n71664), .ZN(
        n93876) );
  NOR4_X1 U79425 ( .A1(n93878), .A2(n93879), .A3(n93880), .A4(n93881), .ZN(
        n93864) );
  NAND2_X1 U79426 ( .A1(n93882), .A2(n93883), .ZN(n93881) );
  AOI22_X1 U79427 ( .A1(n90411), .A2(n108870), .B1(n90412), .B2(n108861), .ZN(
        n93883) );
  AOI22_X1 U79428 ( .A1(n90413), .A2(n108863), .B1(n90414), .B2(n71638), .ZN(
        n93882) );
  NAND2_X1 U79429 ( .A1(n93884), .A2(n93885), .ZN(n93880) );
  AOI22_X1 U79430 ( .A1(n90417), .A2(n108868), .B1(n90418), .B2(n108872), .ZN(
        n93885) );
  AOI22_X1 U79431 ( .A1(n90419), .A2(n108874), .B1(n90420), .B2(n108871), .ZN(
        n93884) );
  NAND2_X1 U79432 ( .A1(n93886), .A2(n93887), .ZN(n93879) );
  AOI22_X1 U79433 ( .A1(n90423), .A2(n71647), .B1(n90424), .B2(n108867), .ZN(
        n93887) );
  AOI22_X1 U79434 ( .A1(n90425), .A2(n108869), .B1(n90426), .B2(n108873), .ZN(
        n93886) );
  NAND2_X1 U79435 ( .A1(n93888), .A2(n93889), .ZN(n93878) );
  AOI22_X1 U79436 ( .A1(n90429), .A2(n108879), .B1(n90430), .B2(n71651), .ZN(
        n93889) );
  AOI22_X1 U79437 ( .A1(n90431), .A2(n71649), .B1(n90432), .B2(n108878), .ZN(
        n93888) );
  NAND2_X1 U79438 ( .A1(n93890), .A2(n93891), .ZN(n93835) );
  NOR4_X1 U79439 ( .A1(n93892), .A2(n93893), .A3(n93894), .A4(n93895), .ZN(
        n93891) );
  NAND2_X1 U79440 ( .A1(n93896), .A2(n93897), .ZN(n93895) );
  AOI22_X1 U79441 ( .A1(n90441), .A2(n71689), .B1(n90442), .B2(n108900), .ZN(
        n93897) );
  AOI22_X1 U79442 ( .A1(n90443), .A2(n108904), .B1(n90444), .B2(n108903), .ZN(
        n93896) );
  NAND2_X1 U79443 ( .A1(n93898), .A2(n93899), .ZN(n93894) );
  AOI22_X1 U79444 ( .A1(n90447), .A2(n108909), .B1(n90448), .B2(n108908), .ZN(
        n93899) );
  AOI22_X1 U79445 ( .A1(n90449), .A2(n108899), .B1(n90450), .B2(n108901), .ZN(
        n93898) );
  NAND2_X1 U79446 ( .A1(n93900), .A2(n93901), .ZN(n93893) );
  AOI22_X1 U79447 ( .A1(n90453), .A2(n108910), .B1(n90454), .B2(n108906), .ZN(
        n93901) );
  AOI22_X1 U79448 ( .A1(n90455), .A2(n71693), .B1(n90456), .B2(n71695), .ZN(
        n93900) );
  NAND2_X1 U79449 ( .A1(n93902), .A2(n93903), .ZN(n93892) );
  AOI22_X1 U79450 ( .A1(n90459), .A2(n108913), .B1(n90460), .B2(n71701), .ZN(
        n93903) );
  AOI22_X1 U79451 ( .A1(n90461), .A2(n108905), .B1(n90462), .B2(n108907), .ZN(
        n93902) );
  NOR4_X1 U79452 ( .A1(n93904), .A2(n93905), .A3(n93906), .A4(n93907), .ZN(
        n93890) );
  NAND2_X1 U79453 ( .A1(n93908), .A2(n93909), .ZN(n93907) );
  AOI22_X1 U79454 ( .A1(n90469), .A2(n108888), .B1(n90470), .B2(n108893), .ZN(
        n93909) );
  AOI22_X1 U79455 ( .A1(n90471), .A2(n108887), .B1(n90472), .B2(n71669), .ZN(
        n93908) );
  NAND2_X1 U79456 ( .A1(n93910), .A2(n93911), .ZN(n93906) );
  AOI22_X1 U79457 ( .A1(n90475), .A2(n71678), .B1(n90476), .B2(n108895), .ZN(
        n93911) );
  AOI22_X1 U79458 ( .A1(n90477), .A2(n108896), .B1(n90478), .B2(n108886), .ZN(
        n93910) );
  NAND2_X1 U79459 ( .A1(n93912), .A2(n93913), .ZN(n93905) );
  AOI22_X1 U79460 ( .A1(n90481), .A2(n108894), .B1(n90482), .B2(n108898), .ZN(
        n93913) );
  AOI22_X1 U79461 ( .A1(n90483), .A2(n108892), .B1(n90484), .B2(n108897), .ZN(
        n93912) );
  NAND2_X1 U79462 ( .A1(n93914), .A2(n93915), .ZN(n93904) );
  AOI22_X1 U79463 ( .A1(n90487), .A2(n71683), .B1(n90488), .B2(n108902), .ZN(
        n93915) );
  AOI22_X1 U79464 ( .A1(n90489), .A2(n71681), .B1(n90490), .B2(n108891), .ZN(
        n93914) );
  NAND2_X1 U79465 ( .A1(n93916), .A2(n93917), .ZN(n93834) );
  NOR4_X1 U79466 ( .A1(n93918), .A2(n93919), .A3(n93920), .A4(n93921), .ZN(
        n93917) );
  NAND2_X1 U79467 ( .A1(n93922), .A2(n93923), .ZN(n93921) );
  AOI22_X1 U79468 ( .A1(n90499), .A2(n108931), .B1(n90500), .B2(n108930), .ZN(
        n93923) );
  AOI22_X1 U79469 ( .A1(n90501), .A2(n71717), .B1(n90502), .B2(n108928), .ZN(
        n93922) );
  NAND2_X1 U79470 ( .A1(n93924), .A2(n93925), .ZN(n93920) );
  AOI22_X1 U79471 ( .A1(n90505), .A2(n108926), .B1(n90506), .B2(n108929), .ZN(
        n93925) );
  AOI22_X1 U79472 ( .A1(n105651), .A2(n71723), .B1(n90508), .B2(n108927), .ZN(
        n93924) );
  NAND2_X1 U79473 ( .A1(n93926), .A2(n93927), .ZN(n93919) );
  AOI22_X1 U79474 ( .A1(n90511), .A2(n108937), .B1(n105649), .B2(n71729), .ZN(
        n93927) );
  AOI22_X1 U79475 ( .A1(n105648), .A2(n108935), .B1(n105647), .B2(n108936), 
        .ZN(n93926) );
  NAND2_X1 U79476 ( .A1(n93928), .A2(n93929), .ZN(n93918) );
  AOI22_X1 U79477 ( .A1(n90517), .A2(n108932), .B1(n105646), .B2(n108934), 
        .ZN(n93929) );
  AOI22_X1 U79478 ( .A1(n105645), .A2(n108938), .B1(n105644), .B2(n108933), 
        .ZN(n93928) );
  NOR4_X1 U79479 ( .A1(n93930), .A2(n93931), .A3(n93932), .A4(n93933), .ZN(
        n93916) );
  NAND2_X1 U79480 ( .A1(n93934), .A2(n93935), .ZN(n93933) );
  AOI22_X1 U79481 ( .A1(n90527), .A2(n108912), .B1(n90528), .B2(n108916), .ZN(
        n93935) );
  AOI22_X1 U79482 ( .A1(n90529), .A2(n108915), .B1(n90530), .B2(n71700), .ZN(
        n93934) );
  NAND2_X1 U79483 ( .A1(n93936), .A2(n93937), .ZN(n93932) );
  AOI22_X1 U79484 ( .A1(n90533), .A2(n108922), .B1(n90534), .B2(n108911), .ZN(
        n93937) );
  AOI22_X1 U79485 ( .A1(n90535), .A2(n108914), .B1(n90536), .B2(n108919), .ZN(
        n93936) );
  NAND2_X1 U79486 ( .A1(n93938), .A2(n93939), .ZN(n93931) );
  AOI22_X1 U79487 ( .A1(n90539), .A2(n108918), .B1(n90540), .B2(n108923), .ZN(
        n93939) );
  AOI22_X1 U79488 ( .A1(n90541), .A2(n108925), .B1(n90542), .B2(n108921), .ZN(
        n93938) );
  NAND2_X1 U79489 ( .A1(n93940), .A2(n93941), .ZN(n93930) );
  AOI22_X1 U79490 ( .A1(n90545), .A2(n71718), .B1(n90546), .B2(n108917), .ZN(
        n93941) );
  AOI22_X1 U79491 ( .A1(n90547), .A2(n108920), .B1(n90548), .B2(n108924), .ZN(
        n93940) );
  AOI21_X1 U79492 ( .B1(n90295), .B2(n89977), .A(n93943), .ZN(n93942) );
  OAI21_X1 U79493 ( .B1(n93944), .B2(n90298), .A(n93945), .ZN(n93943) );
  OAI21_X1 U79494 ( .B1(n93946), .B2(n93947), .A(n105658), .ZN(n93945) );
  OAI21_X1 U79495 ( .B1(n101684), .B2(n105657), .A(n93948), .ZN(n93947) );
  AOI22_X1 U79496 ( .A1(n105656), .A2(n108846), .B1(n105655), .B2(n71615), 
        .ZN(n93948) );
  NAND2_X1 U79497 ( .A1(n93949), .A2(n93950), .ZN(n93946) );
  AOI22_X1 U79498 ( .A1(n105654), .A2(n108851), .B1(n90310), .B2(n108848), 
        .ZN(n93950) );
  AOI22_X1 U79499 ( .A1(n90311), .A2(n71613), .B1(n105652), .B2(n108847), .ZN(
        n93949) );
  NOR4_X1 U79500 ( .A1(n93951), .A2(n93952), .A3(n93953), .A4(n93954), .ZN(
        n93944) );
  NAND2_X1 U79501 ( .A1(n93955), .A2(n93956), .ZN(n93954) );
  NOR4_X1 U79502 ( .A1(n93957), .A2(n93958), .A3(n93959), .A4(n93960), .ZN(
        n93956) );
  NAND2_X1 U79503 ( .A1(n93961), .A2(n93962), .ZN(n93960) );
  AOI22_X1 U79504 ( .A1(n90325), .A2(n108827), .B1(n90326), .B2(n108828), .ZN(
        n93962) );
  AOI22_X1 U79505 ( .A1(n90327), .A2(n108836), .B1(n90328), .B2(n108834), .ZN(
        n93961) );
  NAND2_X1 U79506 ( .A1(n93963), .A2(n93964), .ZN(n93959) );
  AOI22_X1 U79507 ( .A1(n90331), .A2(n71482), .B1(n90332), .B2(n108831), .ZN(
        n93964) );
  AOI22_X1 U79508 ( .A1(n90333), .A2(n71586), .B1(n90334), .B2(n108748), .ZN(
        n93963) );
  NAND2_X1 U79509 ( .A1(n93965), .A2(n93966), .ZN(n93958) );
  AOI22_X1 U79510 ( .A1(n90337), .A2(n108752), .B1(n90338), .B2(n71486), .ZN(
        n93966) );
  AOI22_X1 U79511 ( .A1(n90339), .A2(n108832), .B1(n90340), .B2(n108829), .ZN(
        n93965) );
  NAND2_X1 U79512 ( .A1(n93967), .A2(n93968), .ZN(n93957) );
  AOI22_X1 U79513 ( .A1(n90343), .A2(n108750), .B1(n90344), .B2(n108754), .ZN(
        n93968) );
  AOI22_X1 U79514 ( .A1(n90345), .A2(n108753), .B1(n90346), .B2(n71488), .ZN(
        n93967) );
  NOR4_X1 U79515 ( .A1(n93969), .A2(n93970), .A3(n93971), .A4(n93972), .ZN(
        n93955) );
  NAND2_X1 U79516 ( .A1(n93973), .A2(n93974), .ZN(n93972) );
  AOI22_X1 U79517 ( .A1(n90353), .A2(n108837), .B1(n90354), .B2(n108840), .ZN(
        n93974) );
  AOI22_X1 U79518 ( .A1(n90355), .A2(n108841), .B1(n90356), .B2(n108843), .ZN(
        n93973) );
  NAND2_X1 U79519 ( .A1(n93975), .A2(n93976), .ZN(n93971) );
  AOI22_X1 U79520 ( .A1(n90359), .A2(n108842), .B1(n90360), .B2(n108838), .ZN(
        n93976) );
  AOI22_X1 U79521 ( .A1(n90361), .A2(n108844), .B1(n90362), .B2(n108839), .ZN(
        n93975) );
  NAND2_X1 U79522 ( .A1(n93977), .A2(n93978), .ZN(n93970) );
  AOI22_X1 U79523 ( .A1(n90365), .A2(n71596), .B1(n90366), .B2(n71595), .ZN(
        n93978) );
  AOI22_X1 U79524 ( .A1(n90367), .A2(n71598), .B1(n90368), .B2(n108845), .ZN(
        n93977) );
  NAND2_X1 U79525 ( .A1(n93979), .A2(n93980), .ZN(n93969) );
  AOI22_X1 U79526 ( .A1(n90371), .A2(n108830), .B1(n90372), .B2(n108835), .ZN(
        n93980) );
  AOI22_X1 U79527 ( .A1(n90373), .A2(n71593), .B1(n90374), .B2(n108833), .ZN(
        n93979) );
  NAND2_X1 U79528 ( .A1(n93981), .A2(n93982), .ZN(n93953) );
  NOR4_X1 U79529 ( .A1(n93983), .A2(n93984), .A3(n93985), .A4(n93986), .ZN(
        n93982) );
  NAND2_X1 U79530 ( .A1(n93987), .A2(n93988), .ZN(n93986) );
  AOI22_X1 U79531 ( .A1(n90383), .A2(n108763), .B1(n90384), .B2(n108765), .ZN(
        n93988) );
  AOI22_X1 U79532 ( .A1(n90385), .A2(n71511), .B1(n90386), .B2(n108764), .ZN(
        n93987) );
  NAND2_X1 U79533 ( .A1(n93989), .A2(n93990), .ZN(n93985) );
  AOI22_X1 U79534 ( .A1(n90389), .A2(n71515), .B1(n90390), .B2(n71517), .ZN(
        n93990) );
  AOI22_X1 U79535 ( .A1(n90391), .A2(n108771), .B1(n90392), .B2(n108772), .ZN(
        n93989) );
  NAND2_X1 U79536 ( .A1(n93991), .A2(n93992), .ZN(n93984) );
  AOI22_X1 U79537 ( .A1(n90395), .A2(n108768), .B1(n90396), .B2(n108770), .ZN(
        n93992) );
  AOI22_X1 U79538 ( .A1(n90397), .A2(n108773), .B1(n90398), .B2(n108769), .ZN(
        n93991) );
  NAND2_X1 U79539 ( .A1(n93993), .A2(n93994), .ZN(n93983) );
  AOI22_X1 U79540 ( .A1(n90401), .A2(n108778), .B1(n90402), .B2(n71522), .ZN(
        n93994) );
  AOI22_X1 U79541 ( .A1(n90403), .A2(n108777), .B1(n90404), .B2(n71520), .ZN(
        n93993) );
  NOR4_X1 U79542 ( .A1(n93995), .A2(n93996), .A3(n93997), .A4(n93998), .ZN(
        n93981) );
  NAND2_X1 U79543 ( .A1(n93999), .A2(n94000), .ZN(n93998) );
  AOI22_X1 U79544 ( .A1(n90411), .A2(n108758), .B1(n90412), .B2(n108749), .ZN(
        n94000) );
  AOI22_X1 U79545 ( .A1(n90413), .A2(n108751), .B1(n90414), .B2(n71494), .ZN(
        n93999) );
  NAND2_X1 U79546 ( .A1(n94001), .A2(n94002), .ZN(n93997) );
  AOI22_X1 U79547 ( .A1(n90417), .A2(n108756), .B1(n90418), .B2(n108760), .ZN(
        n94002) );
  AOI22_X1 U79548 ( .A1(n90419), .A2(n108762), .B1(n90420), .B2(n108759), .ZN(
        n94001) );
  NAND2_X1 U79549 ( .A1(n94003), .A2(n94004), .ZN(n93996) );
  AOI22_X1 U79550 ( .A1(n90423), .A2(n71503), .B1(n90424), .B2(n108755), .ZN(
        n94004) );
  AOI22_X1 U79551 ( .A1(n90425), .A2(n108757), .B1(n90426), .B2(n108761), .ZN(
        n94003) );
  NAND2_X1 U79552 ( .A1(n94005), .A2(n94006), .ZN(n93995) );
  AOI22_X1 U79553 ( .A1(n90429), .A2(n108767), .B1(n90430), .B2(n71507), .ZN(
        n94006) );
  AOI22_X1 U79554 ( .A1(n90431), .A2(n71505), .B1(n90432), .B2(n108766), .ZN(
        n94005) );
  NAND2_X1 U79555 ( .A1(n94007), .A2(n94008), .ZN(n93952) );
  NOR4_X1 U79556 ( .A1(n94009), .A2(n94010), .A3(n94011), .A4(n94012), .ZN(
        n94008) );
  NAND2_X1 U79557 ( .A1(n94013), .A2(n94014), .ZN(n94012) );
  AOI22_X1 U79558 ( .A1(n90441), .A2(n71545), .B1(n90442), .B2(n108788), .ZN(
        n94014) );
  AOI22_X1 U79559 ( .A1(n90443), .A2(n108792), .B1(n90444), .B2(n108791), .ZN(
        n94013) );
  NAND2_X1 U79560 ( .A1(n94015), .A2(n94016), .ZN(n94011) );
  AOI22_X1 U79561 ( .A1(n90447), .A2(n108797), .B1(n90448), .B2(n108796), .ZN(
        n94016) );
  AOI22_X1 U79562 ( .A1(n90449), .A2(n108787), .B1(n90450), .B2(n108789), .ZN(
        n94015) );
  NAND2_X1 U79563 ( .A1(n94017), .A2(n94018), .ZN(n94010) );
  AOI22_X1 U79564 ( .A1(n90453), .A2(n108798), .B1(n90454), .B2(n108794), .ZN(
        n94018) );
  AOI22_X1 U79565 ( .A1(n90455), .A2(n71549), .B1(n90456), .B2(n71551), .ZN(
        n94017) );
  NAND2_X1 U79566 ( .A1(n94019), .A2(n94020), .ZN(n94009) );
  AOI22_X1 U79567 ( .A1(n90459), .A2(n108801), .B1(n90460), .B2(n71557), .ZN(
        n94020) );
  AOI22_X1 U79568 ( .A1(n90461), .A2(n108793), .B1(n90462), .B2(n108795), .ZN(
        n94019) );
  NOR4_X1 U79569 ( .A1(n94021), .A2(n94022), .A3(n94023), .A4(n94024), .ZN(
        n94007) );
  NAND2_X1 U79570 ( .A1(n94025), .A2(n94026), .ZN(n94024) );
  AOI22_X1 U79571 ( .A1(n90469), .A2(n108776), .B1(n90470), .B2(n108781), .ZN(
        n94026) );
  AOI22_X1 U79572 ( .A1(n90471), .A2(n108775), .B1(n90472), .B2(n71525), .ZN(
        n94025) );
  NAND2_X1 U79573 ( .A1(n94027), .A2(n94028), .ZN(n94023) );
  AOI22_X1 U79574 ( .A1(n90475), .A2(n71534), .B1(n90476), .B2(n108783), .ZN(
        n94028) );
  AOI22_X1 U79575 ( .A1(n90477), .A2(n108784), .B1(n90478), .B2(n108774), .ZN(
        n94027) );
  NAND2_X1 U79576 ( .A1(n94029), .A2(n94030), .ZN(n94022) );
  AOI22_X1 U79577 ( .A1(n90481), .A2(n108782), .B1(n90482), .B2(n108786), .ZN(
        n94030) );
  AOI22_X1 U79578 ( .A1(n90483), .A2(n108780), .B1(n90484), .B2(n108785), .ZN(
        n94029) );
  NAND2_X1 U79579 ( .A1(n94031), .A2(n94032), .ZN(n94021) );
  AOI22_X1 U79580 ( .A1(n90487), .A2(n71539), .B1(n90488), .B2(n108790), .ZN(
        n94032) );
  AOI22_X1 U79581 ( .A1(n90489), .A2(n71537), .B1(n90490), .B2(n108779), .ZN(
        n94031) );
  NAND2_X1 U79582 ( .A1(n94033), .A2(n94034), .ZN(n93951) );
  NOR4_X1 U79583 ( .A1(n94035), .A2(n94036), .A3(n94037), .A4(n94038), .ZN(
        n94034) );
  NAND2_X1 U79584 ( .A1(n94039), .A2(n94040), .ZN(n94038) );
  AOI22_X1 U79585 ( .A1(n90499), .A2(n108819), .B1(n90500), .B2(n108818), .ZN(
        n94040) );
  AOI22_X1 U79586 ( .A1(n90501), .A2(n71573), .B1(n90502), .B2(n108816), .ZN(
        n94039) );
  NAND2_X1 U79587 ( .A1(n94041), .A2(n94042), .ZN(n94037) );
  AOI22_X1 U79588 ( .A1(n90505), .A2(n108814), .B1(n90506), .B2(n108817), .ZN(
        n94042) );
  AOI22_X1 U79589 ( .A1(n105651), .A2(n71579), .B1(n90508), .B2(n108815), .ZN(
        n94041) );
  NAND2_X1 U79590 ( .A1(n94043), .A2(n94044), .ZN(n94036) );
  AOI22_X1 U79591 ( .A1(n90511), .A2(n108825), .B1(n105649), .B2(n71585), .ZN(
        n94044) );
  AOI22_X1 U79592 ( .A1(n105648), .A2(n108823), .B1(n105647), .B2(n108824), 
        .ZN(n94043) );
  NAND2_X1 U79593 ( .A1(n94045), .A2(n94046), .ZN(n94035) );
  AOI22_X1 U79594 ( .A1(n90517), .A2(n108820), .B1(n105646), .B2(n108822), 
        .ZN(n94046) );
  AOI22_X1 U79595 ( .A1(n105645), .A2(n108826), .B1(n105644), .B2(n108821), 
        .ZN(n94045) );
  NOR4_X1 U79596 ( .A1(n94047), .A2(n94048), .A3(n94049), .A4(n94050), .ZN(
        n94033) );
  NAND2_X1 U79597 ( .A1(n94051), .A2(n94052), .ZN(n94050) );
  AOI22_X1 U79598 ( .A1(n90527), .A2(n108800), .B1(n90528), .B2(n108804), .ZN(
        n94052) );
  AOI22_X1 U79599 ( .A1(n90529), .A2(n108803), .B1(n90530), .B2(n71556), .ZN(
        n94051) );
  NAND2_X1 U79600 ( .A1(n94053), .A2(n94054), .ZN(n94049) );
  AOI22_X1 U79601 ( .A1(n90533), .A2(n108810), .B1(n90534), .B2(n108799), .ZN(
        n94054) );
  AOI22_X1 U79602 ( .A1(n90535), .A2(n108802), .B1(n90536), .B2(n108807), .ZN(
        n94053) );
  NAND2_X1 U79603 ( .A1(n94055), .A2(n94056), .ZN(n94048) );
  AOI22_X1 U79604 ( .A1(n90539), .A2(n108806), .B1(n90540), .B2(n108811), .ZN(
        n94056) );
  AOI22_X1 U79605 ( .A1(n90541), .A2(n108813), .B1(n90542), .B2(n108809), .ZN(
        n94055) );
  NAND2_X1 U79606 ( .A1(n94057), .A2(n94058), .ZN(n94047) );
  AOI22_X1 U79607 ( .A1(n90545), .A2(n71574), .B1(n90546), .B2(n108805), .ZN(
        n94058) );
  AOI22_X1 U79608 ( .A1(n90547), .A2(n108808), .B1(n90548), .B2(n108812), .ZN(
        n94057) );
  OAI21_X1 U79609 ( .B1(n94059), .B2(n105659), .A(n94060), .ZN(
        \DLX_Datapath/RegisterFile/N46424 ) );
  AOI22_X1 U79610 ( .A1(n105658), .A2(n94061), .B1(n90295), .B2(n90096), .ZN(
        n94060) );
  AND2_X2 U79611 ( .A1(n94062), .A2(n94063), .ZN(n90295) );
  AOI22_X1 U79612 ( .A1(n104705), .A2(n107118), .B1(n94064), .B2(n107146), 
        .ZN(n94063) );
  AOI21_X1 U79613 ( .B1(n94067), .B2(n94068), .A(n111056), .ZN(n94062) );
  OR2_X1 U79614 ( .A1(n94069), .A2(n94070), .ZN(n94061) );
  OAI21_X1 U79615 ( .B1(n101666), .B2(n105657), .A(n94071), .ZN(n94070) );
  AOI22_X1 U79616 ( .A1(n105656), .A2(n107175), .B1(n105655), .B2(n69426), 
        .ZN(n94071) );
  NOR2_X1 U79617 ( .A1(n94072), .A2(n94065), .ZN(n90306) );
  NOR2_X1 U79618 ( .A1(n94073), .A2(n59452), .ZN(n90305) );
  OR2_X1 U79619 ( .A1(n94073), .A2(n94065), .ZN(n90303) );
  NAND2_X1 U79620 ( .A1(n107144), .A2(n107145), .ZN(n94073) );
  NAND2_X1 U79621 ( .A1(n94074), .A2(n94075), .ZN(n94069) );
  AOI22_X1 U79622 ( .A1(n105654), .A2(n106767), .B1(n90310), .B2(n107171), 
        .ZN(n94075) );
  NOR2_X1 U79623 ( .A1(n94076), .A2(n59452), .ZN(n90310) );
  NOR2_X1 U79624 ( .A1(n94065), .A2(n94076), .ZN(n90309) );
  NAND2_X1 U79625 ( .A1(n59451), .A2(n107144), .ZN(n94076) );
  NAND2_X1 U79626 ( .A1(n104705), .A2(n59452), .ZN(n94065) );
  AOI22_X1 U79627 ( .A1(n90311), .A2(n69430), .B1(n105652), .B2(n107173), .ZN(
        n94074) );
  NOR2_X1 U79628 ( .A1(n94072), .A2(n59452), .ZN(n90312) );
  NAND2_X1 U79629 ( .A1(n59445), .A2(n107145), .ZN(n94072) );
  AND2_X2 U79630 ( .A1(n94064), .A2(n105061), .ZN(n90311) );
  NOR2_X1 U79631 ( .A1(n107145), .A2(n107144), .ZN(n94064) );
  AOI21_X1 U79632 ( .B1(n69424), .B2(n94066), .A(n94068), .ZN(n90302) );
  NOR4_X1 U79633 ( .A1(n94077), .A2(n94078), .A3(n107119), .A4(n94079), .ZN(
        n94066) );
  NAND3_X2 U79634 ( .A1(n104493), .A2(n94080), .A3(n94082), .ZN(n94079) );
  AOI22_X1 U79635 ( .A1(n90119), .A2(n107145), .B1(n90120), .B2(n107144), .ZN(
        n94083) );
  OAI21_X1 U79636 ( .B1(n111056), .B2(n94067), .A(n94068), .ZN(n90298) );
  NAND2_X1 U79637 ( .A1(n94084), .A2(n94085), .ZN(n94067) );
  NOR4_X1 U79638 ( .A1(n94086), .A2(n94087), .A3(n94078), .A4(n94077), .ZN(
        n94085) );
  NOR2_X1 U79639 ( .A1(n90120), .A2(n107144), .ZN(n94077) );
  NOR2_X1 U79640 ( .A1(n90119), .A2(n107145), .ZN(n94078) );
  NOR2_X1 U79641 ( .A1(n59451), .A2(n107122), .ZN(n94087) );
  OAI21_X1 U79642 ( .B1(n59445), .B2(n107114), .A(n94082), .ZN(n94086) );
  XNOR2_X1 U79643 ( .A(n90127), .B(n59452), .ZN(n94082) );
  NOR4_X1 U79644 ( .A1(n94088), .A2(n90136), .A3(n94089), .A4(n94090), .ZN(
        n94084) );
  XNOR2_X1 U79645 ( .A(\DLX_Datapath/RegisterFile/N46177 ), .B(n94091), .ZN(
        n94090) );
  XOR2_X1 U79646 ( .A(n90133), .B(n94092), .Z(n94089) );
  NAND2_X1 U79648 ( .A1(n94094), .A2(n94080), .ZN(n94088) );
  XNOR2_X1 U79649 ( .A(n107128), .B(n59453), .ZN(n94080) );
  XNOR2_X1 U79650 ( .A(\DLX_Datapath/RegisterFile/N46178 ), .B(n94095), .ZN(
        n94094) );
  NOR4_X1 U79651 ( .A1(n94096), .A2(n94097), .A3(n94098), .A4(n94099), .ZN(
        n94059) );
  NAND2_X1 U79652 ( .A1(n94100), .A2(n94101), .ZN(n94099) );
  NOR4_X1 U79653 ( .A1(n94102), .A2(n94103), .A3(n94104), .A4(n94105), .ZN(
        n94101) );
  NAND2_X1 U79654 ( .A1(n94106), .A2(n94107), .ZN(n94105) );
  AOI22_X1 U79655 ( .A1(n90325), .A2(n107213), .B1(n90326), .B2(n107211), .ZN(
        n94107) );
  AND2_X2 U79656 ( .A1(n94108), .A2(n105143), .ZN(n90326) );
  AND2_X2 U79657 ( .A1(n94110), .A2(n105139), .ZN(n90325) );
  AOI22_X1 U79658 ( .A1(n90327), .A2(n107195), .B1(n90328), .B2(n107199), .ZN(
        n94106) );
  AND2_X2 U79659 ( .A1(n94108), .A2(n105141), .ZN(n90328) );
  AND2_X2 U79660 ( .A1(n94113), .A2(n105138), .ZN(n90327) );
  NAND2_X1 U79661 ( .A1(n94115), .A2(n94116), .ZN(n94104) );
  AOI22_X1 U79662 ( .A1(n90331), .A2(n69591), .B1(n90332), .B2(n107205), .ZN(
        n94116) );
  AND2_X2 U79663 ( .A1(n94117), .A2(n94111), .ZN(n90332) );
  AND2_X2 U79664 ( .A1(n94118), .A2(n94119), .ZN(n90331) );
  AOI22_X1 U79665 ( .A1(n90333), .A2(n69484), .B1(n90334), .B2(n107288), .ZN(
        n94115) );
  AND2_X2 U79666 ( .A1(n94118), .A2(n94120), .ZN(n90334) );
  AND2_X2 U79667 ( .A1(n94110), .A2(n94109), .ZN(n90333) );
  NAND2_X1 U79668 ( .A1(n94121), .A2(n94122), .ZN(n94103) );
  AOI22_X1 U79669 ( .A1(n90337), .A2(n107292), .B1(n90338), .B2(n69595), .ZN(
        n94122) );
  AND2_X2 U79670 ( .A1(n94123), .A2(n94119), .ZN(n90338) );
  AND2_X2 U79671 ( .A1(n94124), .A2(n94120), .ZN(n90337) );
  AOI22_X1 U79672 ( .A1(n90339), .A2(n107203), .B1(n90340), .B2(n107209), .ZN(
        n94121) );
  AND2_X2 U79673 ( .A1(n94108), .A2(n105139), .ZN(n90340) );
  AND2_X2 U79674 ( .A1(n94113), .A2(n105143), .ZN(n90339) );
  NAND2_X1 U79675 ( .A1(n94125), .A2(n94126), .ZN(n94102) );
  AOI22_X1 U79676 ( .A1(n90343), .A2(n107290), .B1(n90344), .B2(n107294), .ZN(
        n94126) );
  AND2_X2 U79677 ( .A1(n94118), .A2(n105142), .ZN(n90344) );
  AND2_X2 U79678 ( .A1(n94128), .A2(n94120), .ZN(n90343) );
  AOI22_X1 U79679 ( .A1(n90345), .A2(n107293), .B1(n90346), .B2(n69597), .ZN(
        n94125) );
  AND2_X2 U79680 ( .A1(n94124), .A2(n94119), .ZN(n90346) );
  AND2_X2 U79681 ( .A1(n94118), .A2(n105140), .ZN(n90345) );
  NOR4_X1 U79682 ( .A1(n94130), .A2(n94131), .A3(n94132), .A4(n94133), .ZN(
        n94100) );
  NAND2_X1 U79683 ( .A1(n94134), .A2(n94135), .ZN(n94133) );
  AOI22_X1 U79684 ( .A1(n90353), .A2(n107193), .B1(n90354), .B2(n107187), .ZN(
        n94135) );
  AND2_X2 U79685 ( .A1(n94108), .A2(n94127), .ZN(n90354) );
  AND2_X2 U79686 ( .A1(n94113), .A2(n94112), .ZN(n90353) );
  AOI22_X1 U79687 ( .A1(n90355), .A2(n107185), .B1(n90356), .B2(n107181), .ZN(
        n94134) );
  AND2_X2 U79688 ( .A1(n94117), .A2(n94129), .ZN(n90356) );
  AND2_X2 U79689 ( .A1(n94108), .A2(n105140), .ZN(n90355) );
  NAND2_X1 U79690 ( .A1(n94136), .A2(n94137), .ZN(n94132) );
  AOI22_X1 U79691 ( .A1(n90359), .A2(n107183), .B1(n90360), .B2(n107191), .ZN(
        n94137) );
  AND2_X2 U79692 ( .A1(n94110), .A2(n105142), .ZN(n90360) );
  AND2_X2 U79693 ( .A1(n94117), .A2(n94127), .ZN(n90359) );
  AOI22_X1 U79694 ( .A1(n90361), .A2(n107179), .B1(n90362), .B2(n107189), .ZN(
        n94136) );
  AND2_X2 U79695 ( .A1(n94110), .A2(n94129), .ZN(n90362) );
  AND2_X2 U79696 ( .A1(n94113), .A2(n105142), .ZN(n90361) );
  NAND2_X1 U79697 ( .A1(n94138), .A2(n94139), .ZN(n94131) );
  AOI22_X1 U79698 ( .A1(n90365), .A2(n69464), .B1(n90366), .B2(n69466), .ZN(
        n94139) );
  AND2_X2 U79699 ( .A1(n94110), .A2(n105141), .ZN(n90366) );
  AND2_X2 U79700 ( .A1(n94108), .A2(n94114), .ZN(n90365) );
  NOR2_X1 U79701 ( .A1(n94140), .A2(n94141), .ZN(n94108) );
  AOI22_X1 U79702 ( .A1(n90367), .A2(n69460), .B1(n90368), .B2(n107177), .ZN(
        n94138) );
  AND2_X2 U79703 ( .A1(n94113), .A2(n105140), .ZN(n90368) );
  AND2_X2 U79704 ( .A1(n94117), .A2(n105138), .ZN(n90367) );
  NAND2_X1 U79705 ( .A1(n94142), .A2(n94143), .ZN(n94130) );
  AOI22_X1 U79706 ( .A1(n90371), .A2(n107207), .B1(n90372), .B2(n107197), .ZN(
        n94143) );
  AND2_X2 U79707 ( .A1(n94117), .A2(n94112), .ZN(n90372) );
  AND2_X2 U79708 ( .A1(n94117), .A2(n94109), .ZN(n90371) );
  NOR2_X1 U79709 ( .A1(n94140), .A2(n94144), .ZN(n94117) );
  AOI22_X1 U79710 ( .A1(n90373), .A2(n69470), .B1(n90374), .B2(n107201), .ZN(
        n94142) );
  AND2_X2 U79711 ( .A1(n94110), .A2(n94114), .ZN(n90374) );
  NOR2_X1 U79712 ( .A1(n94140), .A2(n94145), .ZN(n94110) );
  AND2_X2 U79713 ( .A1(n94113), .A2(n94111), .ZN(n90373) );
  NOR2_X1 U79714 ( .A1(n94140), .A2(n94146), .ZN(n94113) );
  OR2_X1 U79715 ( .A1(n94147), .A2(n107095), .ZN(n94140) );
  NAND2_X1 U79716 ( .A1(n94148), .A2(n94149), .ZN(n94098) );
  NOR4_X1 U79717 ( .A1(n94150), .A2(n94151), .A3(n94152), .A4(n94153), .ZN(
        n94149) );
  NAND2_X1 U79718 ( .A1(n94154), .A2(n94155), .ZN(n94153) );
  AOI22_X1 U79719 ( .A1(n90383), .A2(n107303), .B1(n90384), .B2(n107305), .ZN(
        n94155) );
  AND2_X2 U79720 ( .A1(n94124), .A2(n105141), .ZN(n90384) );
  AND2_X2 U79721 ( .A1(n94128), .A2(n105138), .ZN(n90383) );
  AOI22_X1 U79722 ( .A1(n90385), .A2(n69620), .B1(n90386), .B2(n107304), .ZN(
        n94154) );
  AND2_X2 U79723 ( .A1(n94123), .A2(n94112), .ZN(n90386) );
  AND2_X2 U79724 ( .A1(n94123), .A2(n105143), .ZN(n90385) );
  NAND2_X1 U79725 ( .A1(n94156), .A2(n94157), .ZN(n94152) );
  AOI22_X1 U79726 ( .A1(n90389), .A2(n69624), .B1(n90390), .B2(n69626), .ZN(
        n94157) );
  AND2_X2 U79727 ( .A1(n94158), .A2(n94120), .ZN(n90390) );
  AND2_X2 U79728 ( .A1(n94159), .A2(n94120), .ZN(n90389) );
  AOI22_X1 U79729 ( .A1(n90391), .A2(n107311), .B1(n90392), .B2(n107312), .ZN(
        n94156) );
  AND2_X2 U79730 ( .A1(n94159), .A2(n94119), .ZN(n90392) );
  AND2_X2 U79731 ( .A1(n94124), .A2(n94109), .ZN(n90391) );
  NAND2_X1 U79732 ( .A1(n94160), .A2(n94161), .ZN(n94151) );
  AOI22_X1 U79733 ( .A1(n90395), .A2(n107308), .B1(n90396), .B2(n107310), .ZN(
        n94161) );
  AND2_X2 U79734 ( .A1(n94124), .A2(n105139), .ZN(n90396) );
  AND2_X2 U79735 ( .A1(n94128), .A2(n105143), .ZN(n90395) );
  AOI22_X1 U79736 ( .A1(n90397), .A2(n107313), .B1(n90398), .B2(n107309), .ZN(
        n94160) );
  AND2_X2 U79737 ( .A1(n94123), .A2(n94111), .ZN(n90398) );
  AND2_X2 U79738 ( .A1(n94158), .A2(n94119), .ZN(n90397) );
  NAND2_X1 U79739 ( .A1(n94162), .A2(n94163), .ZN(n94150) );
  AOI22_X1 U79740 ( .A1(n90401), .A2(n107318), .B1(n90402), .B2(n69631), .ZN(
        n94163) );
  AND2_X2 U79741 ( .A1(n94159), .A2(n94129), .ZN(n90402) );
  AND2_X2 U79742 ( .A1(n94158), .A2(n105140), .ZN(n90401) );
  AOI22_X1 U79743 ( .A1(n90403), .A2(n107317), .B1(n90404), .B2(n69629), .ZN(
        n94162) );
  AND2_X2 U79744 ( .A1(n94164), .A2(n94119), .ZN(n90404) );
  AND2_X2 U79745 ( .A1(n94159), .A2(n94127), .ZN(n90403) );
  NOR4_X1 U79746 ( .A1(n94165), .A2(n94166), .A3(n94167), .A4(n94168), .ZN(
        n94148) );
  NAND2_X1 U79747 ( .A1(n94169), .A2(n94170), .ZN(n94168) );
  AOI22_X1 U79748 ( .A1(n90411), .A2(n107298), .B1(n90412), .B2(n107289), .ZN(
        n94170) );
  AND2_X2 U79749 ( .A1(n94128), .A2(n94119), .ZN(n90412) );
  AND2_X2 U79750 ( .A1(n94124), .A2(n94129), .ZN(n90411) );
  AOI22_X1 U79751 ( .A1(n90413), .A2(n107291), .B1(n90414), .B2(n69603), .ZN(
        n94169) );
  AND2_X2 U79752 ( .A1(n94123), .A2(n105140), .ZN(n90414) );
  AND2_X2 U79753 ( .A1(n94123), .A2(n94120), .ZN(n90413) );
  NAND2_X1 U79754 ( .A1(n94171), .A2(n94172), .ZN(n94167) );
  AOI22_X1 U79755 ( .A1(n90417), .A2(n107296), .B1(n90418), .B2(n107300), .ZN(
        n94172) );
  AND2_X2 U79756 ( .A1(n94118), .A2(n105141), .ZN(n90418) );
  AND2_X2 U79757 ( .A1(n94128), .A2(n105142), .ZN(n90417) );
  AOI22_X1 U79758 ( .A1(n90419), .A2(n107302), .B1(n90420), .B2(n107299), .ZN(
        n94171) );
  AND2_X2 U79759 ( .A1(n94124), .A2(n94127), .ZN(n90420) );
  AND2_X2 U79760 ( .A1(n94128), .A2(n94112), .ZN(n90419) );
  NAND2_X1 U79761 ( .A1(n94173), .A2(n94174), .ZN(n94166) );
  AOI22_X1 U79762 ( .A1(n90423), .A2(n69612), .B1(n90424), .B2(n107295), .ZN(
        n94174) );
  AND2_X2 U79763 ( .A1(n94128), .A2(n94129), .ZN(n90424) );
  AND2_X2 U79764 ( .A1(n94123), .A2(n94114), .ZN(n90423) );
  AOI22_X1 U79765 ( .A1(n90425), .A2(n107297), .B1(n90426), .B2(n107301), .ZN(
        n94173) );
  AND2_X2 U79766 ( .A1(n94118), .A2(n105138), .ZN(n90426) );
  AND2_X2 U79767 ( .A1(n94123), .A2(n105142), .ZN(n90425) );
  NOR2_X1 U79768 ( .A1(n94175), .A2(n94147), .ZN(n94123) );
  OR2_X1 U79769 ( .A1(n94141), .A2(n94176), .ZN(n94175) );
  NAND2_X1 U79770 ( .A1(n94177), .A2(n94178), .ZN(n94165) );
  AOI22_X1 U79771 ( .A1(n90429), .A2(n107307), .B1(n90430), .B2(n69616), .ZN(
        n94178) );
  AND2_X2 U79772 ( .A1(n94118), .A2(n94109), .ZN(n90430) );
  AND2_X2 U79773 ( .A1(n94128), .A2(n105139), .ZN(n90429) );
  NOR2_X1 U79774 ( .A1(n94179), .A2(n94147), .ZN(n94128) );
  OR2_X1 U79775 ( .A1(n94144), .A2(n94176), .ZN(n94179) );
  AOI22_X1 U79776 ( .A1(n90431), .A2(n69614), .B1(n90432), .B2(n107306), .ZN(
        n94177) );
  AND2_X2 U79777 ( .A1(n94118), .A2(n94111), .ZN(n90432) );
  NOR2_X1 U79778 ( .A1(n94180), .A2(n94147), .ZN(n94118) );
  OR2_X1 U79779 ( .A1(n94146), .A2(n94176), .ZN(n94180) );
  AND2_X2 U79780 ( .A1(n94124), .A2(n94114), .ZN(n90431) );
  NOR2_X1 U79781 ( .A1(n94181), .A2(n94147), .ZN(n94124) );
  OR2_X1 U79782 ( .A1(n94145), .A2(n94176), .ZN(n94181) );
  NAND2_X1 U79783 ( .A1(n94182), .A2(n94183), .ZN(n94097) );
  NOR4_X1 U79784 ( .A1(n94184), .A2(n94185), .A3(n94186), .A4(n94187), .ZN(
        n94183) );
  NAND2_X1 U79785 ( .A1(n94188), .A2(n94189), .ZN(n94187) );
  AOI22_X1 U79786 ( .A1(n90441), .A2(n69654), .B1(n90442), .B2(n107328), .ZN(
        n94189) );
  AND2_X2 U79787 ( .A1(n94164), .A2(n105141), .ZN(n90442) );
  AND2_X2 U79788 ( .A1(n94164), .A2(n105143), .ZN(n90441) );
  AOI22_X1 U79789 ( .A1(n90443), .A2(n107332), .B1(n90444), .B2(n107331), .ZN(
        n94188) );
  AND2_X2 U79790 ( .A1(n94158), .A2(n94109), .ZN(n90444) );
  AND2_X2 U79791 ( .A1(n94190), .A2(n105139), .ZN(n90443) );
  NAND2_X1 U79792 ( .A1(n94191), .A2(n94192), .ZN(n94186) );
  AOI22_X1 U79793 ( .A1(n90447), .A2(n107337), .B1(n90448), .B2(n107336), .ZN(
        n94192) );
  AND2_X2 U79794 ( .A1(n94120), .A2(n94193), .ZN(n90448) );
  AND2_X2 U79795 ( .A1(n94119), .A2(n94194), .ZN(n90447) );
  AOI22_X1 U79796 ( .A1(n90449), .A2(n107327), .B1(n90450), .B2(n107329), .ZN(
        n94191) );
  AND2_X2 U79797 ( .A1(n94159), .A2(n94111), .ZN(n90450) );
  AND2_X2 U79798 ( .A1(n94190), .A2(n105138), .ZN(n90449) );
  NAND2_X1 U79799 ( .A1(n94195), .A2(n94196), .ZN(n94185) );
  AOI22_X1 U79800 ( .A1(n90453), .A2(n107338), .B1(n90454), .B2(n107334), .ZN(
        n94196) );
  AND2_X2 U79801 ( .A1(n94164), .A2(n105139), .ZN(n90454) );
  AND2_X2 U79802 ( .A1(n94119), .A2(n94197), .ZN(n90453) );
  AOI22_X1 U79803 ( .A1(n90455), .A2(n69658), .B1(n90456), .B2(n69660), .ZN(
        n94195) );
  AND2_X2 U79804 ( .A1(n94120), .A2(n94197), .ZN(n90456) );
  AND2_X2 U79805 ( .A1(n94120), .A2(n94194), .ZN(n90455) );
  NAND2_X1 U79806 ( .A1(n94198), .A2(n94199), .ZN(n94184) );
  AOI22_X1 U79807 ( .A1(n90459), .A2(n107341), .B1(n90460), .B2(n69666), .ZN(
        n94199) );
  AND2_X2 U79808 ( .A1(n105142), .A2(n94194), .ZN(n90460) );
  AND2_X2 U79809 ( .A1(n105140), .A2(n94193), .ZN(n90459) );
  AOI22_X1 U79810 ( .A1(n90461), .A2(n107333), .B1(n90462), .B2(n107335), .ZN(
        n94198) );
  AND2_X2 U79811 ( .A1(n94119), .A2(n94193), .ZN(n90462) );
  AND2_X2 U79812 ( .A1(n94190), .A2(n105143), .ZN(n90461) );
  NOR4_X1 U79813 ( .A1(n94200), .A2(n94201), .A3(n94202), .A4(n94203), .ZN(
        n94182) );
  NAND2_X1 U79814 ( .A1(n94204), .A2(n94205), .ZN(n94203) );
  AOI22_X1 U79815 ( .A1(n90469), .A2(n107316), .B1(n90470), .B2(n107321), .ZN(
        n94205) );
  AND2_X2 U79816 ( .A1(n94164), .A2(n105140), .ZN(n90470) );
  AND2_X2 U79817 ( .A1(n94164), .A2(n94120), .ZN(n90469) );
  AOI22_X1 U79818 ( .A1(n90471), .A2(n107315), .B1(n90472), .B2(n69634), .ZN(
        n94204) );
  AND2_X2 U79819 ( .A1(n94158), .A2(n94127), .ZN(n90472) );
  AND2_X2 U79820 ( .A1(n94190), .A2(n94120), .ZN(n90471) );
  NAND2_X1 U79821 ( .A1(n94206), .A2(n94207), .ZN(n94202) );
  AOI22_X1 U79822 ( .A1(n90475), .A2(n69643), .B1(n90476), .B2(n107323), .ZN(
        n94207) );
  AND2_X2 U79823 ( .A1(n94159), .A2(n94112), .ZN(n90476) );
  AND2_X2 U79824 ( .A1(n94190), .A2(n105141), .ZN(n90475) );
  AOI22_X1 U79825 ( .A1(n90477), .A2(n107324), .B1(n90478), .B2(n107314), .ZN(
        n94206) );
  AND2_X2 U79826 ( .A1(n94190), .A2(n94119), .ZN(n90478) );
  AND2_X2 U79827 ( .A1(n94159), .A2(n94114), .ZN(n90477) );
  NAND2_X1 U79828 ( .A1(n94208), .A2(n94209), .ZN(n94201) );
  AOI22_X1 U79829 ( .A1(n90481), .A2(n107322), .B1(n90482), .B2(n107326), .ZN(
        n94209) );
  AND2_X2 U79830 ( .A1(n94158), .A2(n105138), .ZN(n90482) );
  AND2_X2 U79831 ( .A1(n94164), .A2(n105142), .ZN(n90481) );
  AOI22_X1 U79832 ( .A1(n90483), .A2(n107320), .B1(n90484), .B2(n107325), .ZN(
        n94208) );
  AND2_X2 U79833 ( .A1(n94158), .A2(n94112), .ZN(n90484) );
  AND2_X2 U79834 ( .A1(n94190), .A2(n94127), .ZN(n90483) );
  NAND2_X1 U79835 ( .A1(n94210), .A2(n94211), .ZN(n94200) );
  AOI22_X1 U79836 ( .A1(n90487), .A2(n69648), .B1(n90488), .B2(n107330), .ZN(
        n94211) );
  AND2_X2 U79837 ( .A1(n94158), .A2(n94111), .ZN(n90488) );
  NOR2_X1 U79838 ( .A1(n94212), .A2(n94144), .ZN(n94158) );
  AND2_X2 U79839 ( .A1(n94159), .A2(n94109), .ZN(n90487) );
  NOR2_X1 U79840 ( .A1(n94212), .A2(n94146), .ZN(n94159) );
  AOI22_X1 U79841 ( .A1(n90489), .A2(n69646), .B1(n90490), .B2(n107319), .ZN(
        n94210) );
  AND2_X2 U79842 ( .A1(n94190), .A2(n94129), .ZN(n90490) );
  NOR2_X1 U79843 ( .A1(n94212), .A2(n94141), .ZN(n94190) );
  AND2_X2 U79844 ( .A1(n94164), .A2(n94114), .ZN(n90489) );
  NOR2_X1 U79845 ( .A1(n94212), .A2(n94145), .ZN(n94164) );
  NAND2_X1 U79846 ( .A1(n94176), .A2(n94147), .ZN(n94212) );
  NAND2_X1 U79847 ( .A1(n94213), .A2(n94214), .ZN(n94096) );
  NOR4_X1 U79848 ( .A1(n94215), .A2(n94216), .A3(n94217), .A4(n94218), .ZN(
        n94214) );
  NAND2_X1 U79849 ( .A1(n94219), .A2(n94220), .ZN(n94218) );
  AOI22_X1 U79850 ( .A1(n90499), .A2(n107359), .B1(n90500), .B2(n107358), .ZN(
        n94220) );
  AND2_X2 U79851 ( .A1(n94197), .A2(n105143), .ZN(n90500) );
  AND2_X2 U79852 ( .A1(n94111), .A2(n94221), .ZN(n90499) );
  AOI22_X1 U79853 ( .A1(n90501), .A2(n69682), .B1(n90502), .B2(n107356), .ZN(
        n94219) );
  AND2_X2 U79854 ( .A1(n94193), .A2(n94109), .ZN(n90502) );
  AND2_X2 U79855 ( .A1(n94194), .A2(n105143), .ZN(n90501) );
  NAND2_X1 U79856 ( .A1(n94222), .A2(n94223), .ZN(n94217) );
  AOI22_X1 U79857 ( .A1(n90505), .A2(n107354), .B1(n90506), .B2(n107357), .ZN(
        n94223) );
  AND2_X2 U79858 ( .A1(n94194), .A2(n105139), .ZN(n90506) );
  AND2_X2 U79859 ( .A1(n94114), .A2(n94221), .ZN(n90505) );
  AOI22_X1 U79860 ( .A1(n105651), .A2(n69688), .B1(n90508), .B2(n107355), .ZN(
        n94222) );
  AND2_X2 U79861 ( .A1(n94193), .A2(n94111), .ZN(n90508) );
  NOR2_X1 U79862 ( .A1(n94224), .A2(n94146), .ZN(n90507) );
  NAND2_X1 U79863 ( .A1(n94225), .A2(n94226), .ZN(n94216) );
  AOI22_X1 U79864 ( .A1(n105650), .A2(n107364), .B1(n105649), .B2(n69694), 
        .ZN(n94226) );
  NOR2_X1 U79865 ( .A1(n94224), .A2(n94145), .ZN(n90512) );
  NOR2_X1 U79866 ( .A1(n94141), .A2(n94224), .ZN(n90511) );
  AOI22_X1 U79867 ( .A1(n105648), .A2(n107362), .B1(n105647), .B2(n107363), 
        .ZN(n94225) );
  NOR2_X1 U79868 ( .A1(n94141), .A2(n94227), .ZN(n90514) );
  NOR2_X1 U79869 ( .A1(n94224), .A2(n94144), .ZN(n90513) );
  OR2_X1 U79870 ( .A1(n94228), .A2(n59445), .ZN(n94224) );
  NAND2_X1 U79871 ( .A1(n94229), .A2(n94230), .ZN(n94215) );
  AOI22_X1 U79872 ( .A1(n90517), .A2(n107360), .B1(n105646), .B2(n69689), .ZN(
        n94230) );
  NOR2_X1 U79873 ( .A1(n94144), .A2(n94227), .ZN(n90518) );
  AND2_X2 U79874 ( .A1(n94109), .A2(n94221), .ZN(n90517) );
  NOR2_X1 U79875 ( .A1(n94231), .A2(n107098), .ZN(n94109) );
  AOI22_X1 U79876 ( .A1(n105645), .A2(n107365), .B1(n105644), .B2(n107361), 
        .ZN(n94229) );
  NOR2_X1 U79877 ( .A1(n94146), .A2(n94227), .ZN(n90520) );
  NOR2_X1 U79878 ( .A1(n94227), .A2(n94145), .ZN(n90519) );
  OR2_X1 U79879 ( .A1(n94228), .A2(n107144), .ZN(n94227) );
  NAND2_X1 U79880 ( .A1(n94232), .A2(n94095), .ZN(n94228) );
  NOR4_X1 U79881 ( .A1(n94233), .A2(n94234), .A3(n94235), .A4(n94236), .ZN(
        n94213) );
  NAND2_X1 U79882 ( .A1(n94237), .A2(n94238), .ZN(n94236) );
  AOI22_X1 U79883 ( .A1(n90527), .A2(n107340), .B1(n90528), .B2(n107344), .ZN(
        n94238) );
  AND2_X2 U79884 ( .A1(n94127), .A2(n94197), .ZN(n90528) );
  AND2_X2 U79885 ( .A1(n94120), .A2(n94221), .ZN(n90527) );
  NOR2_X1 U79886 ( .A1(n94239), .A2(n104707), .ZN(n94120) );
  NAND2_X1 U79887 ( .A1(n107144), .A2(n107098), .ZN(n94239) );
  AOI22_X1 U79888 ( .A1(n90529), .A2(n107343), .B1(n90530), .B2(n69665), .ZN(
        n94237) );
  AND2_X2 U79889 ( .A1(n94129), .A2(n94194), .ZN(n90530) );
  AND2_X2 U79890 ( .A1(n105140), .A2(n94197), .ZN(n90529) );
  NAND2_X1 U79891 ( .A1(n94240), .A2(n94241), .ZN(n94235) );
  AOI22_X1 U79892 ( .A1(n90533), .A2(n107350), .B1(n90534), .B2(n107339), .ZN(
        n94241) );
  AND2_X2 U79893 ( .A1(n94119), .A2(n94221), .ZN(n90534) );
  NOR2_X1 U79894 ( .A1(n94242), .A2(n107144), .ZN(n94119) );
  NAND2_X1 U79895 ( .A1(n107098), .A2(n59453), .ZN(n94242) );
  AND2_X2 U79896 ( .A1(n94194), .A2(n105138), .ZN(n90533) );
  AOI22_X1 U79897 ( .A1(n90535), .A2(n107342), .B1(n90536), .B2(n107347), .ZN(
        n94240) );
  AND2_X2 U79898 ( .A1(n105141), .A2(n94193), .ZN(n90536) );
  AND2_X2 U79899 ( .A1(n105142), .A2(n94193), .ZN(n90535) );
  NAND2_X1 U79900 ( .A1(n94243), .A2(n94244), .ZN(n94234) );
  AOI22_X1 U79901 ( .A1(n90539), .A2(n107346), .B1(n90540), .B2(n107351), .ZN(
        n94244) );
  AND2_X2 U79902 ( .A1(n94112), .A2(n94197), .ZN(n90540) );
  AND2_X2 U79903 ( .A1(n94127), .A2(n94221), .ZN(n90539) );
  NOR2_X1 U79904 ( .A1(n94231), .A2(n94245), .ZN(n94127) );
  NAND2_X1 U79905 ( .A1(n104707), .A2(n107144), .ZN(n94231) );
  AOI22_X1 U79906 ( .A1(n90541), .A2(n107353), .B1(n90542), .B2(n107349), .ZN(
        n94243) );
  AND2_X2 U79907 ( .A1(n105141), .A2(n94194), .ZN(n90542) );
  NOR2_X1 U79908 ( .A1(n94144), .A2(n94246), .ZN(n94194) );
  NAND2_X1 U79909 ( .A1(n59452), .A2(n107145), .ZN(n94144) );
  AND2_X2 U79910 ( .A1(n94112), .A2(n94221), .ZN(n90541) );
  NOR2_X1 U79911 ( .A1(n94247), .A2(n107098), .ZN(n94112) );
  NAND2_X1 U79912 ( .A1(n59453), .A2(n59445), .ZN(n94247) );
  NAND2_X1 U79913 ( .A1(n94248), .A2(n94249), .ZN(n94233) );
  AOI22_X1 U79914 ( .A1(n90545), .A2(n69683), .B1(n90546), .B2(n107345), .ZN(
        n94249) );
  AND2_X2 U79915 ( .A1(n94129), .A2(n94221), .ZN(n90546) );
  NOR2_X1 U79916 ( .A1(n94145), .A2(n94246), .ZN(n94221) );
  NAND2_X1 U79917 ( .A1(n105061), .A2(n107145), .ZN(n94145) );
  NOR2_X1 U79918 ( .A1(n94250), .A2(n107144), .ZN(n94129) );
  NAND2_X1 U79919 ( .A1(n104707), .A2(n107098), .ZN(n94250) );
  AND2_X2 U79920 ( .A1(n94197), .A2(n105139), .ZN(n90545) );
  NOR2_X1 U79921 ( .A1(n94251), .A2(n107098), .ZN(n94111) );
  NAND2_X1 U79922 ( .A1(n104707), .A2(n59445), .ZN(n94251) );
  AOI22_X1 U79923 ( .A1(n90547), .A2(n107348), .B1(n90548), .B2(n107352), .ZN(
        n94248) );
  AND2_X2 U79924 ( .A1(n94197), .A2(n94114), .ZN(n90548) );
  NOR2_X1 U79925 ( .A1(n94141), .A2(n94246), .ZN(n94197) );
  NAND2_X1 U79926 ( .A1(n59451), .A2(n105061), .ZN(n94141) );
  AND2_X2 U79927 ( .A1(n94193), .A2(n105138), .ZN(n90547) );
  NOR2_X1 U79928 ( .A1(n94252), .A2(n107098), .ZN(n94114) );
  XOR2_X1 U79929 ( .A(n104707), .B(n94092), .Z(n94245) );
  AOI21_X1 U79930 ( .B1(n104707), .B2(n94253), .A(n94254), .ZN(n94092) );
  NAND2_X1 U79931 ( .A1(n107144), .A2(n59453), .ZN(n94252) );
  NOR2_X1 U79932 ( .A1(n94146), .A2(n94246), .ZN(n94193) );
  NAND2_X1 U79933 ( .A1(n107095), .A2(n94147), .ZN(n94246) );
  XOR2_X1 U79934 ( .A(n94095), .B(n94232), .Z(n94147) );
  NOR2_X1 U79935 ( .A1(n94091), .A2(n107097), .ZN(n94232) );
  XNOR2_X1 U79936 ( .A(n104994), .B(n94256), .ZN(n94095) );
  NOR2_X1 U79937 ( .A1(n104997), .A2(n107097), .ZN(n94256) );
  XOR2_X1 U79938 ( .A(n94091), .B(n94254), .Z(n94176) );
  XNOR2_X1 U79939 ( .A(n104997), .B(n94254), .ZN(n94091) );
  NOR2_X1 U79940 ( .A1(n94253), .A2(n104707), .ZN(n94254) );
  NAND2_X1 U79941 ( .A1(n59451), .A2(n59452), .ZN(n94146) );
  XOR2_X1 U79943 ( .A(n106764), .B(
        \dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .Z(
        \DLX_Datapath/RegisterFile/N27074 ) );
  OAI21_X1 U79975 ( .B1(n103351), .B2(n94260), .A(n94261), .ZN(
        \DLX_Datapath/RegisterFile/N26858 ) );
  NAND2_X1 U79976 ( .A1(n107117), .A2(n86303), .ZN(n94261) );
  OAI21_X1 U79977 ( .B1(n103338), .B2(n94260), .A(n94262), .ZN(
        \DLX_Datapath/RegisterFile/N26857 ) );
  NAND2_X1 U79978 ( .A1(n107117), .A2(n86558), .ZN(n94262) );
  OAI21_X1 U79979 ( .B1(n103327), .B2(n94260), .A(n94263), .ZN(
        \DLX_Datapath/RegisterFile/N26856 ) );
  NAND2_X1 U79980 ( .A1(n107117), .A2(n86676), .ZN(n94263) );
  OAI21_X1 U79981 ( .B1(n103311), .B2(n94260), .A(n94264), .ZN(
        \DLX_Datapath/RegisterFile/N26855 ) );
  NAND2_X1 U79982 ( .A1(n107117), .A2(n86794), .ZN(n94264) );
  OAI21_X1 U79983 ( .B1(n103294), .B2(n94260), .A(n94265), .ZN(
        \DLX_Datapath/RegisterFile/N26854 ) );
  NAND2_X1 U79984 ( .A1(n107117), .A2(n86912), .ZN(n94265) );
  OAI21_X1 U79985 ( .B1(n103275), .B2(n94260), .A(n94266), .ZN(
        \DLX_Datapath/RegisterFile/N26853 ) );
  NAND2_X1 U79986 ( .A1(n107117), .A2(n87030), .ZN(n94266) );
  OAI21_X1 U79987 ( .B1(n103256), .B2(n94260), .A(n94267), .ZN(
        \DLX_Datapath/RegisterFile/N26852 ) );
  NAND2_X1 U79988 ( .A1(n107117), .A2(n87148), .ZN(n94267) );
  OAI21_X1 U79989 ( .B1(n103237), .B2(n94260), .A(n94268), .ZN(
        \DLX_Datapath/RegisterFile/N26851 ) );
  NAND2_X1 U79990 ( .A1(n107117), .A2(n87266), .ZN(n94268) );
  OAI21_X1 U79991 ( .B1(n103218), .B2(n105643), .A(n94269), .ZN(
        \DLX_Datapath/RegisterFile/N26850 ) );
  NAND2_X1 U79992 ( .A1(n105214), .A2(n87384), .ZN(n94269) );
  OAI21_X1 U79993 ( .B1(n103200), .B2(n105643), .A(n94270), .ZN(
        \DLX_Datapath/RegisterFile/N26849 ) );
  NAND2_X1 U79994 ( .A1(n105214), .A2(n87502), .ZN(n94270) );
  OAI21_X1 U79995 ( .B1(n103181), .B2(n105643), .A(n94271), .ZN(
        \DLX_Datapath/RegisterFile/N26848 ) );
  NAND2_X1 U79996 ( .A1(n105214), .A2(n87620), .ZN(n94271) );
  OAI21_X1 U79997 ( .B1(n103162), .B2(n105643), .A(n94272), .ZN(
        \DLX_Datapath/RegisterFile/N26847 ) );
  NAND2_X1 U79998 ( .A1(n105214), .A2(n87738), .ZN(n94272) );
  OAI21_X1 U79999 ( .B1(n103142), .B2(n105643), .A(n94273), .ZN(
        \DLX_Datapath/RegisterFile/N26846 ) );
  NAND2_X1 U80000 ( .A1(n105214), .A2(n87856), .ZN(n94273) );
  OAI21_X1 U80001 ( .B1(n103124), .B2(n105643), .A(n94274), .ZN(
        \DLX_Datapath/RegisterFile/N26845 ) );
  NAND2_X1 U80002 ( .A1(n105214), .A2(n87974), .ZN(n94274) );
  OAI21_X1 U80003 ( .B1(n103104), .B2(n105643), .A(n94275), .ZN(
        \DLX_Datapath/RegisterFile/N26844 ) );
  NAND2_X1 U80004 ( .A1(n105214), .A2(n88092), .ZN(n94275) );
  OAI21_X1 U80005 ( .B1(n103084), .B2(n105643), .A(n94276), .ZN(
        \DLX_Datapath/RegisterFile/N26843 ) );
  NAND2_X1 U80006 ( .A1(n105214), .A2(n88210), .ZN(n94276) );
  OAI21_X1 U80007 ( .B1(n103064), .B2(n105643), .A(n94277), .ZN(
        \DLX_Datapath/RegisterFile/N26842 ) );
  NAND2_X1 U80008 ( .A1(n105214), .A2(n88328), .ZN(n94277) );
  OAI21_X1 U80009 ( .B1(n103044), .B2(n105643), .A(n94278), .ZN(
        \DLX_Datapath/RegisterFile/N26841 ) );
  NAND2_X1 U80010 ( .A1(n105214), .A2(n88446), .ZN(n94278) );
  OAI21_X1 U80011 ( .B1(n103024), .B2(n105643), .A(n94279), .ZN(
        \DLX_Datapath/RegisterFile/N26840 ) );
  NAND2_X1 U80012 ( .A1(n105214), .A2(n88564), .ZN(n94279) );
  OAI21_X1 U80013 ( .B1(n103004), .B2(n105643), .A(n94280), .ZN(
        \DLX_Datapath/RegisterFile/N26839 ) );
  NAND2_X1 U80014 ( .A1(n105214), .A2(n88682), .ZN(n94280) );
  OAI21_X1 U80015 ( .B1(n102984), .B2(n105642), .A(n94281), .ZN(
        \DLX_Datapath/RegisterFile/N26838 ) );
  NAND2_X1 U80016 ( .A1(n105213), .A2(n88800), .ZN(n94281) );
  OAI21_X1 U80017 ( .B1(n102967), .B2(n105642), .A(n94282), .ZN(
        \DLX_Datapath/RegisterFile/N26837 ) );
  NAND2_X1 U80018 ( .A1(n105213), .A2(n88918), .ZN(n94282) );
  OAI21_X1 U80019 ( .B1(n102947), .B2(n105642), .A(n94283), .ZN(
        \DLX_Datapath/RegisterFile/N26836 ) );
  NAND2_X1 U80020 ( .A1(n105213), .A2(n81794), .ZN(n94283) );
  OAI21_X1 U80021 ( .B1(n102927), .B2(n105642), .A(n94284), .ZN(
        \DLX_Datapath/RegisterFile/N26835 ) );
  NAND2_X1 U80022 ( .A1(n105213), .A2(n89153), .ZN(n94284) );
  OAI21_X1 U80023 ( .B1(n102907), .B2(n105642), .A(n94285), .ZN(
        \DLX_Datapath/RegisterFile/N26834 ) );
  NAND2_X1 U80024 ( .A1(n105213), .A2(n89271), .ZN(n94285) );
  OAI21_X1 U80025 ( .B1(n102887), .B2(n105642), .A(n94286), .ZN(
        \DLX_Datapath/RegisterFile/N26833 ) );
  NAND2_X1 U80026 ( .A1(n105213), .A2(n81792), .ZN(n94286) );
  OAI21_X1 U80027 ( .B1(n102867), .B2(n105642), .A(n94287), .ZN(
        \DLX_Datapath/RegisterFile/N26832 ) );
  NAND2_X1 U80028 ( .A1(n105213), .A2(n89506), .ZN(n94287) );
  OAI21_X1 U80029 ( .B1(n102847), .B2(n105642), .A(n94288), .ZN(
        \DLX_Datapath/RegisterFile/N26831 ) );
  NAND2_X1 U80030 ( .A1(n105213), .A2(n89624), .ZN(n94288) );
  OAI21_X1 U80031 ( .B1(n102827), .B2(n105642), .A(n94289), .ZN(
        \DLX_Datapath/RegisterFile/N26830 ) );
  NAND2_X1 U80032 ( .A1(n105213), .A2(n89742), .ZN(n94289) );
  OAI21_X1 U80033 ( .B1(n102807), .B2(n105642), .A(n94290), .ZN(
        \DLX_Datapath/RegisterFile/N26829 ) );
  NAND2_X1 U80034 ( .A1(n105213), .A2(n81790), .ZN(n94290) );
  OAI21_X1 U80035 ( .B1(n102787), .B2(n105642), .A(n94291), .ZN(
        \DLX_Datapath/RegisterFile/N26828 ) );
  NAND2_X1 U80036 ( .A1(n105213), .A2(n89977), .ZN(n94291) );
  OAI21_X1 U80037 ( .B1(n102767), .B2(n105642), .A(n94292), .ZN(
        \DLX_Datapath/RegisterFile/N26827 ) );
  NAND2_X1 U80038 ( .A1(n105213), .A2(n90096), .ZN(n94292) );
  NAND2_X1 U80039 ( .A1(n94294), .A2(n94293), .ZN(n94260) );
  NAND2_X1 U80040 ( .A1(n105137), .A2(n94296), .ZN(n94293) );
  OAI21_X1 U80041 ( .B1(n107945), .B2(n105641), .A(n94298), .ZN(
        \DLX_Datapath/RegisterFile/N26826 ) );
  NAND2_X1 U80042 ( .A1(n107116), .A2(n86303), .ZN(n94298) );
  OAI21_X1 U80043 ( .B1(n108041), .B2(n105641), .A(n94299), .ZN(
        \DLX_Datapath/RegisterFile/N26825 ) );
  NAND2_X1 U80044 ( .A1(n107116), .A2(n86558), .ZN(n94299) );
  OAI21_X1 U80045 ( .B1(n107166), .B2(n105641), .A(n94300), .ZN(
        \DLX_Datapath/RegisterFile/N26824 ) );
  NAND2_X1 U80046 ( .A1(n107116), .A2(n86676), .ZN(n94300) );
  OAI21_X1 U80047 ( .B1(n107850), .B2(n105641), .A(n94301), .ZN(
        \DLX_Datapath/RegisterFile/N26823 ) );
  NAND2_X1 U80048 ( .A1(n107116), .A2(n86794), .ZN(n94301) );
  OAI21_X1 U80049 ( .B1(n110745), .B2(n105641), .A(n94302), .ZN(
        \DLX_Datapath/RegisterFile/N26822 ) );
  NAND2_X1 U80050 ( .A1(n107116), .A2(n86912), .ZN(n94302) );
  OAI21_X1 U80051 ( .B1(n108150), .B2(n105641), .A(n94303), .ZN(
        \DLX_Datapath/RegisterFile/N26821 ) );
  NAND2_X1 U80052 ( .A1(n107116), .A2(n87030), .ZN(n94303) );
  OAI21_X1 U80053 ( .B1(n110848), .B2(n105641), .A(n94304), .ZN(
        \DLX_Datapath/RegisterFile/N26820 ) );
  NAND2_X1 U80054 ( .A1(n107116), .A2(n87148), .ZN(n94304) );
  OAI21_X1 U80055 ( .B1(n110949), .B2(n105641), .A(n94305), .ZN(
        \DLX_Datapath/RegisterFile/N26819 ) );
  NAND2_X1 U80056 ( .A1(n107116), .A2(n87266), .ZN(n94305) );
  OAI21_X1 U80057 ( .B1(n110542), .B2(n105640), .A(n94306), .ZN(
        \DLX_Datapath/RegisterFile/N26818 ) );
  NAND2_X1 U80058 ( .A1(n105212), .A2(n87384), .ZN(n94306) );
  OAI21_X1 U80059 ( .B1(n110327), .B2(n105640), .A(n94307), .ZN(
        \DLX_Datapath/RegisterFile/N26817 ) );
  NAND2_X1 U80060 ( .A1(n105212), .A2(n87502), .ZN(n94307) );
  OAI21_X1 U80061 ( .B1(n110647), .B2(n105640), .A(n94308), .ZN(
        \DLX_Datapath/RegisterFile/N26816 ) );
  NAND2_X1 U80062 ( .A1(n105212), .A2(n87620), .ZN(n94308) );
  OAI21_X1 U80063 ( .B1(n110436), .B2(n105640), .A(n94309), .ZN(
        \DLX_Datapath/RegisterFile/N26815 ) );
  NAND2_X1 U80064 ( .A1(n105212), .A2(n87738), .ZN(n94309) );
  OAI21_X1 U80065 ( .B1(n110114), .B2(n105640), .A(n94310), .ZN(
        \DLX_Datapath/RegisterFile/N26814 ) );
  NAND2_X1 U80066 ( .A1(n105212), .A2(n87856), .ZN(n94310) );
  OAI21_X1 U80067 ( .B1(n110221), .B2(n105640), .A(n94311), .ZN(
        \DLX_Datapath/RegisterFile/N26813 ) );
  NAND2_X1 U80068 ( .A1(n105212), .A2(n87974), .ZN(n94311) );
  OAI21_X1 U80069 ( .B1(n110006), .B2(n105640), .A(n94312), .ZN(
        \DLX_Datapath/RegisterFile/N26812 ) );
  NAND2_X1 U80070 ( .A1(n105212), .A2(n88092), .ZN(n94312) );
  OAI21_X1 U80071 ( .B1(n109889), .B2(n105640), .A(n94313), .ZN(
        \DLX_Datapath/RegisterFile/N26811 ) );
  NAND2_X1 U80072 ( .A1(n105212), .A2(n88210), .ZN(n94313) );
  OAI21_X1 U80073 ( .B1(n108263), .B2(n105640), .A(n94314), .ZN(
        \DLX_Datapath/RegisterFile/N26810 ) );
  NAND2_X1 U80074 ( .A1(n105212), .A2(n88328), .ZN(n94314) );
  OAI21_X1 U80075 ( .B1(n108386), .B2(n105640), .A(n94315), .ZN(
        \DLX_Datapath/RegisterFile/N26809 ) );
  NAND2_X1 U80076 ( .A1(n105212), .A2(n88446), .ZN(n94315) );
  OAI21_X1 U80077 ( .B1(n108497), .B2(n105640), .A(n94316), .ZN(
        \DLX_Datapath/RegisterFile/N26808 ) );
  NAND2_X1 U80078 ( .A1(n105212), .A2(n88564), .ZN(n94316) );
  OAI21_X1 U80079 ( .B1(n107734), .B2(n105640), .A(n94317), .ZN(
        \DLX_Datapath/RegisterFile/N26807 ) );
  NAND2_X1 U80080 ( .A1(n105212), .A2(n88682), .ZN(n94317) );
  OAI21_X1 U80081 ( .B1(n109649), .B2(n105641), .A(n94318), .ZN(
        \DLX_Datapath/RegisterFile/N26806 ) );
  NAND2_X1 U80082 ( .A1(n105211), .A2(n88800), .ZN(n94318) );
  OAI21_X1 U80083 ( .B1(n108611), .B2(n105641), .A(n94319), .ZN(
        \DLX_Datapath/RegisterFile/N26805 ) );
  NAND2_X1 U80084 ( .A1(n105211), .A2(n88918), .ZN(n94319) );
  OAI21_X1 U80085 ( .B1(n109756), .B2(n105641), .A(n94320), .ZN(
        \DLX_Datapath/RegisterFile/N26804 ) );
  NAND2_X1 U80086 ( .A1(n105211), .A2(n81794), .ZN(n94320) );
  OAI21_X1 U80087 ( .B1(n109541), .B2(n105641), .A(n94321), .ZN(
        \DLX_Datapath/RegisterFile/N26803 ) );
  NAND2_X1 U80088 ( .A1(n105211), .A2(n89153), .ZN(n94321) );
  OAI21_X1 U80089 ( .B1(n109079), .B2(n94297), .A(n94322), .ZN(
        \DLX_Datapath/RegisterFile/N26802 ) );
  NAND2_X1 U80090 ( .A1(n105211), .A2(n89271), .ZN(n94322) );
  OAI21_X1 U80091 ( .B1(n109426), .B2(n94297), .A(n94323), .ZN(
        \DLX_Datapath/RegisterFile/N26801 ) );
  NAND2_X1 U80092 ( .A1(n105211), .A2(n81792), .ZN(n94323) );
  OAI21_X1 U80093 ( .B1(n109307), .B2(n94297), .A(n94324), .ZN(
        \DLX_Datapath/RegisterFile/N26800 ) );
  NAND2_X1 U80094 ( .A1(n105211), .A2(n89506), .ZN(n94324) );
  OAI21_X1 U80095 ( .B1(n109199), .B2(n94297), .A(n94325), .ZN(
        \DLX_Datapath/RegisterFile/N26799 ) );
  NAND2_X1 U80096 ( .A1(n105211), .A2(n89624), .ZN(n94325) );
  OAI21_X1 U80097 ( .B1(n108734), .B2(n94297), .A(n94326), .ZN(
        \DLX_Datapath/RegisterFile/N26798 ) );
  NAND2_X1 U80098 ( .A1(n105211), .A2(n89742), .ZN(n94326) );
  OAI21_X1 U80099 ( .B1(n108962), .B2(n94297), .A(n94327), .ZN(
        \DLX_Datapath/RegisterFile/N26797 ) );
  NAND2_X1 U80100 ( .A1(n105211), .A2(n81790), .ZN(n94327) );
  OAI21_X1 U80101 ( .B1(n108850), .B2(n94297), .A(n94328), .ZN(
        \DLX_Datapath/RegisterFile/N26796 ) );
  NAND2_X1 U80102 ( .A1(n105211), .A2(n89977), .ZN(n94328) );
  OAI21_X1 U80103 ( .B1(n107167), .B2(n94297), .A(n94329), .ZN(
        \DLX_Datapath/RegisterFile/N26795 ) );
  NAND2_X1 U80104 ( .A1(n105211), .A2(n90096), .ZN(n94329) );
  NAND2_X1 U80105 ( .A1(n94294), .A2(n94330), .ZN(n94297) );
  NAND2_X1 U80106 ( .A1(n105137), .A2(n94331), .ZN(n94330) );
  AOI22_X1 U80107 ( .A1(n94333), .A2(n107944), .B1(n105639), .B2(n86303), .ZN(
        n94332) );
  AOI22_X1 U80108 ( .A1(n104983), .A2(n108040), .B1(n105639), .B2(n86558), 
        .ZN(n94335) );
  AOI22_X1 U80109 ( .A1(n94333), .A2(n107168), .B1(n105639), .B2(n86676), .ZN(
        n94336) );
  AOI22_X1 U80110 ( .A1(n104984), .A2(n107849), .B1(n105639), .B2(n86794), 
        .ZN(n94337) );
  AOI22_X1 U80111 ( .A1(n94333), .A2(n110744), .B1(n105639), .B2(n86912), .ZN(
        n94338) );
  AOI22_X1 U80112 ( .A1(n104983), .A2(n108149), .B1(n105639), .B2(n87030), 
        .ZN(n94339) );
  AOI22_X1 U80113 ( .A1(n104983), .A2(n110847), .B1(n105639), .B2(n87148), 
        .ZN(n94340) );
  AOI22_X1 U80114 ( .A1(n104984), .A2(n110948), .B1(n105639), .B2(n87266), 
        .ZN(n94341) );
  AOI22_X1 U80115 ( .A1(n104983), .A2(n110541), .B1(n105639), .B2(n87384), 
        .ZN(n94342) );
  AOI22_X1 U80116 ( .A1(n104983), .A2(n110326), .B1(n105638), .B2(n87502), 
        .ZN(n94343) );
  AOI22_X1 U80117 ( .A1(n104983), .A2(n110646), .B1(n105638), .B2(n87620), 
        .ZN(n94344) );
  AOI22_X1 U80118 ( .A1(n104984), .A2(n110435), .B1(n105638), .B2(n87738), 
        .ZN(n94345) );
  AOI22_X1 U80119 ( .A1(n104983), .A2(n110113), .B1(n105638), .B2(n87856), 
        .ZN(n94346) );
  AOI22_X1 U80120 ( .A1(n104984), .A2(n110220), .B1(n105638), .B2(n87974), 
        .ZN(n94347) );
  AOI22_X1 U80121 ( .A1(n104983), .A2(n110005), .B1(n105638), .B2(n88092), 
        .ZN(n94348) );
  AOI22_X1 U80122 ( .A1(n104984), .A2(n109888), .B1(n105638), .B2(n88210), 
        .ZN(n94349) );
  AOI22_X1 U80123 ( .A1(n104984), .A2(n108262), .B1(n105638), .B2(n88328), 
        .ZN(n94350) );
  AOI22_X1 U80124 ( .A1(n104983), .A2(n108385), .B1(n105638), .B2(n88446), 
        .ZN(n94351) );
  AOI22_X1 U80125 ( .A1(n104983), .A2(n108496), .B1(n105638), .B2(n88564), 
        .ZN(n94352) );
  AOI22_X1 U80126 ( .A1(n104983), .A2(n107733), .B1(n105638), .B2(n88682), 
        .ZN(n94353) );
  AOI22_X1 U80127 ( .A1(n104984), .A2(n109648), .B1(n105638), .B2(n88800), 
        .ZN(n94354) );
  AOI22_X1 U80128 ( .A1(n104984), .A2(n108610), .B1(n105639), .B2(n88918), 
        .ZN(n94355) );
  AOI22_X1 U80129 ( .A1(n104984), .A2(n109755), .B1(n105639), .B2(n81794), 
        .ZN(n94356) );
  AOI22_X1 U80130 ( .A1(n104983), .A2(n109540), .B1(n105639), .B2(n89153), 
        .ZN(n94357) );
  AOI22_X1 U80131 ( .A1(n104984), .A2(n109078), .B1(n94334), .B2(n89271), .ZN(
        n94358) );
  AOI22_X1 U80132 ( .A1(n104984), .A2(n109425), .B1(n105639), .B2(n81792), 
        .ZN(n94359) );
  AOI22_X1 U80133 ( .A1(n104984), .A2(n109306), .B1(n105638), .B2(n89506), 
        .ZN(n94360) );
  AOI22_X1 U80134 ( .A1(n104983), .A2(n109198), .B1(n105639), .B2(n89624), 
        .ZN(n94361) );
  AOI22_X1 U80135 ( .A1(n104983), .A2(n108733), .B1(n105639), .B2(n89742), 
        .ZN(n94362) );
  AOI22_X1 U80136 ( .A1(n104984), .A2(n108961), .B1(n105638), .B2(n81790), 
        .ZN(n94363) );
  AOI22_X1 U80137 ( .A1(n94333), .A2(n108849), .B1(n105639), .B2(n89977), .ZN(
        n94364) );
  AOI22_X1 U80138 ( .A1(n104984), .A2(n107169), .B1(n105638), .B2(n90096), 
        .ZN(n94365) );
  AOI21_X1 U80139 ( .B1(n94366), .B2(n105602), .A(n94334), .ZN(n94333) );
  AND2_X2 U80140 ( .A1(n105136), .A2(n94367), .ZN(n94334) );
  OAI21_X1 U80141 ( .B1(n105188), .B2(n104556), .A(n94368), .ZN(
        \DLX_Datapath/RegisterFile/N26762 ) );
  NAND2_X1 U80142 ( .A1(n105904), .A2(n86303), .ZN(n94368) );
  OAI21_X1 U80143 ( .B1(n105189), .B2(n104555), .A(n94369), .ZN(
        \DLX_Datapath/RegisterFile/N26761 ) );
  NAND2_X1 U80144 ( .A1(n105904), .A2(n86558), .ZN(n94369) );
  OAI21_X1 U80145 ( .B1(n105188), .B2(n104554), .A(n94370), .ZN(
        \DLX_Datapath/RegisterFile/N26760 ) );
  NAND2_X1 U80146 ( .A1(n105904), .A2(n86676), .ZN(n94370) );
  OAI21_X1 U80147 ( .B1(n105189), .B2(n104553), .A(n94371), .ZN(
        \DLX_Datapath/RegisterFile/N26759 ) );
  NAND2_X1 U80148 ( .A1(n105904), .A2(n86794), .ZN(n94371) );
  OAI21_X1 U80149 ( .B1(n105188), .B2(n104552), .A(n94372), .ZN(
        \DLX_Datapath/RegisterFile/N26758 ) );
  NAND2_X1 U80150 ( .A1(n105904), .A2(n86912), .ZN(n94372) );
  OAI21_X1 U80151 ( .B1(n105188), .B2(n104551), .A(n94373), .ZN(
        \DLX_Datapath/RegisterFile/N26757 ) );
  NAND2_X1 U80152 ( .A1(n105904), .A2(n87030), .ZN(n94373) );
  OAI21_X1 U80153 ( .B1(n105188), .B2(n104550), .A(n94374), .ZN(
        \DLX_Datapath/RegisterFile/N26756 ) );
  NAND2_X1 U80154 ( .A1(n105904), .A2(n87148), .ZN(n94374) );
  OAI21_X1 U80155 ( .B1(n105189), .B2(n104549), .A(n94375), .ZN(
        \DLX_Datapath/RegisterFile/N26755 ) );
  NAND2_X1 U80156 ( .A1(n105904), .A2(n87266), .ZN(n94375) );
  OAI21_X1 U80157 ( .B1(n105188), .B2(n104548), .A(n94376), .ZN(
        \DLX_Datapath/RegisterFile/N26754 ) );
  NAND2_X1 U80158 ( .A1(n105904), .A2(n87384), .ZN(n94376) );
  OAI21_X1 U80159 ( .B1(n106758), .B2(n104547), .A(n94377), .ZN(
        \DLX_Datapath/RegisterFile/N26753 ) );
  NAND2_X1 U80160 ( .A1(n105904), .A2(n87502), .ZN(n94377) );
  OAI21_X1 U80161 ( .B1(n106758), .B2(n104546), .A(n94378), .ZN(
        \DLX_Datapath/RegisterFile/N26752 ) );
  NAND2_X1 U80162 ( .A1(n105904), .A2(n87620), .ZN(n94378) );
  OAI21_X1 U80163 ( .B1(n106758), .B2(n104545), .A(n94379), .ZN(
        \DLX_Datapath/RegisterFile/N26751 ) );
  NAND2_X1 U80164 ( .A1(n105904), .A2(n87738), .ZN(n94379) );
  OAI21_X1 U80165 ( .B1(n106758), .B2(n104544), .A(n94380), .ZN(
        \DLX_Datapath/RegisterFile/N26750 ) );
  NAND2_X1 U80166 ( .A1(n105904), .A2(n87856), .ZN(n94380) );
  OAI21_X1 U80167 ( .B1(n106758), .B2(n104543), .A(n94381), .ZN(
        \DLX_Datapath/RegisterFile/N26749 ) );
  NAND2_X1 U80168 ( .A1(n105904), .A2(n87974), .ZN(n94381) );
  OAI21_X1 U80169 ( .B1(n106758), .B2(n104542), .A(n94382), .ZN(
        \DLX_Datapath/RegisterFile/N26748 ) );
  NAND2_X1 U80170 ( .A1(n105904), .A2(n88092), .ZN(n94382) );
  OAI21_X1 U80171 ( .B1(n106758), .B2(n104541), .A(n94383), .ZN(
        \DLX_Datapath/RegisterFile/N26747 ) );
  NAND2_X1 U80172 ( .A1(n105904), .A2(n88210), .ZN(n94383) );
  OAI21_X1 U80173 ( .B1(n105188), .B2(n104540), .A(n94384), .ZN(
        \DLX_Datapath/RegisterFile/N26746 ) );
  NAND2_X1 U80174 ( .A1(n105904), .A2(n88328), .ZN(n94384) );
  OAI21_X1 U80175 ( .B1(n105189), .B2(n104539), .A(n94385), .ZN(
        \DLX_Datapath/RegisterFile/N26745 ) );
  NAND2_X1 U80176 ( .A1(n105904), .A2(n88446), .ZN(n94385) );
  OAI21_X1 U80177 ( .B1(n105188), .B2(n104538), .A(n94386), .ZN(
        \DLX_Datapath/RegisterFile/N26744 ) );
  NAND2_X1 U80178 ( .A1(n81789), .A2(n88564), .ZN(n94386) );
  OAI21_X1 U80179 ( .B1(n105189), .B2(n104537), .A(n94387), .ZN(
        \DLX_Datapath/RegisterFile/N26743 ) );
  NAND2_X1 U80180 ( .A1(n81789), .A2(n88682), .ZN(n94387) );
  OAI21_X1 U80181 ( .B1(n105188), .B2(n104536), .A(n94388), .ZN(
        \DLX_Datapath/RegisterFile/N26742 ) );
  NAND2_X1 U80182 ( .A1(n81789), .A2(n88800), .ZN(n94388) );
  OAI21_X1 U80183 ( .B1(n105189), .B2(n104535), .A(n94389), .ZN(
        \DLX_Datapath/RegisterFile/N26741 ) );
  NAND2_X1 U80184 ( .A1(n81789), .A2(n88918), .ZN(n94389) );
  OAI21_X1 U80185 ( .B1(n105188), .B2(n104534), .A(n94390), .ZN(
        \DLX_Datapath/RegisterFile/N26739 ) );
  NAND2_X1 U80186 ( .A1(n81789), .A2(n89153), .ZN(n94390) );
  OAI21_X1 U80187 ( .B1(n105189), .B2(n104533), .A(n94391), .ZN(
        \DLX_Datapath/RegisterFile/N26738 ) );
  NAND2_X1 U80188 ( .A1(n81789), .A2(n89271), .ZN(n94391) );
  OAI21_X1 U80189 ( .B1(n105188), .B2(n104532), .A(n94392), .ZN(
        \DLX_Datapath/RegisterFile/N26736 ) );
  NAND2_X1 U80190 ( .A1(n81789), .A2(n89506), .ZN(n94392) );
  OAI21_X1 U80191 ( .B1(n105189), .B2(n104531), .A(n94393), .ZN(
        \DLX_Datapath/RegisterFile/N26735 ) );
  NAND2_X1 U80192 ( .A1(n81789), .A2(n89624), .ZN(n94393) );
  OAI21_X1 U80193 ( .B1(n105188), .B2(n104530), .A(n94394), .ZN(
        \DLX_Datapath/RegisterFile/N26734 ) );
  NAND2_X1 U80194 ( .A1(n81789), .A2(n89742), .ZN(n94394) );
  OAI21_X1 U80195 ( .B1(n105189), .B2(n104529), .A(n94395), .ZN(
        \DLX_Datapath/RegisterFile/N26732 ) );
  NAND2_X1 U80196 ( .A1(n81789), .A2(n89977), .ZN(n94395) );
  OAI21_X1 U80197 ( .B1(n105188), .B2(n104528), .A(n94396), .ZN(
        \DLX_Datapath/RegisterFile/N26731 ) );
  NAND2_X1 U80198 ( .A1(n81789), .A2(n90096), .ZN(n94396) );
  AOI21_X1 U80199 ( .B1(n94259), .B2(n94398), .A(n81789), .ZN(n94397) );
  AND2_X2 U80200 ( .A1(n105136), .A2(n94399), .ZN(n81789) );
  OAI21_X1 U80201 ( .B1(n103350), .B2(n94400), .A(n94401), .ZN(
        \DLX_Datapath/RegisterFile/N26730 ) );
  NAND2_X1 U80202 ( .A1(n107115), .A2(n86303), .ZN(n94401) );
  OAI21_X1 U80203 ( .B1(n103337), .B2(n94400), .A(n94402), .ZN(
        \DLX_Datapath/RegisterFile/N26729 ) );
  NAND2_X1 U80204 ( .A1(n107115), .A2(n86558), .ZN(n94402) );
  OAI21_X1 U80205 ( .B1(n103326), .B2(n94400), .A(n94403), .ZN(
        \DLX_Datapath/RegisterFile/N26728 ) );
  NAND2_X1 U80206 ( .A1(n107115), .A2(n86676), .ZN(n94403) );
  OAI21_X1 U80207 ( .B1(n103310), .B2(n94400), .A(n94404), .ZN(
        \DLX_Datapath/RegisterFile/N26727 ) );
  NAND2_X1 U80208 ( .A1(n107115), .A2(n86794), .ZN(n94404) );
  OAI21_X1 U80209 ( .B1(n103293), .B2(n94400), .A(n94405), .ZN(
        \DLX_Datapath/RegisterFile/N26726 ) );
  NAND2_X1 U80210 ( .A1(n107115), .A2(n86912), .ZN(n94405) );
  OAI21_X1 U80211 ( .B1(n103274), .B2(n94400), .A(n94406), .ZN(
        \DLX_Datapath/RegisterFile/N26725 ) );
  NAND2_X1 U80212 ( .A1(n107115), .A2(n87030), .ZN(n94406) );
  OAI21_X1 U80213 ( .B1(n103255), .B2(n94400), .A(n94407), .ZN(
        \DLX_Datapath/RegisterFile/N26724 ) );
  NAND2_X1 U80214 ( .A1(n107115), .A2(n87148), .ZN(n94407) );
  OAI21_X1 U80215 ( .B1(n103236), .B2(n94400), .A(n94408), .ZN(
        \DLX_Datapath/RegisterFile/N26723 ) );
  NAND2_X1 U80216 ( .A1(n107115), .A2(n87266), .ZN(n94408) );
  OAI21_X1 U80217 ( .B1(n103217), .B2(n105637), .A(n94409), .ZN(
        \DLX_Datapath/RegisterFile/N26722 ) );
  NAND2_X1 U80218 ( .A1(n105210), .A2(n87384), .ZN(n94409) );
  OAI21_X1 U80219 ( .B1(n103199), .B2(n105637), .A(n94410), .ZN(
        \DLX_Datapath/RegisterFile/N26721 ) );
  NAND2_X1 U80220 ( .A1(n105210), .A2(n87502), .ZN(n94410) );
  OAI21_X1 U80221 ( .B1(n103180), .B2(n105637), .A(n94411), .ZN(
        \DLX_Datapath/RegisterFile/N26720 ) );
  NAND2_X1 U80222 ( .A1(n105210), .A2(n87620), .ZN(n94411) );
  OAI21_X1 U80223 ( .B1(n103161), .B2(n105637), .A(n94412), .ZN(
        \DLX_Datapath/RegisterFile/N26719 ) );
  NAND2_X1 U80224 ( .A1(n105210), .A2(n87738), .ZN(n94412) );
  OAI21_X1 U80225 ( .B1(n103141), .B2(n105637), .A(n94413), .ZN(
        \DLX_Datapath/RegisterFile/N26718 ) );
  NAND2_X1 U80226 ( .A1(n105210), .A2(n87856), .ZN(n94413) );
  OAI21_X1 U80227 ( .B1(n103123), .B2(n105637), .A(n94414), .ZN(
        \DLX_Datapath/RegisterFile/N26717 ) );
  NAND2_X1 U80228 ( .A1(n105210), .A2(n87974), .ZN(n94414) );
  OAI21_X1 U80229 ( .B1(n103103), .B2(n105637), .A(n94415), .ZN(
        \DLX_Datapath/RegisterFile/N26716 ) );
  NAND2_X1 U80230 ( .A1(n105210), .A2(n88092), .ZN(n94415) );
  OAI21_X1 U80231 ( .B1(n103083), .B2(n105637), .A(n94416), .ZN(
        \DLX_Datapath/RegisterFile/N26715 ) );
  NAND2_X1 U80232 ( .A1(n105210), .A2(n88210), .ZN(n94416) );
  OAI21_X1 U80233 ( .B1(n103063), .B2(n105637), .A(n94417), .ZN(
        \DLX_Datapath/RegisterFile/N26714 ) );
  NAND2_X1 U80234 ( .A1(n105210), .A2(n88328), .ZN(n94417) );
  OAI21_X1 U80235 ( .B1(n103043), .B2(n105637), .A(n94418), .ZN(
        \DLX_Datapath/RegisterFile/N26713 ) );
  NAND2_X1 U80236 ( .A1(n105210), .A2(n88446), .ZN(n94418) );
  OAI21_X1 U80237 ( .B1(n103023), .B2(n105637), .A(n94419), .ZN(
        \DLX_Datapath/RegisterFile/N26712 ) );
  NAND2_X1 U80238 ( .A1(n105210), .A2(n88564), .ZN(n94419) );
  OAI21_X1 U80239 ( .B1(n103003), .B2(n105637), .A(n94420), .ZN(
        \DLX_Datapath/RegisterFile/N26711 ) );
  NAND2_X1 U80240 ( .A1(n105210), .A2(n88682), .ZN(n94420) );
  OAI21_X1 U80241 ( .B1(n102983), .B2(n105636), .A(n94421), .ZN(
        \DLX_Datapath/RegisterFile/N26710 ) );
  NAND2_X1 U80242 ( .A1(n105209), .A2(n88800), .ZN(n94421) );
  OAI21_X1 U80243 ( .B1(n102966), .B2(n105636), .A(n94422), .ZN(
        \DLX_Datapath/RegisterFile/N26709 ) );
  NAND2_X1 U80244 ( .A1(n105209), .A2(n88918), .ZN(n94422) );
  OAI21_X1 U80245 ( .B1(n102946), .B2(n105636), .A(n94423), .ZN(
        \DLX_Datapath/RegisterFile/N26708 ) );
  NAND2_X1 U80246 ( .A1(n105209), .A2(n81794), .ZN(n94423) );
  OAI21_X1 U80247 ( .B1(n102926), .B2(n105636), .A(n94424), .ZN(
        \DLX_Datapath/RegisterFile/N26707 ) );
  NAND2_X1 U80248 ( .A1(n105209), .A2(n89153), .ZN(n94424) );
  OAI21_X1 U80249 ( .B1(n102906), .B2(n105636), .A(n94425), .ZN(
        \DLX_Datapath/RegisterFile/N26706 ) );
  NAND2_X1 U80250 ( .A1(n105209), .A2(n89271), .ZN(n94425) );
  OAI21_X1 U80251 ( .B1(n102886), .B2(n105636), .A(n94426), .ZN(
        \DLX_Datapath/RegisterFile/N26705 ) );
  NAND2_X1 U80252 ( .A1(n105209), .A2(n81792), .ZN(n94426) );
  OAI21_X1 U80253 ( .B1(n102866), .B2(n105636), .A(n94427), .ZN(
        \DLX_Datapath/RegisterFile/N26704 ) );
  NAND2_X1 U80254 ( .A1(n105209), .A2(n89506), .ZN(n94427) );
  OAI21_X1 U80255 ( .B1(n102846), .B2(n105636), .A(n94428), .ZN(
        \DLX_Datapath/RegisterFile/N26703 ) );
  NAND2_X1 U80256 ( .A1(n105209), .A2(n89624), .ZN(n94428) );
  OAI21_X1 U80257 ( .B1(n102826), .B2(n105636), .A(n94429), .ZN(
        \DLX_Datapath/RegisterFile/N26702 ) );
  NAND2_X1 U80258 ( .A1(n105209), .A2(n89742), .ZN(n94429) );
  OAI21_X1 U80259 ( .B1(n102806), .B2(n105636), .A(n94430), .ZN(
        \DLX_Datapath/RegisterFile/N26701 ) );
  NAND2_X1 U80260 ( .A1(n105209), .A2(n81790), .ZN(n94430) );
  OAI21_X1 U80261 ( .B1(n102786), .B2(n105636), .A(n94431), .ZN(
        \DLX_Datapath/RegisterFile/N26700 ) );
  NAND2_X1 U80262 ( .A1(n105209), .A2(n89977), .ZN(n94431) );
  OAI21_X1 U80263 ( .B1(n102766), .B2(n105636), .A(n94432), .ZN(
        \DLX_Datapath/RegisterFile/N26699 ) );
  NAND2_X1 U80264 ( .A1(n105209), .A2(n90096), .ZN(n94432) );
  NAND2_X1 U80265 ( .A1(n94294), .A2(n94433), .ZN(n94400) );
  NAND2_X1 U80266 ( .A1(n105137), .A2(n94434), .ZN(n94433) );
  OAI21_X1 U80267 ( .B1(n102747), .B2(n94435), .A(n94436), .ZN(
        \DLX_Datapath/RegisterFile/N26698 ) );
  NAND2_X1 U80268 ( .A1(n107113), .A2(n86303), .ZN(n94436) );
  OAI21_X1 U80269 ( .B1(n102734), .B2(n94435), .A(n94437), .ZN(
        \DLX_Datapath/RegisterFile/N26697 ) );
  NAND2_X1 U80270 ( .A1(n107113), .A2(n86558), .ZN(n94437) );
  OAI21_X1 U80271 ( .B1(n102718), .B2(n94435), .A(n94438), .ZN(
        \DLX_Datapath/RegisterFile/N26696 ) );
  NAND2_X1 U80272 ( .A1(n107113), .A2(n86676), .ZN(n94438) );
  OAI21_X1 U80273 ( .B1(n102702), .B2(n94435), .A(n94439), .ZN(
        \DLX_Datapath/RegisterFile/N26695 ) );
  NAND2_X1 U80274 ( .A1(n107113), .A2(n86794), .ZN(n94439) );
  OAI21_X1 U80275 ( .B1(n102688), .B2(n94435), .A(n94440), .ZN(
        \DLX_Datapath/RegisterFile/N26694 ) );
  NAND2_X1 U80276 ( .A1(n107113), .A2(n86912), .ZN(n94440) );
  OAI21_X1 U80277 ( .B1(n102673), .B2(n94435), .A(n94441), .ZN(
        \DLX_Datapath/RegisterFile/N26693 ) );
  NAND2_X1 U80278 ( .A1(n107113), .A2(n87030), .ZN(n94441) );
  OAI21_X1 U80279 ( .B1(n102655), .B2(n94435), .A(n94442), .ZN(
        \DLX_Datapath/RegisterFile/N26692 ) );
  NAND2_X1 U80280 ( .A1(n107113), .A2(n87148), .ZN(n94442) );
  OAI21_X1 U80281 ( .B1(n102639), .B2(n94435), .A(n94443), .ZN(
        \DLX_Datapath/RegisterFile/N26691 ) );
  NAND2_X1 U80282 ( .A1(n107113), .A2(n87266), .ZN(n94443) );
  OAI21_X1 U80283 ( .B1(n102622), .B2(n105635), .A(n94444), .ZN(
        \DLX_Datapath/RegisterFile/N26690 ) );
  NAND2_X1 U80284 ( .A1(n105208), .A2(n87384), .ZN(n94444) );
  OAI21_X1 U80285 ( .B1(n102608), .B2(n105635), .A(n94445), .ZN(
        \DLX_Datapath/RegisterFile/N26689 ) );
  NAND2_X1 U80286 ( .A1(n105208), .A2(n87502), .ZN(n94445) );
  OAI21_X1 U80287 ( .B1(n102593), .B2(n105635), .A(n94446), .ZN(
        \DLX_Datapath/RegisterFile/N26688 ) );
  NAND2_X1 U80288 ( .A1(n105208), .A2(n87620), .ZN(n94446) );
  OAI21_X1 U80289 ( .B1(n102578), .B2(n105635), .A(n94447), .ZN(
        \DLX_Datapath/RegisterFile/N26687 ) );
  NAND2_X1 U80290 ( .A1(n105208), .A2(n87738), .ZN(n94447) );
  OAI21_X1 U80291 ( .B1(n102562), .B2(n105635), .A(n94448), .ZN(
        \DLX_Datapath/RegisterFile/N26686 ) );
  NAND2_X1 U80292 ( .A1(n105208), .A2(n87856), .ZN(n94448) );
  OAI21_X1 U80293 ( .B1(n102545), .B2(n105635), .A(n94449), .ZN(
        \DLX_Datapath/RegisterFile/N26685 ) );
  NAND2_X1 U80294 ( .A1(n105208), .A2(n87974), .ZN(n94449) );
  OAI21_X1 U80295 ( .B1(n102528), .B2(n105635), .A(n94450), .ZN(
        \DLX_Datapath/RegisterFile/N26684 ) );
  NAND2_X1 U80296 ( .A1(n105208), .A2(n88092), .ZN(n94450) );
  OAI21_X1 U80297 ( .B1(n102509), .B2(n105635), .A(n94451), .ZN(
        \DLX_Datapath/RegisterFile/N26683 ) );
  NAND2_X1 U80298 ( .A1(n105208), .A2(n88210), .ZN(n94451) );
  OAI21_X1 U80299 ( .B1(n102491), .B2(n105635), .A(n94452), .ZN(
        \DLX_Datapath/RegisterFile/N26682 ) );
  NAND2_X1 U80300 ( .A1(n105208), .A2(n88328), .ZN(n94452) );
  OAI21_X1 U80301 ( .B1(n102473), .B2(n105635), .A(n94453), .ZN(
        \DLX_Datapath/RegisterFile/N26681 ) );
  NAND2_X1 U80302 ( .A1(n105208), .A2(n88446), .ZN(n94453) );
  OAI21_X1 U80303 ( .B1(n102453), .B2(n105635), .A(n94454), .ZN(
        \DLX_Datapath/RegisterFile/N26680 ) );
  NAND2_X1 U80304 ( .A1(n105208), .A2(n88564), .ZN(n94454) );
  OAI21_X1 U80305 ( .B1(n102435), .B2(n105635), .A(n94455), .ZN(
        \DLX_Datapath/RegisterFile/N26679 ) );
  NAND2_X1 U80306 ( .A1(n105208), .A2(n88682), .ZN(n94455) );
  OAI21_X1 U80307 ( .B1(n102415), .B2(n105634), .A(n94456), .ZN(
        \DLX_Datapath/RegisterFile/N26678 ) );
  NAND2_X1 U80308 ( .A1(n105207), .A2(n88800), .ZN(n94456) );
  OAI21_X1 U80309 ( .B1(n102395), .B2(n105634), .A(n94457), .ZN(
        \DLX_Datapath/RegisterFile/N26677 ) );
  NAND2_X1 U80310 ( .A1(n105207), .A2(n88918), .ZN(n94457) );
  OAI21_X1 U80311 ( .B1(n102375), .B2(n105634), .A(n94458), .ZN(
        \DLX_Datapath/RegisterFile/N26676 ) );
  NAND2_X1 U80312 ( .A1(n105207), .A2(n81794), .ZN(n94458) );
  OAI21_X1 U80313 ( .B1(n102357), .B2(n105634), .A(n94459), .ZN(
        \DLX_Datapath/RegisterFile/N26675 ) );
  NAND2_X1 U80314 ( .A1(n105207), .A2(n89153), .ZN(n94459) );
  OAI21_X1 U80315 ( .B1(n102337), .B2(n105634), .A(n94460), .ZN(
        \DLX_Datapath/RegisterFile/N26674 ) );
  NAND2_X1 U80316 ( .A1(n105207), .A2(n89271), .ZN(n94460) );
  OAI21_X1 U80317 ( .B1(n102317), .B2(n105634), .A(n94461), .ZN(
        \DLX_Datapath/RegisterFile/N26673 ) );
  NAND2_X1 U80318 ( .A1(n105207), .A2(n81792), .ZN(n94461) );
  OAI21_X1 U80319 ( .B1(n102297), .B2(n105634), .A(n94462), .ZN(
        \DLX_Datapath/RegisterFile/N26672 ) );
  NAND2_X1 U80320 ( .A1(n105207), .A2(n89506), .ZN(n94462) );
  OAI21_X1 U80321 ( .B1(n102278), .B2(n105634), .A(n94463), .ZN(
        \DLX_Datapath/RegisterFile/N26671 ) );
  NAND2_X1 U80322 ( .A1(n105207), .A2(n89624), .ZN(n94463) );
  OAI21_X1 U80323 ( .B1(n102258), .B2(n105634), .A(n94464), .ZN(
        \DLX_Datapath/RegisterFile/N26670 ) );
  NAND2_X1 U80324 ( .A1(n105207), .A2(n89742), .ZN(n94464) );
  OAI21_X1 U80325 ( .B1(n102239), .B2(n105634), .A(n94465), .ZN(
        \DLX_Datapath/RegisterFile/N26669 ) );
  NAND2_X1 U80326 ( .A1(n105207), .A2(n81790), .ZN(n94465) );
  OAI21_X1 U80327 ( .B1(n102219), .B2(n105634), .A(n94466), .ZN(
        \DLX_Datapath/RegisterFile/N26668 ) );
  NAND2_X1 U80328 ( .A1(n105207), .A2(n89977), .ZN(n94466) );
  OAI21_X1 U80329 ( .B1(n102199), .B2(n105634), .A(n94467), .ZN(
        \DLX_Datapath/RegisterFile/N26667 ) );
  NAND2_X1 U80330 ( .A1(n105207), .A2(n90096), .ZN(n94467) );
  NAND2_X1 U80331 ( .A1(n94294), .A2(n94468), .ZN(n94435) );
  NAND2_X1 U80332 ( .A1(n94469), .A2(n105136), .ZN(n94468) );
  NOR2_X1 U80333 ( .A1(n94470), .A2(n94093), .ZN(n94469) );
  NAND2_X1 U80334 ( .A1(n105602), .A2(n94366), .ZN(n94294) );
  AOI22_X1 U80335 ( .A1(n104985), .A2(n107941), .B1(n105633), .B2(n86303), 
        .ZN(n94471) );
  AOI22_X1 U80336 ( .A1(n104985), .A2(n108037), .B1(n105633), .B2(n86558), 
        .ZN(n94474) );
  AOI22_X1 U80337 ( .A1(n104985), .A2(n107174), .B1(n105633), .B2(n86676), 
        .ZN(n94475) );
  AOI22_X1 U80338 ( .A1(n104986), .A2(n107846), .B1(n105633), .B2(n86794), 
        .ZN(n94476) );
  AOI22_X1 U80339 ( .A1(n104985), .A2(n110741), .B1(n105633), .B2(n86912), 
        .ZN(n94477) );
  AOI22_X1 U80340 ( .A1(n104986), .A2(n108146), .B1(n105633), .B2(n87030), 
        .ZN(n94478) );
  AOI22_X1 U80341 ( .A1(n104986), .A2(n110844), .B1(n105633), .B2(n87148), 
        .ZN(n94479) );
  AOI22_X1 U80342 ( .A1(n104986), .A2(n110945), .B1(n105633), .B2(n87266), 
        .ZN(n94480) );
  AOI22_X1 U80343 ( .A1(n104985), .A2(n110538), .B1(n105633), .B2(n87384), 
        .ZN(n94481) );
  AOI22_X1 U80344 ( .A1(n94472), .A2(n110323), .B1(n105632), .B2(n87502), .ZN(
        n94482) );
  AOI22_X1 U80345 ( .A1(n94472), .A2(n110643), .B1(n105632), .B2(n87620), .ZN(
        n94483) );
  AOI22_X1 U80346 ( .A1(n104986), .A2(n110432), .B1(n105632), .B2(n87738), 
        .ZN(n94484) );
  AOI22_X1 U80347 ( .A1(n104985), .A2(n110110), .B1(n105632), .B2(n87856), 
        .ZN(n94485) );
  AOI22_X1 U80348 ( .A1(n104986), .A2(n110217), .B1(n105632), .B2(n87974), 
        .ZN(n94486) );
  AOI22_X1 U80349 ( .A1(n94472), .A2(n110002), .B1(n105632), .B2(n88092), .ZN(
        n94487) );
  AOI22_X1 U80350 ( .A1(n104986), .A2(n109885), .B1(n105632), .B2(n88210), 
        .ZN(n94488) );
  AOI22_X1 U80351 ( .A1(n104985), .A2(n108259), .B1(n105632), .B2(n88328), 
        .ZN(n94489) );
  AOI22_X1 U80352 ( .A1(n104985), .A2(n108382), .B1(n105632), .B2(n88446), 
        .ZN(n94490) );
  AOI22_X1 U80353 ( .A1(n104985), .A2(n108493), .B1(n105632), .B2(n88564), 
        .ZN(n94491) );
  AOI22_X1 U80354 ( .A1(n94472), .A2(n107730), .B1(n105632), .B2(n88682), .ZN(
        n94492) );
  AOI22_X1 U80355 ( .A1(n104986), .A2(n109645), .B1(n105632), .B2(n88800), 
        .ZN(n94493) );
  AOI22_X1 U80356 ( .A1(n104985), .A2(n108607), .B1(n105633), .B2(n88918), 
        .ZN(n94494) );
  AOI22_X1 U80357 ( .A1(n104986), .A2(n109752), .B1(n105633), .B2(n81794), 
        .ZN(n94495) );
  AOI22_X1 U80358 ( .A1(n104986), .A2(n109537), .B1(n105633), .B2(n89153), 
        .ZN(n94496) );
  AOI22_X1 U80359 ( .A1(n104986), .A2(n109075), .B1(n94473), .B2(n89271), .ZN(
        n94497) );
  AOI22_X1 U80360 ( .A1(n104985), .A2(n109422), .B1(n105633), .B2(n81792), 
        .ZN(n94498) );
  AOI22_X1 U80361 ( .A1(n104985), .A2(n109303), .B1(n105632), .B2(n89506), 
        .ZN(n94499) );
  AOI22_X1 U80362 ( .A1(n104985), .A2(n109195), .B1(n105633), .B2(n89624), 
        .ZN(n94500) );
  AOI22_X1 U80363 ( .A1(n104986), .A2(n108730), .B1(n105633), .B2(n89742), 
        .ZN(n94501) );
  AOI22_X1 U80364 ( .A1(n104986), .A2(n108958), .B1(n105632), .B2(n81790), 
        .ZN(n94502) );
  AOI22_X1 U80365 ( .A1(n104985), .A2(n108846), .B1(n105633), .B2(n89977), 
        .ZN(n94503) );
  AOI22_X1 U80366 ( .A1(n104986), .A2(n107175), .B1(n105632), .B2(n90096), 
        .ZN(n94504) );
  AOI21_X1 U80367 ( .B1(n94366), .B2(n105602), .A(n94473), .ZN(n94472) );
  AND2_X2 U80368 ( .A1(n105136), .A2(n94505), .ZN(n94473) );
  OAI21_X1 U80369 ( .B1(n107371), .B2(n105630), .A(n94507), .ZN(
        \DLX_Datapath/RegisterFile/N26634 ) );
  AOI22_X1 U80370 ( .A1(n105628), .A2(n107940), .B1(n104714), .B2(n81360), 
        .ZN(n94507) );
  OAI21_X1 U80371 ( .B1(n107373), .B2(n105629), .A(n94510), .ZN(
        \DLX_Datapath/RegisterFile/N26633 ) );
  AOI22_X1 U80372 ( .A1(n105628), .A2(n108036), .B1(n94511), .B2(n104715), 
        .ZN(n94510) );
  OAI21_X1 U80373 ( .B1(n106832), .B2(n105629), .A(n94512), .ZN(
        \DLX_Datapath/RegisterFile/N26632 ) );
  AOI22_X1 U80374 ( .A1(n105628), .A2(n107176), .B1(n104715), .B2(n81539), 
        .ZN(n94512) );
  OAI21_X1 U80375 ( .B1(n107376), .B2(n105630), .A(n94513), .ZN(
        \DLX_Datapath/RegisterFile/N26631 ) );
  AOI22_X1 U80376 ( .A1(n105628), .A2(n107845), .B1(n104716), .B2(n81301), 
        .ZN(n94513) );
  OAI21_X1 U80377 ( .B1(n107378), .B2(n105629), .A(n94514), .ZN(
        \DLX_Datapath/RegisterFile/N26630 ) );
  AOI22_X1 U80378 ( .A1(n105628), .A2(n110740), .B1(n104714), .B2(n81308), 
        .ZN(n94514) );
  OAI21_X1 U80379 ( .B1(n107380), .B2(n105630), .A(n94515), .ZN(
        \DLX_Datapath/RegisterFile/N26629 ) );
  AOI22_X1 U80380 ( .A1(n105628), .A2(n108145), .B1(n94516), .B2(n104716), 
        .ZN(n94515) );
  OAI21_X1 U80381 ( .B1(n107382), .B2(n105630), .A(n94517), .ZN(
        \DLX_Datapath/RegisterFile/N26628 ) );
  AOI22_X1 U80382 ( .A1(n105628), .A2(n110843), .B1(n104716), .B2(n81272), 
        .ZN(n94517) );
  OAI21_X1 U80383 ( .B1(n107384), .B2(n105629), .A(n94518), .ZN(
        \DLX_Datapath/RegisterFile/N26627 ) );
  AOI22_X1 U80384 ( .A1(n105628), .A2(n110944), .B1(n94519), .B2(n104714), 
        .ZN(n94518) );
  OAI21_X1 U80385 ( .B1(n107386), .B2(n105629), .A(n94520), .ZN(
        \DLX_Datapath/RegisterFile/N26626 ) );
  AOI22_X1 U80386 ( .A1(n105627), .A2(n110537), .B1(n104716), .B2(n80192), 
        .ZN(n94520) );
  OAI21_X1 U80387 ( .B1(n107388), .B2(n105630), .A(n94521), .ZN(
        \DLX_Datapath/RegisterFile/N26625 ) );
  AOI22_X1 U80388 ( .A1(n105627), .A2(n110322), .B1(n104716), .B2(n81474), 
        .ZN(n94521) );
  OAI21_X1 U80389 ( .B1(n107390), .B2(n105630), .A(n94522), .ZN(
        \DLX_Datapath/RegisterFile/N26624 ) );
  AOI22_X1 U80390 ( .A1(n105627), .A2(n110642), .B1(n94523), .B2(n104715), 
        .ZN(n94522) );
  AOI22_X1 U80392 ( .A1(n94508), .A2(n110431), .B1(n104716), .B2(n106061), 
        .ZN(n94524) );
  OAI21_X1 U80393 ( .B1(n107394), .B2(n105630), .A(n94525), .ZN(
        \DLX_Datapath/RegisterFile/N26622 ) );
  AOI22_X1 U80394 ( .A1(n105627), .A2(n110109), .B1(n104716), .B2(n81347), 
        .ZN(n94525) );
  OAI21_X1 U80395 ( .B1(n107396), .B2(n105630), .A(n94526), .ZN(
        \DLX_Datapath/RegisterFile/N26621 ) );
  AOI22_X1 U80396 ( .A1(n105627), .A2(n110216), .B1(n94527), .B2(n104714), 
        .ZN(n94526) );
  OAI21_X1 U80397 ( .B1(n107398), .B2(n105629), .A(n94528), .ZN(
        \DLX_Datapath/RegisterFile/N26620 ) );
  AOI22_X1 U80398 ( .A1(n105627), .A2(n110001), .B1(n104714), .B2(n81297), 
        .ZN(n94528) );
  AOI22_X1 U80400 ( .A1(n105628), .A2(n109884), .B1(n94530), .B2(n104714), 
        .ZN(n94529) );
  OAI21_X1 U80401 ( .B1(n107402), .B2(n105630), .A(n94531), .ZN(
        \DLX_Datapath/RegisterFile/N26618 ) );
  AOI22_X1 U80402 ( .A1(n105627), .A2(n108258), .B1(n104715), .B2(n81286), 
        .ZN(n94531) );
  OAI21_X1 U80403 ( .B1(n107404), .B2(n105629), .A(n94532), .ZN(
        \DLX_Datapath/RegisterFile/N26617 ) );
  AOI22_X1 U80404 ( .A1(n105627), .A2(n108381), .B1(n104715), .B2(n106169), 
        .ZN(n94532) );
  AOI22_X1 U80406 ( .A1(n105628), .A2(n108492), .B1(n104714), .B2(n81283), 
        .ZN(n94533) );
  OAI21_X1 U80407 ( .B1(n107408), .B2(n105630), .A(n94534), .ZN(
        \DLX_Datapath/RegisterFile/N26615 ) );
  AOI22_X1 U80408 ( .A1(n105627), .A2(n107729), .B1(n104714), .B2(n81453), 
        .ZN(n94534) );
  OAI21_X1 U80409 ( .B1(n107410), .B2(n105629), .A(n94535), .ZN(
        \DLX_Datapath/RegisterFile/N26614 ) );
  AOI22_X1 U80410 ( .A1(n105627), .A2(n109644), .B1(n94536), .B2(n104716), 
        .ZN(n94535) );
  AOI22_X1 U80412 ( .A1(n105627), .A2(n108606), .B1(n104715), .B2(n106241), 
        .ZN(n94537) );
  OAI21_X1 U80413 ( .B1(n107367), .B2(n105629), .A(n94538), .ZN(
        \DLX_Datapath/RegisterFile/N26612 ) );
  AOI22_X1 U80414 ( .A1(n105627), .A2(n109751), .B1(n104716), .B2(n81351), 
        .ZN(n94538) );
  OAI21_X1 U80415 ( .B1(n107369), .B2(n105630), .A(n94539), .ZN(
        \DLX_Datapath/RegisterFile/N26611 ) );
  AOI22_X1 U80416 ( .A1(n105627), .A2(n109536), .B1(n104715), .B2(n106020), 
        .ZN(n94539) );
  OAI21_X1 U80417 ( .B1(n108974), .B2(n105630), .A(n94540), .ZN(
        \DLX_Datapath/RegisterFile/N26610 ) );
  AOI22_X1 U80418 ( .A1(n105627), .A2(n109074), .B1(n94541), .B2(n104715), 
        .ZN(n94540) );
  OAI21_X1 U80419 ( .B1(n111063), .B2(n105629), .A(n94542), .ZN(
        \DLX_Datapath/RegisterFile/N26609 ) );
  AOI22_X1 U80420 ( .A1(n105627), .A2(n109421), .B1(n104714), .B2(n81269), 
        .ZN(n94542) );
  OAI21_X1 U80421 ( .B1(n111062), .B2(n105630), .A(n94543), .ZN(
        \DLX_Datapath/RegisterFile/N26608 ) );
  AOI22_X1 U80422 ( .A1(n105627), .A2(n109302), .B1(n105625), .B2(n104714), 
        .ZN(n94543) );
  OAI21_X1 U80423 ( .B1(n111061), .B2(n105630), .A(n94545), .ZN(
        \DLX_Datapath/RegisterFile/N26607 ) );
  AOI22_X1 U80424 ( .A1(n105627), .A2(n109194), .B1(n94546), .B2(n104714), 
        .ZN(n94545) );
  OAI21_X1 U80425 ( .B1(n111060), .B2(n105629), .A(n94547), .ZN(
        \DLX_Datapath/RegisterFile/N26606 ) );
  AOI22_X1 U80426 ( .A1(n105627), .A2(n108729), .B1(n94548), .B2(n104716), 
        .ZN(n94547) );
  OAI21_X1 U80427 ( .B1(n111059), .B2(n105629), .A(n94549), .ZN(
        \DLX_Datapath/RegisterFile/N26605 ) );
  AOI22_X1 U80428 ( .A1(n105627), .A2(n108957), .B1(n104715), .B2(n81783), 
        .ZN(n94549) );
  AOI22_X1 U80430 ( .A1(n105627), .A2(n108845), .B1(n104716), .B2(n80188), 
        .ZN(n94550) );
  OAI21_X1 U80431 ( .B1(n111057), .B2(n105629), .A(n94551), .ZN(
        \DLX_Datapath/RegisterFile/N26603 ) );
  AOI22_X1 U80432 ( .A1(n105627), .A2(n107177), .B1(n104715), .B2(n81265), 
        .ZN(n94551) );
  NOR2_X1 U80433 ( .A1(n94552), .A2(n94553), .ZN(n94509) );
  NAND2_X1 U80434 ( .A1(n94506), .A2(n111026), .ZN(n94552) );
  AOI21_X1 U80435 ( .B1(n94259), .B2(n94554), .A(n105631), .ZN(n94508) );
  NAND2_X1 U80436 ( .A1(n105137), .A2(n94555), .ZN(n94506) );
  OAI21_X1 U80437 ( .B1(n107371), .B2(n105619), .A(n94557), .ZN(
        \DLX_Datapath/RegisterFile/N26602 ) );
  AOI22_X1 U80438 ( .A1(n105617), .A2(n107939), .B1(n94559), .B2(n105614), 
        .ZN(n94557) );
  OAI21_X1 U80439 ( .B1(n107373), .B2(n105618), .A(n94561), .ZN(
        \DLX_Datapath/RegisterFile/N26601 ) );
  AOI22_X1 U80440 ( .A1(n105617), .A2(n108035), .B1(n94562), .B2(n105613), 
        .ZN(n94561) );
  OAI21_X1 U80441 ( .B1(n106832), .B2(n105619), .A(n94563), .ZN(
        \DLX_Datapath/RegisterFile/N26600 ) );
  AOI22_X1 U80442 ( .A1(n105617), .A2(n107178), .B1(n94564), .B2(n105614), 
        .ZN(n94563) );
  OAI21_X1 U80443 ( .B1(n107376), .B2(n105618), .A(n94565), .ZN(
        \DLX_Datapath/RegisterFile/N26599 ) );
  AOI22_X1 U80444 ( .A1(n105617), .A2(n107844), .B1(n94566), .B2(n105613), 
        .ZN(n94565) );
  OAI21_X1 U80445 ( .B1(n107378), .B2(n105619), .A(n94567), .ZN(
        \DLX_Datapath/RegisterFile/N26598 ) );
  AOI22_X1 U80446 ( .A1(n105617), .A2(n110739), .B1(n94568), .B2(n105614), 
        .ZN(n94567) );
  OAI21_X1 U80447 ( .B1(n107380), .B2(n105618), .A(n94569), .ZN(
        \DLX_Datapath/RegisterFile/N26597 ) );
  AOI22_X1 U80448 ( .A1(n105617), .A2(n108144), .B1(n94570), .B2(n105613), 
        .ZN(n94569) );
  OAI21_X1 U80449 ( .B1(n107382), .B2(n105619), .A(n94571), .ZN(
        \DLX_Datapath/RegisterFile/N26596 ) );
  AOI22_X1 U80450 ( .A1(n105617), .A2(n110842), .B1(n94572), .B2(n105614), 
        .ZN(n94571) );
  OAI21_X1 U80451 ( .B1(n107384), .B2(n105618), .A(n94573), .ZN(
        \DLX_Datapath/RegisterFile/N26595 ) );
  AOI22_X1 U80452 ( .A1(n105617), .A2(n110943), .B1(n94574), .B2(n105613), 
        .ZN(n94573) );
  OAI21_X1 U80453 ( .B1(n107386), .B2(n105619), .A(n94575), .ZN(
        \DLX_Datapath/RegisterFile/N26594 ) );
  AOI22_X1 U80454 ( .A1(n105616), .A2(n110536), .B1(n94576), .B2(n105613), 
        .ZN(n94575) );
  OAI21_X1 U80455 ( .B1(n107388), .B2(n105619), .A(n94577), .ZN(
        \DLX_Datapath/RegisterFile/N26593 ) );
  AOI22_X1 U80456 ( .A1(n105616), .A2(n110321), .B1(n94578), .B2(n105614), 
        .ZN(n94577) );
  OAI21_X1 U80457 ( .B1(n107390), .B2(n105618), .A(n94579), .ZN(
        \DLX_Datapath/RegisterFile/N26592 ) );
  AOI22_X1 U80458 ( .A1(n105616), .A2(n110641), .B1(n94580), .B2(n105613), 
        .ZN(n94579) );
  OAI21_X1 U80459 ( .B1(n107392), .B2(n105618), .A(n94581), .ZN(
        \DLX_Datapath/RegisterFile/N26591 ) );
  AOI22_X1 U80460 ( .A1(n105616), .A2(n110430), .B1(n94582), .B2(n105614), 
        .ZN(n94581) );
  OAI21_X1 U80461 ( .B1(n107394), .B2(n105619), .A(n94583), .ZN(
        \DLX_Datapath/RegisterFile/N26590 ) );
  AOI22_X1 U80462 ( .A1(n105616), .A2(n110108), .B1(n94584), .B2(n105613), 
        .ZN(n94583) );
  OAI21_X1 U80463 ( .B1(n107396), .B2(n105618), .A(n94585), .ZN(
        \DLX_Datapath/RegisterFile/N26589 ) );
  AOI22_X1 U80464 ( .A1(n105616), .A2(n110215), .B1(n94586), .B2(n105614), 
        .ZN(n94585) );
  OAI21_X1 U80465 ( .B1(n107398), .B2(n105619), .A(n94587), .ZN(
        \DLX_Datapath/RegisterFile/N26588 ) );
  AOI22_X1 U80466 ( .A1(n105616), .A2(n110000), .B1(n94588), .B2(n105613), 
        .ZN(n94587) );
  OAI21_X1 U80467 ( .B1(n107400), .B2(n105618), .A(n94589), .ZN(
        \DLX_Datapath/RegisterFile/N26587 ) );
  AOI22_X1 U80468 ( .A1(n105616), .A2(n109883), .B1(n94590), .B2(n105614), 
        .ZN(n94589) );
  OAI21_X1 U80469 ( .B1(n107402), .B2(n105619), .A(n94591), .ZN(
        \DLX_Datapath/RegisterFile/N26586 ) );
  AOI22_X1 U80470 ( .A1(n105616), .A2(n108257), .B1(n94592), .B2(n105613), 
        .ZN(n94591) );
  OAI21_X1 U80471 ( .B1(n107404), .B2(n105618), .A(n94593), .ZN(
        \DLX_Datapath/RegisterFile/N26585 ) );
  AOI22_X1 U80472 ( .A1(n105616), .A2(n108380), .B1(n94594), .B2(n105614), 
        .ZN(n94593) );
  OAI21_X1 U80473 ( .B1(n107406), .B2(n105619), .A(n94595), .ZN(
        \DLX_Datapath/RegisterFile/N26584 ) );
  AOI22_X1 U80474 ( .A1(n105616), .A2(n108491), .B1(n94596), .B2(n105613), 
        .ZN(n94595) );
  OAI21_X1 U80475 ( .B1(n107408), .B2(n105618), .A(n94597), .ZN(
        \DLX_Datapath/RegisterFile/N26583 ) );
  AOI22_X1 U80476 ( .A1(n105616), .A2(n107728), .B1(n94598), .B2(n105614), 
        .ZN(n94597) );
  OAI21_X1 U80477 ( .B1(n107410), .B2(n105619), .A(n94599), .ZN(
        \DLX_Datapath/RegisterFile/N26582 ) );
  AOI22_X1 U80478 ( .A1(n105615), .A2(n109643), .B1(n94600), .B2(n105613), 
        .ZN(n94599) );
  OAI21_X1 U80479 ( .B1(n107412), .B2(n105619), .A(n94601), .ZN(
        \DLX_Datapath/RegisterFile/N26581 ) );
  AOI22_X1 U80480 ( .A1(n105615), .A2(n108605), .B1(n94602), .B2(n105612), 
        .ZN(n94601) );
  OAI21_X1 U80481 ( .B1(n107367), .B2(n105618), .A(n94603), .ZN(
        \DLX_Datapath/RegisterFile/N26580 ) );
  AOI22_X1 U80482 ( .A1(n105615), .A2(n109750), .B1(n94604), .B2(n105612), 
        .ZN(n94603) );
  OAI21_X1 U80483 ( .B1(n107369), .B2(n105619), .A(n94605), .ZN(
        \DLX_Datapath/RegisterFile/N26579 ) );
  AOI22_X1 U80484 ( .A1(n105615), .A2(n109535), .B1(n94606), .B2(n105612), 
        .ZN(n94605) );
  OAI21_X1 U80485 ( .B1(n108974), .B2(n105618), .A(n94607), .ZN(
        \DLX_Datapath/RegisterFile/N26578 ) );
  AOI22_X1 U80486 ( .A1(n105615), .A2(n109073), .B1(n94608), .B2(n105612), 
        .ZN(n94607) );
  OAI21_X1 U80487 ( .B1(n111063), .B2(n105618), .A(n94609), .ZN(
        \DLX_Datapath/RegisterFile/N26577 ) );
  AOI22_X1 U80488 ( .A1(n105615), .A2(n109420), .B1(n94610), .B2(n105612), 
        .ZN(n94609) );
  OAI21_X1 U80489 ( .B1(n111062), .B2(n105619), .A(n94611), .ZN(
        \DLX_Datapath/RegisterFile/N26576 ) );
  AOI22_X1 U80490 ( .A1(n105615), .A2(n109301), .B1(n94612), .B2(n105612), 
        .ZN(n94611) );
  OAI21_X1 U80491 ( .B1(n111061), .B2(n105618), .A(n94613), .ZN(
        \DLX_Datapath/RegisterFile/N26575 ) );
  AOI22_X1 U80492 ( .A1(n105615), .A2(n109193), .B1(n94614), .B2(n105612), 
        .ZN(n94613) );
  OAI21_X1 U80493 ( .B1(n111060), .B2(n105619), .A(n94615), .ZN(
        \DLX_Datapath/RegisterFile/N26574 ) );
  AOI22_X1 U80494 ( .A1(n105615), .A2(n108728), .B1(n94616), .B2(n105612), 
        .ZN(n94615) );
  OAI21_X1 U80495 ( .B1(n111059), .B2(n105618), .A(n94617), .ZN(
        \DLX_Datapath/RegisterFile/N26573 ) );
  AOI22_X1 U80496 ( .A1(n105615), .A2(n108956), .B1(n94618), .B2(n105612), 
        .ZN(n94617) );
  OAI21_X1 U80497 ( .B1(n111058), .B2(n105619), .A(n94619), .ZN(
        \DLX_Datapath/RegisterFile/N26572 ) );
  AOI22_X1 U80498 ( .A1(n105615), .A2(n108844), .B1(n94620), .B2(n105612), 
        .ZN(n94619) );
  OAI21_X1 U80499 ( .B1(n111057), .B2(n105618), .A(n94621), .ZN(
        \DLX_Datapath/RegisterFile/N26571 ) );
  AOI22_X1 U80500 ( .A1(n105615), .A2(n107179), .B1(n94622), .B2(n105612), 
        .ZN(n94621) );
  NAND2_X1 U80502 ( .A1(n94556), .A2(n111026), .ZN(n94623) );
  NOR2_X1 U80503 ( .A1(n94624), .A2(n105620), .ZN(n94558) );
  NAND2_X1 U80504 ( .A1(n105137), .A2(n94625), .ZN(n94556) );
  OAI21_X1 U80505 ( .B1(n107371), .B2(n105610), .A(n94627), .ZN(
        \DLX_Datapath/RegisterFile/N26570 ) );
  AOI22_X1 U80506 ( .A1(n105608), .A2(n107938), .B1(n105603), .B2(n81521), 
        .ZN(n94627) );
  OAI21_X1 U80507 ( .B1(n107373), .B2(n105610), .A(n94630), .ZN(
        \DLX_Datapath/RegisterFile/N26569 ) );
  AOI22_X1 U80508 ( .A1(n105608), .A2(n108034), .B1(n105604), .B2(n81653), 
        .ZN(n94630) );
  OAI21_X1 U80509 ( .B1(n106832), .B2(n105609), .A(n94631), .ZN(
        \DLX_Datapath/RegisterFile/N26568 ) );
  AOI22_X1 U80510 ( .A1(n105608), .A2(n107180), .B1(n105603), .B2(n81380), 
        .ZN(n94631) );
  OAI21_X1 U80511 ( .B1(n107376), .B2(n105609), .A(n94632), .ZN(
        \DLX_Datapath/RegisterFile/N26567 ) );
  AOI22_X1 U80512 ( .A1(n105608), .A2(n107843), .B1(n105604), .B2(n81377), 
        .ZN(n94632) );
  OAI21_X1 U80513 ( .B1(n107378), .B2(n105610), .A(n94633), .ZN(
        \DLX_Datapath/RegisterFile/N26566 ) );
  AOI22_X1 U80514 ( .A1(n105608), .A2(n110738), .B1(n105605), .B2(n81428), 
        .ZN(n94633) );
  OAI21_X1 U80515 ( .B1(n107380), .B2(n105610), .A(n94634), .ZN(
        \DLX_Datapath/RegisterFile/N26565 ) );
  AOI22_X1 U80516 ( .A1(n105608), .A2(n108143), .B1(n105605), .B2(n81410), 
        .ZN(n94634) );
  OAI21_X1 U80517 ( .B1(n107382), .B2(n105610), .A(n94635), .ZN(
        \DLX_Datapath/RegisterFile/N26564 ) );
  AOI22_X1 U80518 ( .A1(n105608), .A2(n110841), .B1(n105604), .B2(n81700), 
        .ZN(n94635) );
  OAI21_X1 U80519 ( .B1(n107384), .B2(n105610), .A(n94636), .ZN(
        \DLX_Datapath/RegisterFile/N26563 ) );
  AOI22_X1 U80520 ( .A1(n105608), .A2(n110942), .B1(n105603), .B2(n81632), 
        .ZN(n94636) );
  OAI21_X1 U80521 ( .B1(n107386), .B2(n105609), .A(n94637), .ZN(
        \DLX_Datapath/RegisterFile/N26562 ) );
  AOI22_X1 U80522 ( .A1(n105607), .A2(n110535), .B1(n105603), .B2(n81414), 
        .ZN(n94637) );
  OAI21_X1 U80523 ( .B1(n107388), .B2(n105609), .A(n94638), .ZN(
        \DLX_Datapath/RegisterFile/N26561 ) );
  AOI22_X1 U80524 ( .A1(n105607), .A2(n110320), .B1(n105605), .B2(n81317), 
        .ZN(n94638) );
  OAI21_X1 U80525 ( .B1(n107390), .B2(n105610), .A(n94639), .ZN(
        \DLX_Datapath/RegisterFile/N26560 ) );
  AOI22_X1 U80526 ( .A1(n105607), .A2(n110640), .B1(n105604), .B2(n81386), 
        .ZN(n94639) );
  OAI21_X1 U80527 ( .B1(n107392), .B2(n105609), .A(n94640), .ZN(
        \DLX_Datapath/RegisterFile/N26559 ) );
  AOI22_X1 U80528 ( .A1(n105607), .A2(n110429), .B1(n105603), .B2(n81320), 
        .ZN(n94640) );
  OAI21_X1 U80529 ( .B1(n107394), .B2(n105609), .A(n94641), .ZN(
        \DLX_Datapath/RegisterFile/N26558 ) );
  AOI22_X1 U80530 ( .A1(n105607), .A2(n110107), .B1(n105605), .B2(n81604), 
        .ZN(n94641) );
  OAI21_X1 U80531 ( .B1(n107396), .B2(n105609), .A(n94642), .ZN(
        \DLX_Datapath/RegisterFile/N26557 ) );
  AOI22_X1 U80532 ( .A1(n105607), .A2(n110214), .B1(n105604), .B2(n81405), 
        .ZN(n94642) );
  OAI21_X1 U80533 ( .B1(n107398), .B2(n105610), .A(n94643), .ZN(
        \DLX_Datapath/RegisterFile/N26556 ) );
  AOI22_X1 U80534 ( .A1(n105607), .A2(n109999), .B1(n105605), .B2(n81402), 
        .ZN(n94643) );
  OAI21_X1 U80535 ( .B1(n107400), .B2(n105610), .A(n94644), .ZN(
        \DLX_Datapath/RegisterFile/N26555 ) );
  AOI22_X1 U80536 ( .A1(n105607), .A2(n109882), .B1(n105603), .B2(n81400), 
        .ZN(n94644) );
  OAI21_X1 U80537 ( .B1(n107402), .B2(n105609), .A(n94645), .ZN(
        \DLX_Datapath/RegisterFile/N26554 ) );
  AOI22_X1 U80538 ( .A1(n105607), .A2(n108256), .B1(n105603), .B2(n81332), 
        .ZN(n94645) );
  OAI21_X1 U80539 ( .B1(n107404), .B2(n105609), .A(n94646), .ZN(
        \DLX_Datapath/RegisterFile/N26553 ) );
  AOI22_X1 U80540 ( .A1(n105607), .A2(n108379), .B1(n105604), .B2(n81373), 
        .ZN(n94646) );
  OAI21_X1 U80541 ( .B1(n107406), .B2(n105610), .A(n94647), .ZN(
        \DLX_Datapath/RegisterFile/N26552 ) );
  AOI22_X1 U80542 ( .A1(n105607), .A2(n108490), .B1(n105604), .B2(n81322), 
        .ZN(n94647) );
  OAI21_X1 U80543 ( .B1(n107408), .B2(n105609), .A(n94648), .ZN(
        \DLX_Datapath/RegisterFile/N26551 ) );
  AOI22_X1 U80544 ( .A1(n105607), .A2(n107727), .B1(n105605), .B2(n81506), 
        .ZN(n94648) );
  OAI21_X1 U80545 ( .B1(n107410), .B2(n105610), .A(n94649), .ZN(
        \DLX_Datapath/RegisterFile/N26550 ) );
  AOI22_X1 U80546 ( .A1(n105606), .A2(n109642), .B1(n105603), .B2(n81313), 
        .ZN(n94649) );
  OAI21_X1 U80547 ( .B1(n107412), .B2(n105609), .A(n94650), .ZN(
        \DLX_Datapath/RegisterFile/N26549 ) );
  AOI22_X1 U80548 ( .A1(n105606), .A2(n108604), .B1(n105604), .B2(n81330), 
        .ZN(n94650) );
  OAI21_X1 U80549 ( .B1(n107367), .B2(n105610), .A(n94651), .ZN(
        \DLX_Datapath/RegisterFile/N26548 ) );
  AOI22_X1 U80550 ( .A1(n105606), .A2(n109749), .B1(n105603), .B2(n81425), 
        .ZN(n94651) );
  OAI21_X1 U80551 ( .B1(n107369), .B2(n105609), .A(n94652), .ZN(
        \DLX_Datapath/RegisterFile/N26547 ) );
  AOI22_X1 U80552 ( .A1(n105606), .A2(n109534), .B1(n105605), .B2(n81396), 
        .ZN(n94652) );
  OAI21_X1 U80553 ( .B1(n108974), .B2(n105610), .A(n94653), .ZN(
        \DLX_Datapath/RegisterFile/N26546 ) );
  AOI22_X1 U80554 ( .A1(n105606), .A2(n109072), .B1(n105603), .B2(n81590), 
        .ZN(n94653) );
  OAI21_X1 U80555 ( .B1(n111063), .B2(n105609), .A(n94654), .ZN(
        \DLX_Datapath/RegisterFile/N26545 ) );
  AOI22_X1 U80556 ( .A1(n105606), .A2(n109419), .B1(n105604), .B2(n81423), 
        .ZN(n94654) );
  OAI21_X1 U80557 ( .B1(n111062), .B2(n105610), .A(n94655), .ZN(
        \DLX_Datapath/RegisterFile/N26544 ) );
  AOI22_X1 U80558 ( .A1(n105606), .A2(n109300), .B1(n105604), .B2(n81511), 
        .ZN(n94655) );
  OAI21_X1 U80559 ( .B1(n111061), .B2(n105610), .A(n94656), .ZN(
        \DLX_Datapath/RegisterFile/N26543 ) );
  AOI22_X1 U80560 ( .A1(n105606), .A2(n109192), .B1(n105605), .B2(n81503), 
        .ZN(n94656) );
  OAI21_X1 U80561 ( .B1(n111060), .B2(n105609), .A(n94657), .ZN(
        \DLX_Datapath/RegisterFile/N26542 ) );
  AOI22_X1 U80562 ( .A1(n105606), .A2(n108727), .B1(n105603), .B2(n81417), 
        .ZN(n94657) );
  OAI21_X1 U80563 ( .B1(n111059), .B2(n105610), .A(n94658), .ZN(
        \DLX_Datapath/RegisterFile/N26541 ) );
  AOI22_X1 U80564 ( .A1(n105606), .A2(n108955), .B1(n105605), .B2(n81500), 
        .ZN(n94658) );
  OAI21_X1 U80565 ( .B1(n111058), .B2(n105609), .A(n94659), .ZN(
        \DLX_Datapath/RegisterFile/N26540 ) );
  AOI22_X1 U80566 ( .A1(n105606), .A2(n108843), .B1(n105604), .B2(n81335), 
        .ZN(n94659) );
  OAI21_X1 U80567 ( .B1(n111057), .B2(n105609), .A(n94660), .ZN(
        \DLX_Datapath/RegisterFile/N26539 ) );
  AOI22_X1 U80568 ( .A1(n105606), .A2(n107181), .B1(n105605), .B2(n81327), 
        .ZN(n94660) );
  NAND2_X1 U80570 ( .A1(n94626), .A2(n111026), .ZN(n94661) );
  NOR2_X1 U80571 ( .A1(n105611), .A2(n94624), .ZN(n94628) );
  AOI21_X1 U80572 ( .B1(n105206), .B2(n94662), .A(n94663), .ZN(n94624) );
  OR2_X1 U80573 ( .A1(n86230), .A2(n94553), .ZN(n94662) );
  NAND2_X1 U80574 ( .A1(n105137), .A2(n94664), .ZN(n94626) );
  OAI21_X1 U80575 ( .B1(n107371), .B2(n105600), .A(n94666), .ZN(
        \DLX_Datapath/RegisterFile/N26538 ) );
  AOI22_X1 U80576 ( .A1(n94667), .A2(n105002), .B1(n105187), .B2(n107937), 
        .ZN(n94666) );
  OAI21_X1 U80577 ( .B1(n107373), .B2(n105600), .A(n94669), .ZN(
        \DLX_Datapath/RegisterFile/N26537 ) );
  AOI22_X1 U80578 ( .A1(n94670), .A2(n105003), .B1(n105186), .B2(n108033), 
        .ZN(n94669) );
  OAI21_X1 U80579 ( .B1(n106832), .B2(n105600), .A(n94671), .ZN(
        \DLX_Datapath/RegisterFile/N26536 ) );
  AOI22_X1 U80580 ( .A1(n94672), .A2(n105003), .B1(n105187), .B2(n107182), 
        .ZN(n94671) );
  OAI21_X1 U80581 ( .B1(n107376), .B2(n105600), .A(n94673), .ZN(
        \DLX_Datapath/RegisterFile/N26535 ) );
  AOI22_X1 U80582 ( .A1(n94674), .A2(n105002), .B1(n105187), .B2(n107842), 
        .ZN(n94673) );
  OAI21_X1 U80583 ( .B1(n107378), .B2(n105600), .A(n94675), .ZN(
        \DLX_Datapath/RegisterFile/N26534 ) );
  AOI22_X1 U80584 ( .A1(n94676), .A2(n105003), .B1(n105186), .B2(n110737), 
        .ZN(n94675) );
  OAI21_X1 U80585 ( .B1(n107380), .B2(n105600), .A(n94677), .ZN(
        \DLX_Datapath/RegisterFile/N26533 ) );
  AOI22_X1 U80586 ( .A1(n94678), .A2(n105002), .B1(n105186), .B2(n108142), 
        .ZN(n94677) );
  OAI21_X1 U80587 ( .B1(n107382), .B2(n105600), .A(n94679), .ZN(
        \DLX_Datapath/RegisterFile/N26532 ) );
  AOI22_X1 U80588 ( .A1(n94680), .A2(n105002), .B1(n105187), .B2(n110840), 
        .ZN(n94679) );
  OAI21_X1 U80589 ( .B1(n107384), .B2(n105600), .A(n94681), .ZN(
        \DLX_Datapath/RegisterFile/N26531 ) );
  AOI22_X1 U80590 ( .A1(n94682), .A2(n105002), .B1(n105186), .B2(n110941), 
        .ZN(n94681) );
  OAI21_X1 U80591 ( .B1(n107386), .B2(n105600), .A(n94683), .ZN(
        \DLX_Datapath/RegisterFile/N26530 ) );
  AOI22_X1 U80592 ( .A1(n94684), .A2(n105003), .B1(n105186), .B2(n110534), 
        .ZN(n94683) );
  OAI21_X1 U80593 ( .B1(n107388), .B2(n105600), .A(n94685), .ZN(
        \DLX_Datapath/RegisterFile/N26529 ) );
  AOI22_X1 U80594 ( .A1(n94686), .A2(n105003), .B1(n105187), .B2(n110319), 
        .ZN(n94685) );
  OAI21_X1 U80595 ( .B1(n107390), .B2(n105600), .A(n94687), .ZN(
        \DLX_Datapath/RegisterFile/N26528 ) );
  AOI22_X1 U80596 ( .A1(n94688), .A2(n105003), .B1(n106756), .B2(n110639), 
        .ZN(n94687) );
  OAI21_X1 U80597 ( .B1(n107392), .B2(n105600), .A(n94689), .ZN(
        \DLX_Datapath/RegisterFile/N26527 ) );
  AOI22_X1 U80598 ( .A1(n94690), .A2(n105003), .B1(n106756), .B2(n110428), 
        .ZN(n94689) );
  OAI21_X1 U80599 ( .B1(n107394), .B2(n105600), .A(n94691), .ZN(
        \DLX_Datapath/RegisterFile/N26526 ) );
  AOI22_X1 U80600 ( .A1(n94692), .A2(n105002), .B1(n106756), .B2(n110106), 
        .ZN(n94691) );
  OAI21_X1 U80601 ( .B1(n107396), .B2(n105600), .A(n94693), .ZN(
        \DLX_Datapath/RegisterFile/N26525 ) );
  AOI22_X1 U80602 ( .A1(n94694), .A2(n105003), .B1(n106756), .B2(n110213), 
        .ZN(n94693) );
  OAI21_X1 U80603 ( .B1(n107398), .B2(n105600), .A(n94695), .ZN(
        \DLX_Datapath/RegisterFile/N26524 ) );
  AOI22_X1 U80604 ( .A1(n94696), .A2(n105002), .B1(n105186), .B2(n109998), 
        .ZN(n94695) );
  OAI21_X1 U80605 ( .B1(n107400), .B2(n105600), .A(n94697), .ZN(
        \DLX_Datapath/RegisterFile/N26523 ) );
  AOI22_X1 U80606 ( .A1(n94698), .A2(n105002), .B1(n106756), .B2(n109881), 
        .ZN(n94697) );
  OAI21_X1 U80607 ( .B1(n107402), .B2(n105600), .A(n94699), .ZN(
        \DLX_Datapath/RegisterFile/N26522 ) );
  AOI22_X1 U80608 ( .A1(n94700), .A2(n105003), .B1(n106756), .B2(n108255), 
        .ZN(n94699) );
  OAI21_X1 U80609 ( .B1(n107404), .B2(n105600), .A(n94701), .ZN(
        \DLX_Datapath/RegisterFile/N26521 ) );
  AOI22_X1 U80610 ( .A1(n94702), .A2(n105003), .B1(n105187), .B2(n108378), 
        .ZN(n94701) );
  OAI21_X1 U80611 ( .B1(n107406), .B2(n105600), .A(n94703), .ZN(
        \DLX_Datapath/RegisterFile/N26520 ) );
  AOI22_X1 U80612 ( .A1(n94704), .A2(n94668), .B1(n106756), .B2(n108489), .ZN(
        n94703) );
  OAI21_X1 U80613 ( .B1(n107408), .B2(n105600), .A(n94705), .ZN(
        \DLX_Datapath/RegisterFile/N26519 ) );
  AOI22_X1 U80614 ( .A1(n94706), .A2(n105003), .B1(n105187), .B2(n107726), 
        .ZN(n94705) );
  OAI21_X1 U80615 ( .B1(n107410), .B2(n105600), .A(n94707), .ZN(
        \DLX_Datapath/RegisterFile/N26518 ) );
  AOI22_X1 U80616 ( .A1(n94708), .A2(n105002), .B1(n106756), .B2(n109641), 
        .ZN(n94707) );
  OAI21_X1 U80617 ( .B1(n107412), .B2(n105600), .A(n94709), .ZN(
        \DLX_Datapath/RegisterFile/N26517 ) );
  AOI22_X1 U80618 ( .A1(n94710), .A2(n105002), .B1(n105187), .B2(n108603), 
        .ZN(n94709) );
  OAI21_X1 U80619 ( .B1(n107367), .B2(n105600), .A(n94711), .ZN(
        \DLX_Datapath/RegisterFile/N26516 ) );
  AOI22_X1 U80620 ( .A1(n94712), .A2(n105002), .B1(n105186), .B2(n109748), 
        .ZN(n94711) );
  OAI21_X1 U80621 ( .B1(n107369), .B2(n105600), .A(n94713), .ZN(
        \DLX_Datapath/RegisterFile/N26515 ) );
  AOI22_X1 U80622 ( .A1(n94714), .A2(n105003), .B1(n105186), .B2(n109533), 
        .ZN(n94713) );
  OAI21_X1 U80623 ( .B1(n108974), .B2(n105600), .A(n94715), .ZN(
        \DLX_Datapath/RegisterFile/N26514 ) );
  AOI22_X1 U80624 ( .A1(n105002), .A2(n81259), .B1(n105187), .B2(n109071), 
        .ZN(n94715) );
  OAI21_X1 U80625 ( .B1(n111063), .B2(n105600), .A(n94716), .ZN(
        \DLX_Datapath/RegisterFile/N26513 ) );
  AOI22_X1 U80626 ( .A1(n94717), .A2(n94668), .B1(n105187), .B2(n109418), .ZN(
        n94716) );
  OAI21_X1 U80627 ( .B1(n111062), .B2(n105600), .A(n94718), .ZN(
        \DLX_Datapath/RegisterFile/N26512 ) );
  AOI22_X1 U80628 ( .A1(n94719), .A2(n105002), .B1(n105186), .B2(n109299), 
        .ZN(n94718) );
  OAI21_X1 U80629 ( .B1(n111061), .B2(n105600), .A(n94720), .ZN(
        \DLX_Datapath/RegisterFile/N26511 ) );
  AOI22_X1 U80630 ( .A1(n94721), .A2(n105002), .B1(n105186), .B2(n109191), 
        .ZN(n94720) );
  OAI21_X1 U80631 ( .B1(n111060), .B2(n105600), .A(n94722), .ZN(
        \DLX_Datapath/RegisterFile/N26510 ) );
  AOI22_X1 U80632 ( .A1(n94723), .A2(n105003), .B1(n105187), .B2(n108726), 
        .ZN(n94722) );
  OAI21_X1 U80633 ( .B1(n111059), .B2(n105600), .A(n94724), .ZN(
        \DLX_Datapath/RegisterFile/N26509 ) );
  AOI22_X1 U80634 ( .A1(n94725), .A2(n94668), .B1(n105186), .B2(n108954), .ZN(
        n94724) );
  OAI21_X1 U80635 ( .B1(n111058), .B2(n105600), .A(n94726), .ZN(
        \DLX_Datapath/RegisterFile/N26508 ) );
  AOI22_X1 U80636 ( .A1(n94727), .A2(n94668), .B1(n105187), .B2(n108842), .ZN(
        n94726) );
  OAI21_X1 U80637 ( .B1(n111057), .B2(n105600), .A(n94728), .ZN(
        \DLX_Datapath/RegisterFile/N26507 ) );
  AOI22_X1 U80638 ( .A1(n94729), .A2(n105003), .B1(n105186), .B2(n107183), 
        .ZN(n94728) );
  OAI21_X1 U80639 ( .B1(n94731), .B2(n94663), .A(n94665), .ZN(n94730) );
  AOI21_X1 U80640 ( .B1(n94732), .B2(n111026), .A(n94366), .ZN(n94731) );
  NOR2_X1 U80641 ( .A1(n94733), .A2(n106754), .ZN(n94668) );
  NAND2_X1 U80642 ( .A1(n94665), .A2(n111026), .ZN(n94733) );
  NAND2_X1 U80643 ( .A1(n105137), .A2(n94734), .ZN(n94665) );
  OAI21_X1 U80644 ( .B1(n107371), .B2(n105598), .A(n94736), .ZN(
        \DLX_Datapath/RegisterFile/N26506 ) );
  AOI22_X1 U80645 ( .A1(n105597), .A2(n107936), .B1(n105594), .B2(n81360), 
        .ZN(n94736) );
  OAI21_X1 U80646 ( .B1(n107373), .B2(n105598), .A(n94739), .ZN(
        \DLX_Datapath/RegisterFile/N26505 ) );
  AOI22_X1 U80647 ( .A1(n105597), .A2(n108032), .B1(n105593), .B2(n94511), 
        .ZN(n94739) );
  OAI21_X1 U80648 ( .B1(n106832), .B2(n105599), .A(n94740), .ZN(
        \DLX_Datapath/RegisterFile/N26504 ) );
  AOI22_X1 U80649 ( .A1(n105597), .A2(n107184), .B1(n105593), .B2(n81539), 
        .ZN(n94740) );
  OAI21_X1 U80650 ( .B1(n107376), .B2(n105598), .A(n94741), .ZN(
        \DLX_Datapath/RegisterFile/N26503 ) );
  AOI22_X1 U80651 ( .A1(n105597), .A2(n107841), .B1(n105593), .B2(n81301), 
        .ZN(n94741) );
  OAI21_X1 U80652 ( .B1(n107378), .B2(n105598), .A(n94742), .ZN(
        \DLX_Datapath/RegisterFile/N26502 ) );
  AOI22_X1 U80653 ( .A1(n105597), .A2(n110736), .B1(n105594), .B2(n81308), 
        .ZN(n94742) );
  OAI21_X1 U80654 ( .B1(n107380), .B2(n105598), .A(n94743), .ZN(
        \DLX_Datapath/RegisterFile/N26501 ) );
  AOI22_X1 U80655 ( .A1(n105597), .A2(n108141), .B1(n105594), .B2(n94516), 
        .ZN(n94743) );
  OAI21_X1 U80656 ( .B1(n107382), .B2(n105599), .A(n94744), .ZN(
        \DLX_Datapath/RegisterFile/N26500 ) );
  AOI22_X1 U80657 ( .A1(n105597), .A2(n110839), .B1(n105594), .B2(n81272), 
        .ZN(n94744) );
  OAI21_X1 U80658 ( .B1(n107384), .B2(n105599), .A(n94745), .ZN(
        \DLX_Datapath/RegisterFile/N26499 ) );
  AOI22_X1 U80659 ( .A1(n105597), .A2(n110940), .B1(n105593), .B2(n94519), 
        .ZN(n94745) );
  OAI21_X1 U80660 ( .B1(n107386), .B2(n105598), .A(n94746), .ZN(
        \DLX_Datapath/RegisterFile/N26498 ) );
  AOI22_X1 U80661 ( .A1(n105596), .A2(n110533), .B1(n105593), .B2(n80192), 
        .ZN(n94746) );
  OAI21_X1 U80662 ( .B1(n107388), .B2(n105599), .A(n94747), .ZN(
        \DLX_Datapath/RegisterFile/N26497 ) );
  AOI22_X1 U80663 ( .A1(n105596), .A2(n110318), .B1(n105594), .B2(n81474), 
        .ZN(n94747) );
  OAI21_X1 U80664 ( .B1(n107390), .B2(n105599), .A(n94748), .ZN(
        \DLX_Datapath/RegisterFile/N26496 ) );
  AOI22_X1 U80665 ( .A1(n105596), .A2(n110638), .B1(n105593), .B2(n94523), 
        .ZN(n94748) );
  OAI21_X1 U80666 ( .B1(n107392), .B2(n105598), .A(n94749), .ZN(
        \DLX_Datapath/RegisterFile/N26495 ) );
  AOI22_X1 U80667 ( .A1(n105596), .A2(n110427), .B1(n105594), .B2(n106061), 
        .ZN(n94749) );
  OAI21_X1 U80668 ( .B1(n107394), .B2(n105599), .A(n94750), .ZN(
        \DLX_Datapath/RegisterFile/N26494 ) );
  AOI22_X1 U80669 ( .A1(n105596), .A2(n110105), .B1(n105593), .B2(n81347), 
        .ZN(n94750) );
  OAI21_X1 U80670 ( .B1(n107396), .B2(n105599), .A(n94751), .ZN(
        \DLX_Datapath/RegisterFile/N26493 ) );
  AOI22_X1 U80671 ( .A1(n105596), .A2(n110212), .B1(n105594), .B2(n94527), 
        .ZN(n94751) );
  OAI21_X1 U80672 ( .B1(n107398), .B2(n105598), .A(n94752), .ZN(
        \DLX_Datapath/RegisterFile/N26492 ) );
  AOI22_X1 U80673 ( .A1(n105596), .A2(n109997), .B1(n105593), .B2(n81297), 
        .ZN(n94752) );
  OAI21_X1 U80674 ( .B1(n107400), .B2(n105599), .A(n94753), .ZN(
        \DLX_Datapath/RegisterFile/N26491 ) );
  AOI22_X1 U80675 ( .A1(n105596), .A2(n109880), .B1(n105594), .B2(n94530), 
        .ZN(n94753) );
  OAI21_X1 U80676 ( .B1(n107402), .B2(n105598), .A(n94754), .ZN(
        \DLX_Datapath/RegisterFile/N26490 ) );
  AOI22_X1 U80677 ( .A1(n105596), .A2(n108254), .B1(n105593), .B2(n81286), 
        .ZN(n94754) );
  OAI21_X1 U80678 ( .B1(n107404), .B2(n105598), .A(n94755), .ZN(
        \DLX_Datapath/RegisterFile/N26489 ) );
  AOI22_X1 U80679 ( .A1(n105596), .A2(n108377), .B1(n105594), .B2(n106169), 
        .ZN(n94755) );
  OAI21_X1 U80680 ( .B1(n107406), .B2(n105599), .A(n94756), .ZN(
        \DLX_Datapath/RegisterFile/N26488 ) );
  AOI22_X1 U80681 ( .A1(n105596), .A2(n108488), .B1(n105593), .B2(n81283), 
        .ZN(n94756) );
  OAI21_X1 U80682 ( .B1(n107408), .B2(n105599), .A(n94757), .ZN(
        \DLX_Datapath/RegisterFile/N26487 ) );
  AOI22_X1 U80683 ( .A1(n105596), .A2(n107725), .B1(n105594), .B2(n81453), 
        .ZN(n94757) );
  OAI21_X1 U80684 ( .B1(n107410), .B2(n105599), .A(n94758), .ZN(
        \DLX_Datapath/RegisterFile/N26486 ) );
  AOI22_X1 U80685 ( .A1(n105595), .A2(n109640), .B1(n105593), .B2(n94536), 
        .ZN(n94758) );
  OAI21_X1 U80686 ( .B1(n107412), .B2(n105599), .A(n94759), .ZN(
        \DLX_Datapath/RegisterFile/N26485 ) );
  AOI22_X1 U80687 ( .A1(n105595), .A2(n108602), .B1(n105592), .B2(n106241), 
        .ZN(n94759) );
  OAI21_X1 U80688 ( .B1(n107367), .B2(n105599), .A(n94760), .ZN(
        \DLX_Datapath/RegisterFile/N26484 ) );
  AOI22_X1 U80689 ( .A1(n105595), .A2(n109747), .B1(n105592), .B2(n81351), 
        .ZN(n94760) );
  OAI21_X1 U80690 ( .B1(n107369), .B2(n105598), .A(n94761), .ZN(
        \DLX_Datapath/RegisterFile/N26483 ) );
  AOI22_X1 U80691 ( .A1(n105595), .A2(n109532), .B1(n105592), .B2(n106020), 
        .ZN(n94761) );
  OAI21_X1 U80692 ( .B1(n108974), .B2(n105599), .A(n94762), .ZN(
        \DLX_Datapath/RegisterFile/N26482 ) );
  AOI22_X1 U80693 ( .A1(n105595), .A2(n109070), .B1(n105592), .B2(n94541), 
        .ZN(n94762) );
  OAI21_X1 U80694 ( .B1(n111063), .B2(n105598), .A(n94763), .ZN(
        \DLX_Datapath/RegisterFile/N26481 ) );
  AOI22_X1 U80695 ( .A1(n105595), .A2(n109417), .B1(n105592), .B2(n81269), 
        .ZN(n94763) );
  OAI21_X1 U80696 ( .B1(n111062), .B2(n105599), .A(n94764), .ZN(
        \DLX_Datapath/RegisterFile/N26480 ) );
  AOI22_X1 U80697 ( .A1(n105595), .A2(n109298), .B1(n105592), .B2(n105624), 
        .ZN(n94764) );
  OAI21_X1 U80698 ( .B1(n111061), .B2(n105598), .A(n94765), .ZN(
        \DLX_Datapath/RegisterFile/N26479 ) );
  AOI22_X1 U80699 ( .A1(n105595), .A2(n109190), .B1(n105592), .B2(n94546), 
        .ZN(n94765) );
  OAI21_X1 U80700 ( .B1(n111060), .B2(n105598), .A(n94766), .ZN(
        \DLX_Datapath/RegisterFile/N26478 ) );
  AOI22_X1 U80701 ( .A1(n105595), .A2(n108725), .B1(n105592), .B2(n94548), 
        .ZN(n94766) );
  OAI21_X1 U80702 ( .B1(n111059), .B2(n105598), .A(n94767), .ZN(
        \DLX_Datapath/RegisterFile/N26477 ) );
  AOI22_X1 U80703 ( .A1(n105595), .A2(n108953), .B1(n105592), .B2(n81783), 
        .ZN(n94767) );
  OAI21_X1 U80704 ( .B1(n111058), .B2(n105598), .A(n94768), .ZN(
        \DLX_Datapath/RegisterFile/N26476 ) );
  AOI22_X1 U80705 ( .A1(n105595), .A2(n108841), .B1(n105592), .B2(n80188), 
        .ZN(n94768) );
  OAI21_X1 U80706 ( .B1(n111057), .B2(n105599), .A(n94769), .ZN(
        \DLX_Datapath/RegisterFile/N26475 ) );
  AOI22_X1 U80707 ( .A1(n105595), .A2(n107185), .B1(n105592), .B2(n81265), 
        .ZN(n94769) );
  NAND2_X1 U80709 ( .A1(n94735), .A2(n111024), .ZN(n94770) );
  AOI21_X1 U80710 ( .B1(n94259), .B2(n94771), .A(n105011), .ZN(n94737) );
  NAND2_X1 U80711 ( .A1(n94553), .A2(n105205), .ZN(n94259) );
  NAND2_X1 U80712 ( .A1(n105137), .A2(n94772), .ZN(n94735) );
  OAI21_X1 U80713 ( .B1(n107371), .B2(n105590), .A(n94774), .ZN(
        \DLX_Datapath/RegisterFile/N26474 ) );
  AOI22_X1 U80714 ( .A1(n105589), .A2(n107935), .B1(n94776), .B2(n94559), .ZN(
        n94774) );
  OAI21_X1 U80715 ( .B1(n107373), .B2(n105590), .A(n94777), .ZN(
        \DLX_Datapath/RegisterFile/N26473 ) );
  AOI22_X1 U80716 ( .A1(n105589), .A2(n108031), .B1(n104813), .B2(n94562), 
        .ZN(n94777) );
  OAI21_X1 U80717 ( .B1(n106832), .B2(n105590), .A(n94778), .ZN(
        \DLX_Datapath/RegisterFile/N26472 ) );
  AOI22_X1 U80718 ( .A1(n105589), .A2(n107186), .B1(n104813), .B2(n94564), 
        .ZN(n94778) );
  OAI21_X1 U80719 ( .B1(n107376), .B2(n105590), .A(n94779), .ZN(
        \DLX_Datapath/RegisterFile/N26471 ) );
  AOI22_X1 U80720 ( .A1(n105589), .A2(n107840), .B1(n104812), .B2(n94566), 
        .ZN(n94779) );
  OAI21_X1 U80721 ( .B1(n107378), .B2(n105590), .A(n94780), .ZN(
        \DLX_Datapath/RegisterFile/N26470 ) );
  AOI22_X1 U80722 ( .A1(n105589), .A2(n110735), .B1(n104813), .B2(n94568), 
        .ZN(n94780) );
  OAI21_X1 U80723 ( .B1(n107380), .B2(n105590), .A(n94781), .ZN(
        \DLX_Datapath/RegisterFile/N26469 ) );
  AOI22_X1 U80724 ( .A1(n105589), .A2(n108140), .B1(n104812), .B2(n94570), 
        .ZN(n94781) );
  OAI21_X1 U80725 ( .B1(n107382), .B2(n105590), .A(n94782), .ZN(
        \DLX_Datapath/RegisterFile/N26468 ) );
  AOI22_X1 U80726 ( .A1(n105589), .A2(n110838), .B1(n104813), .B2(n94572), 
        .ZN(n94782) );
  OAI21_X1 U80727 ( .B1(n107384), .B2(n105590), .A(n94783), .ZN(
        \DLX_Datapath/RegisterFile/N26467 ) );
  AOI22_X1 U80728 ( .A1(n105589), .A2(n110939), .B1(n104813), .B2(n94574), 
        .ZN(n94783) );
  OAI21_X1 U80729 ( .B1(n107386), .B2(n105590), .A(n94784), .ZN(
        \DLX_Datapath/RegisterFile/N26466 ) );
  AOI22_X1 U80730 ( .A1(n105588), .A2(n110532), .B1(n104812), .B2(n94576), 
        .ZN(n94784) );
  OAI21_X1 U80731 ( .B1(n107388), .B2(n105590), .A(n94785), .ZN(
        \DLX_Datapath/RegisterFile/N26465 ) );
  AOI22_X1 U80732 ( .A1(n105588), .A2(n110317), .B1(n104813), .B2(n94578), 
        .ZN(n94785) );
  OAI21_X1 U80733 ( .B1(n107390), .B2(n105590), .A(n94786), .ZN(
        \DLX_Datapath/RegisterFile/N26464 ) );
  AOI22_X1 U80734 ( .A1(n105588), .A2(n110637), .B1(n104812), .B2(n94580), 
        .ZN(n94786) );
  OAI21_X1 U80735 ( .B1(n107392), .B2(n105590), .A(n94787), .ZN(
        \DLX_Datapath/RegisterFile/N26463 ) );
  AOI22_X1 U80736 ( .A1(n105588), .A2(n110426), .B1(n94776), .B2(n94582), .ZN(
        n94787) );
  OAI21_X1 U80737 ( .B1(n107394), .B2(n105590), .A(n94788), .ZN(
        \DLX_Datapath/RegisterFile/N26462 ) );
  AOI22_X1 U80738 ( .A1(n105588), .A2(n110104), .B1(n104812), .B2(n94584), 
        .ZN(n94788) );
  OAI21_X1 U80739 ( .B1(n107396), .B2(n105590), .A(n94789), .ZN(
        \DLX_Datapath/RegisterFile/N26461 ) );
  AOI22_X1 U80740 ( .A1(n105588), .A2(n110211), .B1(n104813), .B2(n94586), 
        .ZN(n94789) );
  OAI21_X1 U80741 ( .B1(n107398), .B2(n105590), .A(n94790), .ZN(
        \DLX_Datapath/RegisterFile/N26460 ) );
  AOI22_X1 U80742 ( .A1(n105588), .A2(n109996), .B1(n104813), .B2(n94588), 
        .ZN(n94790) );
  OAI21_X1 U80743 ( .B1(n107400), .B2(n105590), .A(n94791), .ZN(
        \DLX_Datapath/RegisterFile/N26459 ) );
  AOI22_X1 U80744 ( .A1(n105588), .A2(n109879), .B1(n104813), .B2(n94590), 
        .ZN(n94791) );
  OAI21_X1 U80745 ( .B1(n107402), .B2(n105590), .A(n94792), .ZN(
        \DLX_Datapath/RegisterFile/N26458 ) );
  AOI22_X1 U80746 ( .A1(n105588), .A2(n108253), .B1(n104812), .B2(n94592), 
        .ZN(n94792) );
  OAI21_X1 U80747 ( .B1(n107404), .B2(n105590), .A(n94793), .ZN(
        \DLX_Datapath/RegisterFile/N26457 ) );
  AOI22_X1 U80748 ( .A1(n105588), .A2(n108376), .B1(n94776), .B2(n94594), .ZN(
        n94793) );
  OAI21_X1 U80749 ( .B1(n107406), .B2(n105590), .A(n94794), .ZN(
        \DLX_Datapath/RegisterFile/N26456 ) );
  AOI22_X1 U80750 ( .A1(n105588), .A2(n108487), .B1(n94776), .B2(n94596), .ZN(
        n94794) );
  OAI21_X1 U80751 ( .B1(n107408), .B2(n105590), .A(n94795), .ZN(
        \DLX_Datapath/RegisterFile/N26455 ) );
  AOI22_X1 U80752 ( .A1(n105588), .A2(n107724), .B1(n104813), .B2(n94598), 
        .ZN(n94795) );
  OAI21_X1 U80753 ( .B1(n107410), .B2(n105590), .A(n94796), .ZN(
        \DLX_Datapath/RegisterFile/N26454 ) );
  AOI22_X1 U80754 ( .A1(n105587), .A2(n109639), .B1(n94776), .B2(n94600), .ZN(
        n94796) );
  OAI21_X1 U80755 ( .B1(n107412), .B2(n105590), .A(n94797), .ZN(
        \DLX_Datapath/RegisterFile/N26453 ) );
  AOI22_X1 U80756 ( .A1(n105587), .A2(n108601), .B1(n94776), .B2(n94602), .ZN(
        n94797) );
  OAI21_X1 U80757 ( .B1(n107367), .B2(n105590), .A(n94798), .ZN(
        \DLX_Datapath/RegisterFile/N26452 ) );
  AOI22_X1 U80758 ( .A1(n105587), .A2(n109746), .B1(n94776), .B2(n94604), .ZN(
        n94798) );
  OAI21_X1 U80759 ( .B1(n107369), .B2(n105590), .A(n94799), .ZN(
        \DLX_Datapath/RegisterFile/N26451 ) );
  AOI22_X1 U80760 ( .A1(n105587), .A2(n109531), .B1(n94776), .B2(n94606), .ZN(
        n94799) );
  OAI21_X1 U80761 ( .B1(n108974), .B2(n105590), .A(n94800), .ZN(
        \DLX_Datapath/RegisterFile/N26450 ) );
  AOI22_X1 U80762 ( .A1(n105587), .A2(n109069), .B1(n94776), .B2(n94608), .ZN(
        n94800) );
  OAI21_X1 U80763 ( .B1(n111063), .B2(n105590), .A(n94801), .ZN(
        \DLX_Datapath/RegisterFile/N26449 ) );
  AOI22_X1 U80764 ( .A1(n105587), .A2(n109416), .B1(n94776), .B2(n94610), .ZN(
        n94801) );
  OAI21_X1 U80765 ( .B1(n111062), .B2(n105590), .A(n94802), .ZN(
        \DLX_Datapath/RegisterFile/N26448 ) );
  AOI22_X1 U80766 ( .A1(n105587), .A2(n109297), .B1(n104813), .B2(n94612), 
        .ZN(n94802) );
  OAI21_X1 U80767 ( .B1(n111061), .B2(n105590), .A(n94803), .ZN(
        \DLX_Datapath/RegisterFile/N26447 ) );
  AOI22_X1 U80768 ( .A1(n105587), .A2(n109189), .B1(n104812), .B2(n94614), 
        .ZN(n94803) );
  OAI21_X1 U80769 ( .B1(n111060), .B2(n105590), .A(n94804), .ZN(
        \DLX_Datapath/RegisterFile/N26446 ) );
  AOI22_X1 U80770 ( .A1(n105587), .A2(n108724), .B1(n94776), .B2(n94616), .ZN(
        n94804) );
  OAI21_X1 U80771 ( .B1(n111059), .B2(n105590), .A(n94805), .ZN(
        \DLX_Datapath/RegisterFile/N26445 ) );
  AOI22_X1 U80772 ( .A1(n105587), .A2(n108952), .B1(n104812), .B2(n94618), 
        .ZN(n94805) );
  OAI21_X1 U80773 ( .B1(n111058), .B2(n105590), .A(n94806), .ZN(
        \DLX_Datapath/RegisterFile/N26444 ) );
  AOI22_X1 U80774 ( .A1(n105587), .A2(n108840), .B1(n104812), .B2(n94620), 
        .ZN(n94806) );
  OAI21_X1 U80775 ( .B1(n111057), .B2(n105590), .A(n94807), .ZN(
        \DLX_Datapath/RegisterFile/N26443 ) );
  AOI22_X1 U80776 ( .A1(n105587), .A2(n107187), .B1(n104812), .B2(n94622), 
        .ZN(n94807) );
  NOR2_X1 U80777 ( .A1(n94808), .A2(n94553), .ZN(n94776) );
  NAND2_X1 U80778 ( .A1(n94773), .A2(n111024), .ZN(n94808) );
  NOR2_X1 U80779 ( .A1(n94809), .A2(n105591), .ZN(n94775) );
  NAND2_X1 U80780 ( .A1(n105136), .A2(n94810), .ZN(n94773) );
  OAI21_X1 U80781 ( .B1(n107371), .B2(n105585), .A(n94812), .ZN(
        \DLX_Datapath/RegisterFile/N26442 ) );
  AOI22_X1 U80782 ( .A1(n105584), .A2(n107934), .B1(n105581), .B2(n81521), 
        .ZN(n94812) );
  OAI21_X1 U80783 ( .B1(n107373), .B2(n105585), .A(n94815), .ZN(
        \DLX_Datapath/RegisterFile/N26441 ) );
  AOI22_X1 U80784 ( .A1(n105584), .A2(n108030), .B1(n105580), .B2(n81653), 
        .ZN(n94815) );
  OAI21_X1 U80785 ( .B1(n106832), .B2(n105585), .A(n94816), .ZN(
        \DLX_Datapath/RegisterFile/N26440 ) );
  AOI22_X1 U80786 ( .A1(n105584), .A2(n107188), .B1(n105581), .B2(n81380), 
        .ZN(n94816) );
  OAI21_X1 U80787 ( .B1(n107376), .B2(n105585), .A(n94817), .ZN(
        \DLX_Datapath/RegisterFile/N26439 ) );
  AOI22_X1 U80788 ( .A1(n105584), .A2(n107839), .B1(n105580), .B2(n81377), 
        .ZN(n94817) );
  OAI21_X1 U80789 ( .B1(n107378), .B2(n105585), .A(n94818), .ZN(
        \DLX_Datapath/RegisterFile/N26438 ) );
  AOI22_X1 U80790 ( .A1(n105584), .A2(n110734), .B1(n105581), .B2(n81428), 
        .ZN(n94818) );
  OAI21_X1 U80791 ( .B1(n107380), .B2(n105585), .A(n94819), .ZN(
        \DLX_Datapath/RegisterFile/N26437 ) );
  AOI22_X1 U80792 ( .A1(n105584), .A2(n108139), .B1(n105580), .B2(n81410), 
        .ZN(n94819) );
  OAI21_X1 U80793 ( .B1(n107382), .B2(n105585), .A(n94820), .ZN(
        \DLX_Datapath/RegisterFile/N26436 ) );
  AOI22_X1 U80794 ( .A1(n105584), .A2(n110837), .B1(n105580), .B2(n81700), 
        .ZN(n94820) );
  OAI21_X1 U80795 ( .B1(n107384), .B2(n105585), .A(n94821), .ZN(
        \DLX_Datapath/RegisterFile/N26435 ) );
  AOI22_X1 U80796 ( .A1(n105584), .A2(n110938), .B1(n105581), .B2(n81632), 
        .ZN(n94821) );
  OAI21_X1 U80797 ( .B1(n107386), .B2(n105585), .A(n94822), .ZN(
        \DLX_Datapath/RegisterFile/N26434 ) );
  AOI22_X1 U80798 ( .A1(n105583), .A2(n110531), .B1(n105580), .B2(n81414), 
        .ZN(n94822) );
  OAI21_X1 U80799 ( .B1(n107388), .B2(n105585), .A(n94823), .ZN(
        \DLX_Datapath/RegisterFile/N26433 ) );
  AOI22_X1 U80800 ( .A1(n105583), .A2(n110316), .B1(n105581), .B2(n81317), 
        .ZN(n94823) );
  AOI22_X1 U80802 ( .A1(n105583), .A2(n110636), .B1(n105580), .B2(n81386), 
        .ZN(n94824) );
  OAI21_X1 U80803 ( .B1(n107392), .B2(n105586), .A(n94825), .ZN(
        \DLX_Datapath/RegisterFile/N26431 ) );
  AOI22_X1 U80804 ( .A1(n105583), .A2(n110425), .B1(n105581), .B2(n81320), 
        .ZN(n94825) );
  AOI22_X1 U80806 ( .A1(n105583), .A2(n110103), .B1(n105580), .B2(n81604), 
        .ZN(n94826) );
  OAI21_X1 U80807 ( .B1(n107396), .B2(n105585), .A(n94827), .ZN(
        \DLX_Datapath/RegisterFile/N26429 ) );
  AOI22_X1 U80808 ( .A1(n105583), .A2(n110210), .B1(n105581), .B2(n81405), 
        .ZN(n94827) );
  OAI21_X1 U80809 ( .B1(n107398), .B2(n105585), .A(n94828), .ZN(
        \DLX_Datapath/RegisterFile/N26428 ) );
  AOI22_X1 U80810 ( .A1(n105583), .A2(n109995), .B1(n105580), .B2(n81402), 
        .ZN(n94828) );
  OAI21_X1 U80811 ( .B1(n107400), .B2(n105585), .A(n94829), .ZN(
        \DLX_Datapath/RegisterFile/N26427 ) );
  AOI22_X1 U80812 ( .A1(n105583), .A2(n109878), .B1(n105581), .B2(n81400), 
        .ZN(n94829) );
  OAI21_X1 U80813 ( .B1(n107402), .B2(n105585), .A(n94830), .ZN(
        \DLX_Datapath/RegisterFile/N26426 ) );
  AOI22_X1 U80814 ( .A1(n105583), .A2(n108252), .B1(n105580), .B2(n81332), 
        .ZN(n94830) );
  OAI21_X1 U80815 ( .B1(n107404), .B2(n105585), .A(n94831), .ZN(
        \DLX_Datapath/RegisterFile/N26425 ) );
  AOI22_X1 U80816 ( .A1(n105583), .A2(n108375), .B1(n105581), .B2(n81373), 
        .ZN(n94831) );
  OAI21_X1 U80817 ( .B1(n107406), .B2(n105586), .A(n94832), .ZN(
        \DLX_Datapath/RegisterFile/N26424 ) );
  AOI22_X1 U80818 ( .A1(n105583), .A2(n108486), .B1(n105580), .B2(n81322), 
        .ZN(n94832) );
  OAI21_X1 U80819 ( .B1(n107408), .B2(n105585), .A(n94833), .ZN(
        \DLX_Datapath/RegisterFile/N26423 ) );
  AOI22_X1 U80820 ( .A1(n105583), .A2(n107723), .B1(n105581), .B2(n81506), 
        .ZN(n94833) );
  OAI21_X1 U80821 ( .B1(n107410), .B2(n105585), .A(n94834), .ZN(
        \DLX_Datapath/RegisterFile/N26422 ) );
  AOI22_X1 U80822 ( .A1(n105582), .A2(n109638), .B1(n105580), .B2(n81313), 
        .ZN(n94834) );
  OAI21_X1 U80823 ( .B1(n107412), .B2(n105586), .A(n94835), .ZN(
        \DLX_Datapath/RegisterFile/N26421 ) );
  AOI22_X1 U80824 ( .A1(n105582), .A2(n108600), .B1(n105579), .B2(n81330), 
        .ZN(n94835) );
  AOI22_X1 U80826 ( .A1(n105582), .A2(n109745), .B1(n105579), .B2(n81425), 
        .ZN(n94836) );
  AOI22_X1 U80828 ( .A1(n105582), .A2(n109530), .B1(n105579), .B2(n81396), 
        .ZN(n94837) );
  OAI21_X1 U80829 ( .B1(n108974), .B2(n105585), .A(n94838), .ZN(
        \DLX_Datapath/RegisterFile/N26418 ) );
  AOI22_X1 U80830 ( .A1(n105582), .A2(n109068), .B1(n105579), .B2(n81590), 
        .ZN(n94838) );
  AOI22_X1 U80832 ( .A1(n105582), .A2(n109415), .B1(n105579), .B2(n81423), 
        .ZN(n94839) );
  OAI21_X1 U80833 ( .B1(n111062), .B2(n105585), .A(n94840), .ZN(
        \DLX_Datapath/RegisterFile/N26416 ) );
  AOI22_X1 U80834 ( .A1(n105582), .A2(n109296), .B1(n105579), .B2(n81511), 
        .ZN(n94840) );
  OAI21_X1 U80835 ( .B1(n111061), .B2(n105585), .A(n94841), .ZN(
        \DLX_Datapath/RegisterFile/N26415 ) );
  AOI22_X1 U80836 ( .A1(n105582), .A2(n109188), .B1(n105579), .B2(n81503), 
        .ZN(n94841) );
  OAI21_X1 U80837 ( .B1(n111060), .B2(n105585), .A(n94842), .ZN(
        \DLX_Datapath/RegisterFile/N26414 ) );
  AOI22_X1 U80838 ( .A1(n105582), .A2(n108723), .B1(n105579), .B2(n81417), 
        .ZN(n94842) );
  OAI21_X1 U80839 ( .B1(n111059), .B2(n105586), .A(n94843), .ZN(
        \DLX_Datapath/RegisterFile/N26413 ) );
  AOI22_X1 U80840 ( .A1(n105582), .A2(n108951), .B1(n105579), .B2(n81500), 
        .ZN(n94843) );
  OAI21_X1 U80841 ( .B1(n111058), .B2(n105585), .A(n94844), .ZN(
        \DLX_Datapath/RegisterFile/N26412 ) );
  AOI22_X1 U80842 ( .A1(n105582), .A2(n108839), .B1(n105579), .B2(n81335), 
        .ZN(n94844) );
  OAI21_X1 U80843 ( .B1(n111057), .B2(n105586), .A(n94845), .ZN(
        \DLX_Datapath/RegisterFile/N26411 ) );
  AOI22_X1 U80844 ( .A1(n105582), .A2(n107189), .B1(n105579), .B2(n81327), 
        .ZN(n94845) );
  NOR2_X1 U80847 ( .A1(n104923), .A2(n94809), .ZN(n94813) );
  AOI21_X1 U80848 ( .B1(n105206), .B2(n94847), .A(n94663), .ZN(n94809) );
  OR2_X1 U80849 ( .A1(n94848), .A2(n94553), .ZN(n94847) );
  NAND2_X1 U80850 ( .A1(n94849), .A2(n94850), .ZN(n94553) );
  NOR2_X1 U80851 ( .A1(n94851), .A2(n94852), .ZN(n94849) );
  OAI21_X1 U80853 ( .B1(n107371), .B2(n105578), .A(n94855), .ZN(
        \DLX_Datapath/RegisterFile/N26410 ) );
  AOI22_X1 U80854 ( .A1(n105577), .A2(n94667), .B1(n106755), .B2(n107933), 
        .ZN(n94855) );
  OAI21_X1 U80855 ( .B1(n107373), .B2(n105578), .A(n94857), .ZN(
        \DLX_Datapath/RegisterFile/N26409 ) );
  AOI22_X1 U80856 ( .A1(n105576), .A2(n94670), .B1(n105185), .B2(n108029), 
        .ZN(n94857) );
  OAI21_X1 U80857 ( .B1(n106832), .B2(n105578), .A(n94858), .ZN(
        \DLX_Datapath/RegisterFile/N26408 ) );
  AOI22_X1 U80858 ( .A1(n105577), .A2(n94672), .B1(n106755), .B2(n107190), 
        .ZN(n94858) );
  OAI21_X1 U80859 ( .B1(n107376), .B2(n105578), .A(n94859), .ZN(
        \DLX_Datapath/RegisterFile/N26407 ) );
  AOI22_X1 U80860 ( .A1(n105576), .A2(n94674), .B1(n105185), .B2(n107838), 
        .ZN(n94859) );
  OAI21_X1 U80861 ( .B1(n107378), .B2(n105578), .A(n94860), .ZN(
        \DLX_Datapath/RegisterFile/N26406 ) );
  AOI22_X1 U80862 ( .A1(n105577), .A2(n94676), .B1(n106755), .B2(n110733), 
        .ZN(n94860) );
  OAI21_X1 U80863 ( .B1(n107380), .B2(n105578), .A(n94861), .ZN(
        \DLX_Datapath/RegisterFile/N26405 ) );
  AOI22_X1 U80864 ( .A1(n105576), .A2(n94678), .B1(n105185), .B2(n108138), 
        .ZN(n94861) );
  OAI21_X1 U80865 ( .B1(n107382), .B2(n105578), .A(n94862), .ZN(
        \DLX_Datapath/RegisterFile/N26404 ) );
  AOI22_X1 U80866 ( .A1(n105577), .A2(n94680), .B1(n106755), .B2(n110836), 
        .ZN(n94862) );
  OAI21_X1 U80867 ( .B1(n107384), .B2(n105578), .A(n94863), .ZN(
        \DLX_Datapath/RegisterFile/N26403 ) );
  AOI22_X1 U80868 ( .A1(n105576), .A2(n94682), .B1(n105185), .B2(n110937), 
        .ZN(n94863) );
  OAI21_X1 U80869 ( .B1(n107386), .B2(n105578), .A(n94864), .ZN(
        \DLX_Datapath/RegisterFile/N26402 ) );
  AOI22_X1 U80870 ( .A1(n105576), .A2(n94684), .B1(n105185), .B2(n110530), 
        .ZN(n94864) );
  OAI21_X1 U80871 ( .B1(n107388), .B2(n105578), .A(n94865), .ZN(
        \DLX_Datapath/RegisterFile/N26401 ) );
  AOI22_X1 U80872 ( .A1(n105577), .A2(n94686), .B1(n106755), .B2(n110315), 
        .ZN(n94865) );
  OAI21_X1 U80873 ( .B1(n107390), .B2(n105578), .A(n94866), .ZN(
        \DLX_Datapath/RegisterFile/N26400 ) );
  AOI22_X1 U80874 ( .A1(n94856), .A2(n94688), .B1(n105184), .B2(n110635), .ZN(
        n94866) );
  OAI21_X1 U80875 ( .B1(n107392), .B2(n105578), .A(n94867), .ZN(
        \DLX_Datapath/RegisterFile/N26399 ) );
  AOI22_X1 U80876 ( .A1(n105577), .A2(n94690), .B1(n105184), .B2(n110424), 
        .ZN(n94867) );
  OAI21_X1 U80877 ( .B1(n107394), .B2(n105578), .A(n94868), .ZN(
        \DLX_Datapath/RegisterFile/N26398 ) );
  AOI22_X1 U80878 ( .A1(n105576), .A2(n94692), .B1(n105184), .B2(n110102), 
        .ZN(n94868) );
  OAI21_X1 U80879 ( .B1(n107396), .B2(n105578), .A(n94869), .ZN(
        \DLX_Datapath/RegisterFile/N26397 ) );
  AOI22_X1 U80880 ( .A1(n94856), .A2(n94694), .B1(n105184), .B2(n110209), .ZN(
        n94869) );
  OAI21_X1 U80881 ( .B1(n107398), .B2(n105578), .A(n94870), .ZN(
        \DLX_Datapath/RegisterFile/N26396 ) );
  AOI22_X1 U80882 ( .A1(n105576), .A2(n94696), .B1(n105184), .B2(n109994), 
        .ZN(n94870) );
  OAI21_X1 U80883 ( .B1(n107400), .B2(n105578), .A(n94871), .ZN(
        \DLX_Datapath/RegisterFile/N26395 ) );
  AOI22_X1 U80884 ( .A1(n94856), .A2(n94698), .B1(n105184), .B2(n109877), .ZN(
        n94871) );
  OAI21_X1 U80885 ( .B1(n107402), .B2(n105578), .A(n94872), .ZN(
        \DLX_Datapath/RegisterFile/N26394 ) );
  AOI22_X1 U80886 ( .A1(n94856), .A2(n94700), .B1(n105184), .B2(n108251), .ZN(
        n94872) );
  OAI21_X1 U80887 ( .B1(n107404), .B2(n105578), .A(n94873), .ZN(
        \DLX_Datapath/RegisterFile/N26393 ) );
  AOI22_X1 U80888 ( .A1(n105577), .A2(n94702), .B1(n105184), .B2(n108374), 
        .ZN(n94873) );
  OAI21_X1 U80889 ( .B1(n107406), .B2(n105578), .A(n94874), .ZN(
        \DLX_Datapath/RegisterFile/N26392 ) );
  AOI22_X1 U80890 ( .A1(n105576), .A2(n94704), .B1(n105184), .B2(n108485), 
        .ZN(n94874) );
  OAI21_X1 U80891 ( .B1(n107408), .B2(n105578), .A(n94875), .ZN(
        \DLX_Datapath/RegisterFile/N26391 ) );
  AOI22_X1 U80892 ( .A1(n105577), .A2(n94706), .B1(n105184), .B2(n107722), 
        .ZN(n94875) );
  OAI21_X1 U80893 ( .B1(n107410), .B2(n105578), .A(n94876), .ZN(
        \DLX_Datapath/RegisterFile/N26390 ) );
  AOI22_X1 U80894 ( .A1(n105577), .A2(n94708), .B1(n105184), .B2(n109637), 
        .ZN(n94876) );
  OAI21_X1 U80895 ( .B1(n107412), .B2(n105578), .A(n94877), .ZN(
        \DLX_Datapath/RegisterFile/N26389 ) );
  AOI22_X1 U80896 ( .A1(n105576), .A2(n94710), .B1(n105185), .B2(n108599), 
        .ZN(n94877) );
  OAI21_X1 U80897 ( .B1(n107367), .B2(n105578), .A(n94878), .ZN(
        \DLX_Datapath/RegisterFile/N26388 ) );
  AOI22_X1 U80898 ( .A1(n105577), .A2(n94712), .B1(n106755), .B2(n109744), 
        .ZN(n94878) );
  OAI21_X1 U80899 ( .B1(n107369), .B2(n105578), .A(n94879), .ZN(
        \DLX_Datapath/RegisterFile/N26387 ) );
  AOI22_X1 U80900 ( .A1(n105576), .A2(n94714), .B1(n105185), .B2(n109529), 
        .ZN(n94879) );
  OAI21_X1 U80901 ( .B1(n108974), .B2(n105578), .A(n94880), .ZN(
        \DLX_Datapath/RegisterFile/N26386 ) );
  AOI22_X1 U80902 ( .A1(n105577), .A2(n81259), .B1(n105185), .B2(n109067), 
        .ZN(n94880) );
  OAI21_X1 U80903 ( .B1(n111063), .B2(n105578), .A(n94881), .ZN(
        \DLX_Datapath/RegisterFile/N26385 ) );
  AOI22_X1 U80904 ( .A1(n105576), .A2(n94717), .B1(n105185), .B2(n109414), 
        .ZN(n94881) );
  OAI21_X1 U80905 ( .B1(n111062), .B2(n105578), .A(n94882), .ZN(
        \DLX_Datapath/RegisterFile/N26384 ) );
  AOI22_X1 U80906 ( .A1(n105577), .A2(n94719), .B1(n105184), .B2(n109295), 
        .ZN(n94882) );
  OAI21_X1 U80907 ( .B1(n111061), .B2(n105578), .A(n94883), .ZN(
        \DLX_Datapath/RegisterFile/N26383 ) );
  AOI22_X1 U80908 ( .A1(n105576), .A2(n94721), .B1(n105185), .B2(n109187), 
        .ZN(n94883) );
  OAI21_X1 U80909 ( .B1(n111060), .B2(n105578), .A(n94884), .ZN(
        \DLX_Datapath/RegisterFile/N26382 ) );
  AOI22_X1 U80910 ( .A1(n105577), .A2(n94723), .B1(n106755), .B2(n108722), 
        .ZN(n94884) );
  OAI21_X1 U80911 ( .B1(n111059), .B2(n105578), .A(n94885), .ZN(
        \DLX_Datapath/RegisterFile/N26381 ) );
  AOI22_X1 U80912 ( .A1(n105576), .A2(n94725), .B1(n105185), .B2(n108950), 
        .ZN(n94885) );
  OAI21_X1 U80913 ( .B1(n111058), .B2(n105578), .A(n94886), .ZN(
        \DLX_Datapath/RegisterFile/N26380 ) );
  AOI22_X1 U80914 ( .A1(n105577), .A2(n94727), .B1(n106755), .B2(n108838), 
        .ZN(n94886) );
  OAI21_X1 U80915 ( .B1(n111057), .B2(n105578), .A(n94887), .ZN(
        \DLX_Datapath/RegisterFile/N26379 ) );
  AOI22_X1 U80916 ( .A1(n105576), .A2(n94729), .B1(n105185), .B2(n107191), 
        .ZN(n94887) );
  OAI21_X1 U80917 ( .B1(n94889), .B2(n94663), .A(n94854), .ZN(n94888) );
  AOI21_X1 U80918 ( .B1(n94732), .B2(n111024), .A(n94366), .ZN(n94889) );
  NOR2_X1 U80919 ( .A1(n94890), .A2(n106754), .ZN(n94856) );
  NAND2_X1 U80922 ( .A1(n94854), .A2(n111024), .ZN(n94890) );
  NAND2_X1 U80923 ( .A1(n105136), .A2(n94892), .ZN(n94854) );
  OAI21_X1 U80926 ( .B1(n107371), .B2(n105574), .A(n94897), .ZN(
        \DLX_Datapath/RegisterFile/N26378 ) );
  AOI22_X1 U80927 ( .A1(n105572), .A2(n107932), .B1(n105569), .B2(n81360), 
        .ZN(n94897) );
  OAI21_X1 U80928 ( .B1(n107373), .B2(n105573), .A(n94900), .ZN(
        \DLX_Datapath/RegisterFile/N26377 ) );
  AOI22_X1 U80929 ( .A1(n105572), .A2(n108028), .B1(n105569), .B2(n94511), 
        .ZN(n94900) );
  OAI21_X1 U80930 ( .B1(n106832), .B2(n105574), .A(n94901), .ZN(
        \DLX_Datapath/RegisterFile/N26376 ) );
  AOI22_X1 U80931 ( .A1(n105572), .A2(n107192), .B1(n105568), .B2(n81539), 
        .ZN(n94901) );
  OAI21_X1 U80932 ( .B1(n107376), .B2(n105573), .A(n94902), .ZN(
        \DLX_Datapath/RegisterFile/N26375 ) );
  AOI22_X1 U80933 ( .A1(n105572), .A2(n107837), .B1(n105569), .B2(n81301), 
        .ZN(n94902) );
  OAI21_X1 U80934 ( .B1(n107378), .B2(n105574), .A(n94903), .ZN(
        \DLX_Datapath/RegisterFile/N26374 ) );
  AOI22_X1 U80935 ( .A1(n105572), .A2(n110732), .B1(n105568), .B2(n81308), 
        .ZN(n94903) );
  OAI21_X1 U80936 ( .B1(n107380), .B2(n105573), .A(n94904), .ZN(
        \DLX_Datapath/RegisterFile/N26373 ) );
  AOI22_X1 U80937 ( .A1(n105572), .A2(n108137), .B1(n105568), .B2(n94516), 
        .ZN(n94904) );
  OAI21_X1 U80938 ( .B1(n107382), .B2(n105574), .A(n94905), .ZN(
        \DLX_Datapath/RegisterFile/N26372 ) );
  AOI22_X1 U80939 ( .A1(n105572), .A2(n110835), .B1(n105568), .B2(n81272), 
        .ZN(n94905) );
  OAI21_X1 U80940 ( .B1(n107384), .B2(n105573), .A(n94906), .ZN(
        \DLX_Datapath/RegisterFile/N26371 ) );
  AOI22_X1 U80941 ( .A1(n105572), .A2(n110936), .B1(n105569), .B2(n94519), 
        .ZN(n94906) );
  OAI21_X1 U80942 ( .B1(n107386), .B2(n105574), .A(n94907), .ZN(
        \DLX_Datapath/RegisterFile/N26370 ) );
  AOI22_X1 U80943 ( .A1(n105571), .A2(n110529), .B1(n105567), .B2(n80192), 
        .ZN(n94907) );
  OAI21_X1 U80944 ( .B1(n107388), .B2(n105574), .A(n94908), .ZN(
        \DLX_Datapath/RegisterFile/N26369 ) );
  AOI22_X1 U80945 ( .A1(n105571), .A2(n110314), .B1(n105567), .B2(n81474), 
        .ZN(n94908) );
  OAI21_X1 U80946 ( .B1(n107390), .B2(n105574), .A(n94909), .ZN(
        \DLX_Datapath/RegisterFile/N26368 ) );
  AOI22_X1 U80947 ( .A1(n105571), .A2(n110634), .B1(n105569), .B2(n94523), 
        .ZN(n94909) );
  OAI21_X1 U80948 ( .B1(n107392), .B2(n105574), .A(n94910), .ZN(
        \DLX_Datapath/RegisterFile/N26367 ) );
  AOI22_X1 U80949 ( .A1(n105571), .A2(n110423), .B1(n105567), .B2(n106061), 
        .ZN(n94910) );
  OAI21_X1 U80950 ( .B1(n107394), .B2(n105574), .A(n94911), .ZN(
        \DLX_Datapath/RegisterFile/N26366 ) );
  AOI22_X1 U80951 ( .A1(n105571), .A2(n110101), .B1(n105567), .B2(n81347), 
        .ZN(n94911) );
  OAI21_X1 U80952 ( .B1(n107396), .B2(n105574), .A(n94912), .ZN(
        \DLX_Datapath/RegisterFile/N26365 ) );
  AOI22_X1 U80953 ( .A1(n105571), .A2(n110208), .B1(n105568), .B2(n94527), 
        .ZN(n94912) );
  OAI21_X1 U80954 ( .B1(n107398), .B2(n105574), .A(n94913), .ZN(
        \DLX_Datapath/RegisterFile/N26364 ) );
  AOI22_X1 U80955 ( .A1(n105571), .A2(n109993), .B1(n105567), .B2(n81297), 
        .ZN(n94913) );
  OAI21_X1 U80956 ( .B1(n107400), .B2(n105574), .A(n94914), .ZN(
        \DLX_Datapath/RegisterFile/N26363 ) );
  AOI22_X1 U80957 ( .A1(n105571), .A2(n109876), .B1(n105569), .B2(n94530), 
        .ZN(n94914) );
  OAI21_X1 U80958 ( .B1(n107402), .B2(n105574), .A(n94915), .ZN(
        \DLX_Datapath/RegisterFile/N26362 ) );
  AOI22_X1 U80959 ( .A1(n105571), .A2(n108250), .B1(n105567), .B2(n81286), 
        .ZN(n94915) );
  OAI21_X1 U80960 ( .B1(n107404), .B2(n105574), .A(n94916), .ZN(
        \DLX_Datapath/RegisterFile/N26361 ) );
  AOI22_X1 U80961 ( .A1(n105571), .A2(n108373), .B1(n105568), .B2(n106169), 
        .ZN(n94916) );
  OAI21_X1 U80962 ( .B1(n107406), .B2(n105574), .A(n94917), .ZN(
        \DLX_Datapath/RegisterFile/N26360 ) );
  AOI22_X1 U80963 ( .A1(n105571), .A2(n108484), .B1(n105567), .B2(n81283), 
        .ZN(n94917) );
  OAI21_X1 U80964 ( .B1(n107408), .B2(n105574), .A(n94918), .ZN(
        \DLX_Datapath/RegisterFile/N26359 ) );
  AOI22_X1 U80965 ( .A1(n105571), .A2(n107721), .B1(n105568), .B2(n81453), 
        .ZN(n94918) );
  OAI21_X1 U80966 ( .B1(n107410), .B2(n105573), .A(n94919), .ZN(
        \DLX_Datapath/RegisterFile/N26358 ) );
  AOI22_X1 U80967 ( .A1(n105570), .A2(n109636), .B1(n105568), .B2(n94536), 
        .ZN(n94919) );
  OAI21_X1 U80968 ( .B1(n107412), .B2(n105573), .A(n94920), .ZN(
        \DLX_Datapath/RegisterFile/N26357 ) );
  AOI22_X1 U80969 ( .A1(n105570), .A2(n108598), .B1(n105567), .B2(n106241), 
        .ZN(n94920) );
  OAI21_X1 U80970 ( .B1(n107367), .B2(n105573), .A(n94921), .ZN(
        \DLX_Datapath/RegisterFile/N26356 ) );
  AOI22_X1 U80971 ( .A1(n105570), .A2(n109743), .B1(n105569), .B2(n81351), 
        .ZN(n94921) );
  OAI21_X1 U80972 ( .B1(n107369), .B2(n105573), .A(n94922), .ZN(
        \DLX_Datapath/RegisterFile/N26355 ) );
  AOI22_X1 U80973 ( .A1(n105570), .A2(n109528), .B1(n105567), .B2(n106020), 
        .ZN(n94922) );
  OAI21_X1 U80974 ( .B1(n108974), .B2(n105573), .A(n94923), .ZN(
        \DLX_Datapath/RegisterFile/N26354 ) );
  AOI22_X1 U80975 ( .A1(n105570), .A2(n109066), .B1(n105569), .B2(n94541), 
        .ZN(n94923) );
  OAI21_X1 U80976 ( .B1(n111063), .B2(n105573), .A(n94924), .ZN(
        \DLX_Datapath/RegisterFile/N26353 ) );
  AOI22_X1 U80977 ( .A1(n105570), .A2(n109413), .B1(n105567), .B2(n81269), 
        .ZN(n94924) );
  OAI21_X1 U80978 ( .B1(n111062), .B2(n105573), .A(n94925), .ZN(
        \DLX_Datapath/RegisterFile/N26352 ) );
  AOI22_X1 U80979 ( .A1(n105570), .A2(n109294), .B1(n105568), .B2(n105624), 
        .ZN(n94925) );
  OAI21_X1 U80980 ( .B1(n111061), .B2(n105573), .A(n94926), .ZN(
        \DLX_Datapath/RegisterFile/N26351 ) );
  AOI22_X1 U80981 ( .A1(n105570), .A2(n109186), .B1(n105569), .B2(n94546), 
        .ZN(n94926) );
  OAI21_X1 U80982 ( .B1(n111060), .B2(n105573), .A(n94927), .ZN(
        \DLX_Datapath/RegisterFile/N26350 ) );
  AOI22_X1 U80983 ( .A1(n105570), .A2(n108721), .B1(n105568), .B2(n94548), 
        .ZN(n94927) );
  OAI21_X1 U80984 ( .B1(n111059), .B2(n105573), .A(n94928), .ZN(
        \DLX_Datapath/RegisterFile/N26349 ) );
  AOI22_X1 U80985 ( .A1(n105570), .A2(n108949), .B1(n105569), .B2(n81783), 
        .ZN(n94928) );
  OAI21_X1 U80986 ( .B1(n111058), .B2(n105573), .A(n94929), .ZN(
        \DLX_Datapath/RegisterFile/N26348 ) );
  AOI22_X1 U80987 ( .A1(n105570), .A2(n108837), .B1(n105567), .B2(n80188), 
        .ZN(n94929) );
  OAI21_X1 U80988 ( .B1(n111057), .B2(n105573), .A(n94930), .ZN(
        \DLX_Datapath/RegisterFile/N26347 ) );
  AOI22_X1 U80989 ( .A1(n105570), .A2(n107193), .B1(n105568), .B2(n81265), 
        .ZN(n94930) );
  NOR2_X1 U80990 ( .A1(n94931), .A2(n105575), .ZN(n94899) );
  AOI21_X1 U80991 ( .B1(n94932), .B2(n94258), .A(n105575), .ZN(n94898) );
  NAND2_X1 U80992 ( .A1(n94933), .A2(n94934), .ZN(n94896) );
  OAI21_X1 U80993 ( .B1(n107371), .B2(n105565), .A(n94936), .ZN(
        \DLX_Datapath/RegisterFile/N26346 ) );
  AOI22_X1 U80994 ( .A1(n105563), .A2(n94559), .B1(n105560), .B2(n107931), 
        .ZN(n94936) );
  OAI21_X1 U80995 ( .B1(n107373), .B2(n105564), .A(n94939), .ZN(
        \DLX_Datapath/RegisterFile/N26345 ) );
  AOI22_X1 U80996 ( .A1(n105562), .A2(n94562), .B1(n105559), .B2(n108027), 
        .ZN(n94939) );
  OAI21_X1 U80997 ( .B1(n106832), .B2(n105565), .A(n94940), .ZN(
        \DLX_Datapath/RegisterFile/N26344 ) );
  AOI22_X1 U80998 ( .A1(n105563), .A2(n94564), .B1(n105560), .B2(n107194), 
        .ZN(n94940) );
  OAI21_X1 U80999 ( .B1(n107376), .B2(n105564), .A(n94941), .ZN(
        \DLX_Datapath/RegisterFile/N26343 ) );
  AOI22_X1 U81000 ( .A1(n105562), .A2(n94566), .B1(n105559), .B2(n107836), 
        .ZN(n94941) );
  OAI21_X1 U81001 ( .B1(n107378), .B2(n105565), .A(n94942), .ZN(
        \DLX_Datapath/RegisterFile/N26342 ) );
  AOI22_X1 U81002 ( .A1(n105563), .A2(n94568), .B1(n105560), .B2(n110731), 
        .ZN(n94942) );
  OAI21_X1 U81003 ( .B1(n107380), .B2(n105564), .A(n94943), .ZN(
        \DLX_Datapath/RegisterFile/N26341 ) );
  AOI22_X1 U81004 ( .A1(n105562), .A2(n94570), .B1(n105559), .B2(n108136), 
        .ZN(n94943) );
  OAI21_X1 U81005 ( .B1(n107382), .B2(n105565), .A(n94944), .ZN(
        \DLX_Datapath/RegisterFile/N26340 ) );
  AOI22_X1 U81006 ( .A1(n105563), .A2(n94572), .B1(n105560), .B2(n110834), 
        .ZN(n94944) );
  OAI21_X1 U81007 ( .B1(n107384), .B2(n105564), .A(n94945), .ZN(
        \DLX_Datapath/RegisterFile/N26339 ) );
  AOI22_X1 U81008 ( .A1(n105562), .A2(n94574), .B1(n105559), .B2(n110935), 
        .ZN(n94945) );
  OAI21_X1 U81009 ( .B1(n107386), .B2(n105565), .A(n94946), .ZN(
        \DLX_Datapath/RegisterFile/N26338 ) );
  AOI22_X1 U81010 ( .A1(n105561), .A2(n94576), .B1(n105558), .B2(n110528), 
        .ZN(n94946) );
  OAI21_X1 U81011 ( .B1(n107388), .B2(n105565), .A(n94947), .ZN(
        \DLX_Datapath/RegisterFile/N26337 ) );
  AOI22_X1 U81012 ( .A1(n105561), .A2(n94578), .B1(n105558), .B2(n110313), 
        .ZN(n94947) );
  OAI21_X1 U81013 ( .B1(n107390), .B2(n105565), .A(n94948), .ZN(
        \DLX_Datapath/RegisterFile/N26336 ) );
  AOI22_X1 U81014 ( .A1(n105561), .A2(n94580), .B1(n105558), .B2(n110633), 
        .ZN(n94948) );
  OAI21_X1 U81015 ( .B1(n107392), .B2(n105565), .A(n94949), .ZN(
        \DLX_Datapath/RegisterFile/N26335 ) );
  AOI22_X1 U81016 ( .A1(n105561), .A2(n94582), .B1(n105558), .B2(n110422), 
        .ZN(n94949) );
  OAI21_X1 U81017 ( .B1(n107394), .B2(n105565), .A(n94950), .ZN(
        \DLX_Datapath/RegisterFile/N26334 ) );
  AOI22_X1 U81018 ( .A1(n105561), .A2(n94584), .B1(n105558), .B2(n110100), 
        .ZN(n94950) );
  OAI21_X1 U81019 ( .B1(n107396), .B2(n105565), .A(n94951), .ZN(
        \DLX_Datapath/RegisterFile/N26333 ) );
  AOI22_X1 U81020 ( .A1(n105561), .A2(n94586), .B1(n105558), .B2(n110207), 
        .ZN(n94951) );
  OAI21_X1 U81021 ( .B1(n107398), .B2(n105565), .A(n94952), .ZN(
        \DLX_Datapath/RegisterFile/N26332 ) );
  AOI22_X1 U81022 ( .A1(n105561), .A2(n94588), .B1(n105558), .B2(n109992), 
        .ZN(n94952) );
  OAI21_X1 U81023 ( .B1(n107400), .B2(n105565), .A(n94953), .ZN(
        \DLX_Datapath/RegisterFile/N26331 ) );
  AOI22_X1 U81024 ( .A1(n105561), .A2(n94590), .B1(n105558), .B2(n109875), 
        .ZN(n94953) );
  OAI21_X1 U81025 ( .B1(n107402), .B2(n105565), .A(n94954), .ZN(
        \DLX_Datapath/RegisterFile/N26330 ) );
  AOI22_X1 U81026 ( .A1(n105561), .A2(n94592), .B1(n105558), .B2(n108249), 
        .ZN(n94954) );
  OAI21_X1 U81027 ( .B1(n107404), .B2(n105565), .A(n94955), .ZN(
        \DLX_Datapath/RegisterFile/N26329 ) );
  AOI22_X1 U81028 ( .A1(n105561), .A2(n94594), .B1(n105558), .B2(n108372), 
        .ZN(n94955) );
  OAI21_X1 U81029 ( .B1(n107406), .B2(n105565), .A(n94956), .ZN(
        \DLX_Datapath/RegisterFile/N26328 ) );
  AOI22_X1 U81030 ( .A1(n105561), .A2(n94596), .B1(n105558), .B2(n108483), 
        .ZN(n94956) );
  OAI21_X1 U81031 ( .B1(n107408), .B2(n105565), .A(n94957), .ZN(
        \DLX_Datapath/RegisterFile/N26327 ) );
  AOI22_X1 U81032 ( .A1(n105562), .A2(n94598), .B1(n105559), .B2(n107720), 
        .ZN(n94957) );
  OAI21_X1 U81033 ( .B1(n107410), .B2(n105564), .A(n94958), .ZN(
        \DLX_Datapath/RegisterFile/N26326 ) );
  AOI22_X1 U81034 ( .A1(n105563), .A2(n94600), .B1(n105560), .B2(n109635), 
        .ZN(n94958) );
  OAI21_X1 U81035 ( .B1(n107412), .B2(n105564), .A(n94959), .ZN(
        \DLX_Datapath/RegisterFile/N26325 ) );
  AOI22_X1 U81036 ( .A1(n105562), .A2(n94602), .B1(n105559), .B2(n108597), 
        .ZN(n94959) );
  OAI21_X1 U81037 ( .B1(n107367), .B2(n105564), .A(n94960), .ZN(
        \DLX_Datapath/RegisterFile/N26324 ) );
  AOI22_X1 U81038 ( .A1(n105563), .A2(n94604), .B1(n105560), .B2(n109742), 
        .ZN(n94960) );
  OAI21_X1 U81039 ( .B1(n107369), .B2(n105564), .A(n94961), .ZN(
        \DLX_Datapath/RegisterFile/N26323 ) );
  AOI22_X1 U81040 ( .A1(n105562), .A2(n94606), .B1(n105559), .B2(n109527), 
        .ZN(n94961) );
  OAI21_X1 U81041 ( .B1(n108974), .B2(n105564), .A(n94962), .ZN(
        \DLX_Datapath/RegisterFile/N26322 ) );
  AOI22_X1 U81042 ( .A1(n105562), .A2(n94608), .B1(n105559), .B2(n109065), 
        .ZN(n94962) );
  OAI21_X1 U81043 ( .B1(n111063), .B2(n105564), .A(n94963), .ZN(
        \DLX_Datapath/RegisterFile/N26321 ) );
  AOI22_X1 U81044 ( .A1(n105563), .A2(n94610), .B1(n105560), .B2(n109412), 
        .ZN(n94963) );
  OAI21_X1 U81045 ( .B1(n111062), .B2(n105564), .A(n94964), .ZN(
        \DLX_Datapath/RegisterFile/N26320 ) );
  AOI22_X1 U81046 ( .A1(n105562), .A2(n94612), .B1(n105559), .B2(n109293), 
        .ZN(n94964) );
  OAI21_X1 U81047 ( .B1(n111061), .B2(n105564), .A(n94965), .ZN(
        \DLX_Datapath/RegisterFile/N26319 ) );
  AOI22_X1 U81048 ( .A1(n105563), .A2(n94614), .B1(n105560), .B2(n109185), 
        .ZN(n94965) );
  OAI21_X1 U81049 ( .B1(n111060), .B2(n105564), .A(n94966), .ZN(
        \DLX_Datapath/RegisterFile/N26318 ) );
  AOI22_X1 U81050 ( .A1(n105562), .A2(n94616), .B1(n105559), .B2(n108720), 
        .ZN(n94966) );
  OAI21_X1 U81051 ( .B1(n111059), .B2(n105564), .A(n94967), .ZN(
        \DLX_Datapath/RegisterFile/N26317 ) );
  AOI22_X1 U81052 ( .A1(n105563), .A2(n94618), .B1(n105560), .B2(n108948), 
        .ZN(n94967) );
  OAI21_X1 U81053 ( .B1(n111058), .B2(n105564), .A(n94968), .ZN(
        \DLX_Datapath/RegisterFile/N26316 ) );
  AOI22_X1 U81054 ( .A1(n105562), .A2(n94620), .B1(n105559), .B2(n108836), 
        .ZN(n94968) );
  OAI21_X1 U81055 ( .B1(n111057), .B2(n105564), .A(n94969), .ZN(
        \DLX_Datapath/RegisterFile/N26315 ) );
  AOI22_X1 U81056 ( .A1(n105563), .A2(n94622), .B1(n105560), .B2(n107195), 
        .ZN(n94969) );
  NOR2_X1 U81057 ( .A1(n94970), .A2(n105566), .ZN(n94938) );
  NOR2_X1 U81058 ( .A1(n94931), .A2(n105566), .ZN(n94937) );
  NAND2_X1 U81059 ( .A1(n104908), .A2(n94296), .ZN(n94935) );
  OAI21_X1 U81060 ( .B1(n107371), .B2(n105953), .A(n94971), .ZN(
        \DLX_Datapath/RegisterFile/N26314 ) );
  AOI22_X1 U81061 ( .A1(n104688), .A2(n107930), .B1(n104963), .B2(n81521), 
        .ZN(n94971) );
  OAI21_X1 U81062 ( .B1(n107373), .B2(n105952), .A(n94972), .ZN(
        \DLX_Datapath/RegisterFile/N26313 ) );
  AOI22_X1 U81063 ( .A1(n104688), .A2(n108026), .B1(n104964), .B2(n81653), 
        .ZN(n94972) );
  OAI21_X1 U81064 ( .B1(n106832), .B2(n105953), .A(n94973), .ZN(
        \DLX_Datapath/RegisterFile/N26312 ) );
  AOI22_X1 U81065 ( .A1(n81682), .A2(n107196), .B1(n104963), .B2(n81380), .ZN(
        n94973) );
  OAI21_X1 U81066 ( .B1(n107376), .B2(n105953), .A(n94974), .ZN(
        \DLX_Datapath/RegisterFile/N26311 ) );
  AOI22_X1 U81067 ( .A1(n81682), .A2(n107835), .B1(n104962), .B2(n81377), .ZN(
        n94974) );
  OAI21_X1 U81068 ( .B1(n107378), .B2(n105953), .A(n94975), .ZN(
        \DLX_Datapath/RegisterFile/N26310 ) );
  AOI22_X1 U81069 ( .A1(n81682), .A2(n110730), .B1(n104962), .B2(n81428), .ZN(
        n94975) );
  OAI21_X1 U81070 ( .B1(n107380), .B2(n105953), .A(n94976), .ZN(
        \DLX_Datapath/RegisterFile/N26309 ) );
  AOI22_X1 U81071 ( .A1(n81682), .A2(n108135), .B1(n104963), .B2(n81410), .ZN(
        n94976) );
  OAI21_X1 U81072 ( .B1(n107382), .B2(n105953), .A(n94977), .ZN(
        \DLX_Datapath/RegisterFile/N26308 ) );
  AOI22_X1 U81073 ( .A1(n104689), .A2(n110833), .B1(n81700), .B2(n104964), 
        .ZN(n94977) );
  OAI21_X1 U81074 ( .B1(n107384), .B2(n105953), .A(n94978), .ZN(
        \DLX_Datapath/RegisterFile/N26307 ) );
  AOI22_X1 U81075 ( .A1(n104689), .A2(n110934), .B1(n104964), .B2(n81632), 
        .ZN(n94978) );
  OAI21_X1 U81076 ( .B1(n107386), .B2(n105953), .A(n94979), .ZN(
        \DLX_Datapath/RegisterFile/N26306 ) );
  AOI22_X1 U81077 ( .A1(n104688), .A2(n110527), .B1(n104963), .B2(n81414), 
        .ZN(n94979) );
  OAI21_X1 U81078 ( .B1(n107388), .B2(n105953), .A(n94980), .ZN(
        \DLX_Datapath/RegisterFile/N26305 ) );
  AOI22_X1 U81079 ( .A1(n104689), .A2(n110312), .B1(n104962), .B2(n81317), 
        .ZN(n94980) );
  OAI21_X1 U81080 ( .B1(n107390), .B2(n105953), .A(n94981), .ZN(
        \DLX_Datapath/RegisterFile/N26304 ) );
  AOI22_X1 U81081 ( .A1(n104688), .A2(n110632), .B1(n104963), .B2(n81386), 
        .ZN(n94981) );
  OAI21_X1 U81082 ( .B1(n107392), .B2(n105953), .A(n94982), .ZN(
        \DLX_Datapath/RegisterFile/N26303 ) );
  AOI22_X1 U81083 ( .A1(n104689), .A2(n110421), .B1(n104962), .B2(n81320), 
        .ZN(n94982) );
  OAI21_X1 U81084 ( .B1(n107394), .B2(n105953), .A(n94983), .ZN(
        \DLX_Datapath/RegisterFile/N26302 ) );
  AOI22_X1 U81085 ( .A1(n104688), .A2(n110099), .B1(n104964), .B2(n81604), 
        .ZN(n94983) );
  OAI21_X1 U81086 ( .B1(n107396), .B2(n105953), .A(n94984), .ZN(
        \DLX_Datapath/RegisterFile/N26301 ) );
  AOI22_X1 U81087 ( .A1(n104688), .A2(n110206), .B1(n104964), .B2(n81405), 
        .ZN(n94984) );
  OAI21_X1 U81088 ( .B1(n107398), .B2(n105953), .A(n94985), .ZN(
        \DLX_Datapath/RegisterFile/N26300 ) );
  AOI22_X1 U81089 ( .A1(n104689), .A2(n109991), .B1(n104963), .B2(n81402), 
        .ZN(n94985) );
  OAI21_X1 U81090 ( .B1(n107400), .B2(n105952), .A(n94986), .ZN(
        \DLX_Datapath/RegisterFile/N26299 ) );
  AOI22_X1 U81091 ( .A1(n81682), .A2(n109874), .B1(n104963), .B2(n81400), .ZN(
        n94986) );
  OAI21_X1 U81092 ( .B1(n107410), .B2(n105952), .A(n94987), .ZN(
        \DLX_Datapath/RegisterFile/N26294 ) );
  AOI22_X1 U81093 ( .A1(n81682), .A2(n109634), .B1(n104962), .B2(n81313), .ZN(
        n94987) );
  OAI21_X1 U81094 ( .B1(n107367), .B2(n105952), .A(n94988), .ZN(
        \DLX_Datapath/RegisterFile/N26292 ) );
  AOI22_X1 U81095 ( .A1(n104689), .A2(n109741), .B1(n104964), .B2(n81425), 
        .ZN(n94988) );
  OAI21_X1 U81096 ( .B1(n107369), .B2(n105952), .A(n94989), .ZN(
        \DLX_Datapath/RegisterFile/N26291 ) );
  AOI22_X1 U81097 ( .A1(n104689), .A2(n109526), .B1(n104963), .B2(n81396), 
        .ZN(n94989) );
  OAI21_X1 U81098 ( .B1(n108974), .B2(n105952), .A(n94990), .ZN(
        \DLX_Datapath/RegisterFile/N26290 ) );
  AOI22_X1 U81099 ( .A1(n104689), .A2(n109064), .B1(n104962), .B2(n81590), 
        .ZN(n94990) );
  OAI21_X1 U81100 ( .B1(n111063), .B2(n105952), .A(n94991), .ZN(
        \DLX_Datapath/RegisterFile/N26289 ) );
  AOI22_X1 U81101 ( .A1(n104688), .A2(n109411), .B1(n104964), .B2(n81423), 
        .ZN(n94991) );
  OAI21_X1 U81102 ( .B1(n111062), .B2(n105952), .A(n94992), .ZN(
        \DLX_Datapath/RegisterFile/N26288 ) );
  AOI22_X1 U81103 ( .A1(n104688), .A2(n109292), .B1(n104962), .B2(n81511), 
        .ZN(n94992) );
  OAI21_X1 U81104 ( .B1(n111061), .B2(n105952), .A(n94993), .ZN(
        \DLX_Datapath/RegisterFile/N26287 ) );
  AOI22_X1 U81105 ( .A1(n104689), .A2(n109184), .B1(n104964), .B2(n81503), 
        .ZN(n94993) );
  OAI21_X1 U81106 ( .B1(n111060), .B2(n105952), .A(n94994), .ZN(
        \DLX_Datapath/RegisterFile/N26286 ) );
  AOI22_X1 U81107 ( .A1(n104688), .A2(n108719), .B1(n104963), .B2(n81417), 
        .ZN(n94994) );
  OAI21_X1 U81108 ( .B1(n111059), .B2(n105952), .A(n94995), .ZN(
        \DLX_Datapath/RegisterFile/N26285 ) );
  AOI22_X1 U81109 ( .A1(n104689), .A2(n108947), .B1(n104962), .B2(n81500), 
        .ZN(n94995) );
  OAI21_X1 U81110 ( .B1(n111058), .B2(n105952), .A(n94996), .ZN(
        \DLX_Datapath/RegisterFile/N26284 ) );
  AOI22_X1 U81111 ( .A1(n104688), .A2(n108835), .B1(n104963), .B2(n81335), 
        .ZN(n94996) );
  OAI21_X1 U81112 ( .B1(n111057), .B2(n105952), .A(n94997), .ZN(
        \DLX_Datapath/RegisterFile/N26283 ) );
  AOI22_X1 U81113 ( .A1(n104688), .A2(n107197), .B1(n104962), .B2(n81327), 
        .ZN(n94997) );
  NOR2_X1 U81115 ( .A1(n94970), .A2(n105954), .ZN(n81682) );
  AOI21_X1 U81116 ( .B1(n105206), .B2(n94931), .A(n94663), .ZN(n94970) );
  OR2_X1 U81117 ( .A1(n94998), .A2(n94999), .ZN(n94931) );
  NAND2_X1 U81118 ( .A1(n104909), .A2(n94331), .ZN(n81680) );
  OAI21_X1 U81119 ( .B1(n107371), .B2(n104993), .A(n95001), .ZN(
        \DLX_Datapath/RegisterFile/N26282 ) );
  AOI22_X1 U81120 ( .A1(n105557), .A2(n94667), .B1(n105039), .B2(n70407), .ZN(
        n95001) );
  OAI21_X1 U81121 ( .B1(n107373), .B2(n104992), .A(n95003), .ZN(
        \DLX_Datapath/RegisterFile/N26281 ) );
  AOI22_X1 U81122 ( .A1(n105556), .A2(n94670), .B1(n105182), .B2(n70549), .ZN(
        n95003) );
  OAI21_X1 U81123 ( .B1(n106832), .B2(n104993), .A(n95004), .ZN(
        \DLX_Datapath/RegisterFile/N26280 ) );
  AOI22_X1 U81124 ( .A1(n105557), .A2(n94672), .B1(n105183), .B2(n69459), .ZN(
        n95004) );
  OAI21_X1 U81125 ( .B1(n107376), .B2(n104992), .A(n95005), .ZN(
        \DLX_Datapath/RegisterFile/N26279 ) );
  AOI22_X1 U81126 ( .A1(n105556), .A2(n94674), .B1(n105039), .B2(n70263), .ZN(
        n95005) );
  OAI21_X1 U81127 ( .B1(n107378), .B2(n104993), .A(n95006), .ZN(
        \DLX_Datapath/RegisterFile/N26278 ) );
  AOI22_X1 U81128 ( .A1(n105557), .A2(n94676), .B1(n105182), .B2(n74109), .ZN(
        n95006) );
  OAI21_X1 U81129 ( .B1(n107380), .B2(n104992), .A(n95007), .ZN(
        \DLX_Datapath/RegisterFile/N26277 ) );
  AOI22_X1 U81130 ( .A1(n105556), .A2(n94678), .B1(n105182), .B2(n70696), .ZN(
        n95007) );
  OAI21_X1 U81131 ( .B1(n107382), .B2(n104993), .A(n95008), .ZN(
        \DLX_Datapath/RegisterFile/N26276 ) );
  AOI22_X1 U81132 ( .A1(n105557), .A2(n94680), .B1(n105038), .B2(n74250), .ZN(
        n95008) );
  OAI21_X1 U81133 ( .B1(n107384), .B2(n104992), .A(n95009), .ZN(
        \DLX_Datapath/RegisterFile/N26275 ) );
  AOI22_X1 U81134 ( .A1(n105556), .A2(n94682), .B1(n105183), .B2(n74390), .ZN(
        n95009) );
  OAI21_X1 U81135 ( .B1(n107386), .B2(n104992), .A(n95010), .ZN(
        \DLX_Datapath/RegisterFile/N26274 ) );
  AOI22_X1 U81136 ( .A1(n105556), .A2(n94684), .B1(n105038), .B2(n73826), .ZN(
        n95010) );
  OAI21_X1 U81137 ( .B1(n107388), .B2(n104993), .A(n95011), .ZN(
        \DLX_Datapath/RegisterFile/N26273 ) );
  AOI22_X1 U81138 ( .A1(n105557), .A2(n94686), .B1(n105183), .B2(n73530), .ZN(
        n95011) );
  AOI22_X1 U81140 ( .A1(n105555), .A2(n94688), .B1(n105038), .B2(n73967), .ZN(
        n95012) );
  OAI21_X1 U81141 ( .B1(n107392), .B2(n104993), .A(n95013), .ZN(
        \DLX_Datapath/RegisterFile/N26271 ) );
  AOI22_X1 U81142 ( .A1(n105555), .A2(n94690), .B1(n105039), .B2(n73679), .ZN(
        n95013) );
  OAI21_X1 U81143 ( .B1(n107394), .B2(n104992), .A(n95014), .ZN(
        \DLX_Datapath/RegisterFile/N26270 ) );
  AOI22_X1 U81144 ( .A1(n105555), .A2(n94692), .B1(n105039), .B2(n73241), .ZN(
        n95014) );
  OAI21_X1 U81145 ( .B1(n107396), .B2(n104993), .A(n95015), .ZN(
        \DLX_Datapath/RegisterFile/N26269 ) );
  AOI22_X1 U81146 ( .A1(n105555), .A2(n94694), .B1(n105039), .B2(n73383), .ZN(
        n95015) );
  OAI21_X1 U81147 ( .B1(n107398), .B2(n104992), .A(n95016), .ZN(
        \DLX_Datapath/RegisterFile/N26268 ) );
  AOI22_X1 U81148 ( .A1(n105555), .A2(n94696), .B1(n105039), .B2(n73099), .ZN(
        n95016) );
  OAI21_X1 U81149 ( .B1(n107400), .B2(n104993), .A(n95017), .ZN(
        \DLX_Datapath/RegisterFile/N26267 ) );
  AOI22_X1 U81150 ( .A1(n105555), .A2(n94698), .B1(n105182), .B2(n72949), .ZN(
        n95017) );
  OAI21_X1 U81151 ( .B1(n107402), .B2(n104992), .A(n95018), .ZN(
        \DLX_Datapath/RegisterFile/N26266 ) );
  AOI22_X1 U81152 ( .A1(n105555), .A2(n94700), .B1(n105039), .B2(n70845), .ZN(
        n95018) );
  OAI21_X1 U81153 ( .B1(n107404), .B2(n104993), .A(n95019), .ZN(
        \DLX_Datapath/RegisterFile/N26265 ) );
  AOI22_X1 U81154 ( .A1(n105555), .A2(n94702), .B1(n105182), .B2(n71004), .ZN(
        n95019) );
  OAI21_X1 U81155 ( .B1(n107406), .B2(n104992), .A(n95020), .ZN(
        \DLX_Datapath/RegisterFile/N26264 ) );
  AOI22_X1 U81156 ( .A1(n105555), .A2(n94704), .B1(n105182), .B2(n71149), .ZN(
        n95020) );
  OAI21_X1 U81157 ( .B1(n107408), .B2(n104993), .A(n95021), .ZN(
        \DLX_Datapath/RegisterFile/N26263 ) );
  AOI22_X1 U81158 ( .A1(n105555), .A2(n94706), .B1(n105038), .B2(n70110), .ZN(
        n95021) );
  OAI21_X1 U81159 ( .B1(n107410), .B2(n104992), .A(n95022), .ZN(
        \DLX_Datapath/RegisterFile/N26262 ) );
  AOI22_X1 U81160 ( .A1(n105555), .A2(n94708), .B1(n105182), .B2(n72639), .ZN(
        n95022) );
  OAI21_X1 U81161 ( .B1(n107412), .B2(n104993), .A(n95023), .ZN(
        \DLX_Datapath/RegisterFile/N26261 ) );
  AOI22_X1 U81162 ( .A1(n105556), .A2(n94710), .B1(n105182), .B2(n71298), .ZN(
        n95023) );
  OAI21_X1 U81163 ( .B1(n107367), .B2(n104992), .A(n95024), .ZN(
        \DLX_Datapath/RegisterFile/N26260 ) );
  AOI22_X1 U81164 ( .A1(n105557), .A2(n94712), .B1(n105039), .B2(n72781), .ZN(
        n95024) );
  OAI21_X1 U81165 ( .B1(n107369), .B2(n104993), .A(n95025), .ZN(
        \DLX_Datapath/RegisterFile/N26259 ) );
  AOI22_X1 U81166 ( .A1(n105556), .A2(n94714), .B1(n105038), .B2(n72491), .ZN(
        n95025) );
  OAI21_X1 U81167 ( .B1(n108974), .B2(n104992), .A(n95026), .ZN(
        \DLX_Datapath/RegisterFile/N26258 ) );
  AOI22_X1 U81168 ( .A1(n105557), .A2(n81259), .B1(n105039), .B2(n71891), .ZN(
        n95026) );
  OAI21_X1 U81169 ( .B1(n111063), .B2(n104992), .A(n95027), .ZN(
        \DLX_Datapath/RegisterFile/N26257 ) );
  AOI22_X1 U81170 ( .A1(n105556), .A2(n94717), .B1(n105182), .B2(n72340), .ZN(
        n95027) );
  OAI21_X1 U81171 ( .B1(n111062), .B2(n104993), .A(n95028), .ZN(
        \DLX_Datapath/RegisterFile/N26256 ) );
  AOI22_X1 U81172 ( .A1(n105557), .A2(n94719), .B1(n105182), .B2(n72189), .ZN(
        n95028) );
  OAI21_X1 U81173 ( .B1(n111061), .B2(n104992), .A(n95029), .ZN(
        \DLX_Datapath/RegisterFile/N26255 ) );
  AOI22_X1 U81174 ( .A1(n105556), .A2(n94721), .B1(n105182), .B2(n72045), .ZN(
        n95029) );
  OAI21_X1 U81175 ( .B1(n111060), .B2(n104993), .A(n95030), .ZN(
        \DLX_Datapath/RegisterFile/N26254 ) );
  AOI22_X1 U81176 ( .A1(n105557), .A2(n94723), .B1(n105039), .B2(n71447), .ZN(
        n95030) );
  OAI21_X1 U81177 ( .B1(n111059), .B2(n104992), .A(n95031), .ZN(
        \DLX_Datapath/RegisterFile/N26253 ) );
  AOI22_X1 U81178 ( .A1(n105556), .A2(n94725), .B1(n105183), .B2(n71742), .ZN(
        n95031) );
  OAI21_X1 U81179 ( .B1(n111058), .B2(n104993), .A(n95032), .ZN(
        \DLX_Datapath/RegisterFile/N26252 ) );
  AOI22_X1 U81180 ( .A1(n105557), .A2(n94727), .B1(n105183), .B2(n71598), .ZN(
        n95032) );
  OAI21_X1 U81181 ( .B1(n111057), .B2(n104993), .A(n95033), .ZN(
        \DLX_Datapath/RegisterFile/N26251 ) );
  AOI22_X1 U81182 ( .A1(n105556), .A2(n94729), .B1(n105039), .B2(n69460), .ZN(
        n95033) );
  OAI21_X1 U81183 ( .B1(n95035), .B2(n94663), .A(n95000), .ZN(n95034) );
  AOI21_X1 U81184 ( .B1(n95036), .B2(n111025), .A(n94366), .ZN(n95035) );
  NAND2_X1 U81186 ( .A1(n95000), .A2(n111025), .ZN(n95037) );
  NAND2_X1 U81187 ( .A1(n104909), .A2(n94367), .ZN(n95000) );
  OAI21_X1 U81188 ( .B1(n107371), .B2(n105553), .A(n95039), .ZN(
        \DLX_Datapath/RegisterFile/N26250 ) );
  AOI22_X1 U81189 ( .A1(n105550), .A2(n81360), .B1(n105547), .B2(n107929), 
        .ZN(n95039) );
  OAI21_X1 U81190 ( .B1(n107373), .B2(n105553), .A(n95042), .ZN(
        \DLX_Datapath/RegisterFile/N26249 ) );
  AOI22_X1 U81191 ( .A1(n105550), .A2(n94511), .B1(n105547), .B2(n108025), 
        .ZN(n95042) );
  OAI21_X1 U81192 ( .B1(n106832), .B2(n105553), .A(n95043), .ZN(
        \DLX_Datapath/RegisterFile/N26248 ) );
  AOI22_X1 U81193 ( .A1(n105551), .A2(n81539), .B1(n105548), .B2(n107198), 
        .ZN(n95043) );
  OAI21_X1 U81194 ( .B1(n107376), .B2(n105553), .A(n95044), .ZN(
        \DLX_Datapath/RegisterFile/N26247 ) );
  AOI22_X1 U81195 ( .A1(n105550), .A2(n81301), .B1(n105547), .B2(n107834), 
        .ZN(n95044) );
  OAI21_X1 U81196 ( .B1(n107378), .B2(n105553), .A(n95045), .ZN(
        \DLX_Datapath/RegisterFile/N26246 ) );
  AOI22_X1 U81197 ( .A1(n105551), .A2(n81308), .B1(n105548), .B2(n110729), 
        .ZN(n95045) );
  OAI21_X1 U81198 ( .B1(n107380), .B2(n105553), .A(n95046), .ZN(
        \DLX_Datapath/RegisterFile/N26245 ) );
  AOI22_X1 U81199 ( .A1(n105551), .A2(n94516), .B1(n105548), .B2(n108134), 
        .ZN(n95046) );
  OAI21_X1 U81200 ( .B1(n107382), .B2(n105553), .A(n95047), .ZN(
        \DLX_Datapath/RegisterFile/N26244 ) );
  AOI22_X1 U81201 ( .A1(n105551), .A2(n81272), .B1(n105548), .B2(n110832), 
        .ZN(n95047) );
  OAI21_X1 U81202 ( .B1(n107384), .B2(n105553), .A(n95048), .ZN(
        \DLX_Datapath/RegisterFile/N26243 ) );
  AOI22_X1 U81203 ( .A1(n105550), .A2(n94519), .B1(n105547), .B2(n110933), 
        .ZN(n95048) );
  OAI21_X1 U81204 ( .B1(n107386), .B2(n105552), .A(n95049), .ZN(
        \DLX_Datapath/RegisterFile/N26242 ) );
  AOI22_X1 U81205 ( .A1(n105549), .A2(n80192), .B1(n105546), .B2(n110526), 
        .ZN(n95049) );
  OAI21_X1 U81206 ( .B1(n107388), .B2(n105552), .A(n95050), .ZN(
        \DLX_Datapath/RegisterFile/N26241 ) );
  AOI22_X1 U81207 ( .A1(n105550), .A2(n81474), .B1(n105547), .B2(n110311), 
        .ZN(n95050) );
  OAI21_X1 U81208 ( .B1(n107390), .B2(n105552), .A(n95051), .ZN(
        \DLX_Datapath/RegisterFile/N26240 ) );
  AOI22_X1 U81209 ( .A1(n105550), .A2(n94523), .B1(n105547), .B2(n110631), 
        .ZN(n95051) );
  OAI21_X1 U81210 ( .B1(n107392), .B2(n105552), .A(n95052), .ZN(
        \DLX_Datapath/RegisterFile/N26239 ) );
  AOI22_X1 U81211 ( .A1(n105551), .A2(n106060), .B1(n105548), .B2(n110420), 
        .ZN(n95052) );
  OAI21_X1 U81212 ( .B1(n107394), .B2(n105552), .A(n95053), .ZN(
        \DLX_Datapath/RegisterFile/N26238 ) );
  AOI22_X1 U81213 ( .A1(n105549), .A2(n81347), .B1(n105546), .B2(n110098), 
        .ZN(n95053) );
  OAI21_X1 U81214 ( .B1(n107396), .B2(n105552), .A(n95054), .ZN(
        \DLX_Datapath/RegisterFile/N26237 ) );
  AOI22_X1 U81215 ( .A1(n105551), .A2(n94527), .B1(n105548), .B2(n110205), 
        .ZN(n95054) );
  OAI21_X1 U81216 ( .B1(n107398), .B2(n105552), .A(n95055), .ZN(
        \DLX_Datapath/RegisterFile/N26236 ) );
  AOI22_X1 U81217 ( .A1(n105549), .A2(n81297), .B1(n105546), .B2(n109990), 
        .ZN(n95055) );
  OAI21_X1 U81218 ( .B1(n107400), .B2(n105552), .A(n95056), .ZN(
        \DLX_Datapath/RegisterFile/N26235 ) );
  AOI22_X1 U81219 ( .A1(n105550), .A2(n94530), .B1(n105547), .B2(n109873), 
        .ZN(n95056) );
  OAI21_X1 U81220 ( .B1(n107402), .B2(n105552), .A(n95057), .ZN(
        \DLX_Datapath/RegisterFile/N26234 ) );
  AOI22_X1 U81221 ( .A1(n105549), .A2(n81286), .B1(n105546), .B2(n108247), 
        .ZN(n95057) );
  OAI21_X1 U81222 ( .B1(n107404), .B2(n105552), .A(n95058), .ZN(
        \DLX_Datapath/RegisterFile/N26233 ) );
  AOI22_X1 U81223 ( .A1(n105549), .A2(n106167), .B1(n105546), .B2(n108370), 
        .ZN(n95058) );
  OAI21_X1 U81224 ( .B1(n107406), .B2(n105552), .A(n95059), .ZN(
        \DLX_Datapath/RegisterFile/N26232 ) );
  AOI22_X1 U81225 ( .A1(n105549), .A2(n81283), .B1(n105546), .B2(n108481), 
        .ZN(n95059) );
  OAI21_X1 U81226 ( .B1(n107408), .B2(n105552), .A(n95060), .ZN(
        \DLX_Datapath/RegisterFile/N26231 ) );
  AOI22_X1 U81227 ( .A1(n105550), .A2(n81453), .B1(n105547), .B2(n107718), 
        .ZN(n95060) );
  OAI21_X1 U81228 ( .B1(n107410), .B2(n105553), .A(n95061), .ZN(
        \DLX_Datapath/RegisterFile/N26230 ) );
  AOI22_X1 U81229 ( .A1(n105551), .A2(n105626), .B1(n105548), .B2(n109633), 
        .ZN(n95061) );
  OAI21_X1 U81230 ( .B1(n107412), .B2(n105553), .A(n95062), .ZN(
        \DLX_Datapath/RegisterFile/N26229 ) );
  AOI22_X1 U81231 ( .A1(n105549), .A2(n106240), .B1(n105546), .B2(n108595), 
        .ZN(n95062) );
  OAI21_X1 U81232 ( .B1(n107367), .B2(n105553), .A(n95063), .ZN(
        \DLX_Datapath/RegisterFile/N26228 ) );
  AOI22_X1 U81233 ( .A1(n105549), .A2(n81351), .B1(n105546), .B2(n109740), 
        .ZN(n95063) );
  OAI21_X1 U81234 ( .B1(n107369), .B2(n105552), .A(n95064), .ZN(
        \DLX_Datapath/RegisterFile/N26227 ) );
  AOI22_X1 U81235 ( .A1(n105551), .A2(n106019), .B1(n105548), .B2(n109525), 
        .ZN(n95064) );
  OAI21_X1 U81236 ( .B1(n108974), .B2(n105553), .A(n95065), .ZN(
        \DLX_Datapath/RegisterFile/N26226 ) );
  AOI22_X1 U81237 ( .A1(n105550), .A2(n94541), .B1(n105547), .B2(n109063), 
        .ZN(n95065) );
  OAI21_X1 U81238 ( .B1(n111063), .B2(n105553), .A(n95066), .ZN(
        \DLX_Datapath/RegisterFile/N26225 ) );
  AOI22_X1 U81239 ( .A1(n105549), .A2(n81269), .B1(n105546), .B2(n109410), 
        .ZN(n95066) );
  OAI21_X1 U81240 ( .B1(n111062), .B2(n105552), .A(n95067), .ZN(
        \DLX_Datapath/RegisterFile/N26224 ) );
  AOI22_X1 U81241 ( .A1(n105551), .A2(n105623), .B1(n105548), .B2(n109291), 
        .ZN(n95067) );
  OAI21_X1 U81242 ( .B1(n111061), .B2(n105553), .A(n95068), .ZN(
        \DLX_Datapath/RegisterFile/N26223 ) );
  AOI22_X1 U81243 ( .A1(n105550), .A2(n105622), .B1(n105547), .B2(n109183), 
        .ZN(n95068) );
  OAI21_X1 U81244 ( .B1(n111060), .B2(n105552), .A(n95069), .ZN(
        \DLX_Datapath/RegisterFile/N26222 ) );
  AOI22_X1 U81245 ( .A1(n105551), .A2(n105621), .B1(n105548), .B2(n108718), 
        .ZN(n95069) );
  OAI21_X1 U81246 ( .B1(n111059), .B2(n105553), .A(n95070), .ZN(
        \DLX_Datapath/RegisterFile/N26221 ) );
  AOI22_X1 U81247 ( .A1(n105550), .A2(n105911), .B1(n105547), .B2(n108946), 
        .ZN(n95070) );
  OAI21_X1 U81248 ( .B1(n111058), .B2(n105552), .A(n95071), .ZN(
        \DLX_Datapath/RegisterFile/N26220 ) );
  AOI22_X1 U81249 ( .A1(n105549), .A2(n80188), .B1(n105546), .B2(n108834), 
        .ZN(n95071) );
  OAI21_X1 U81250 ( .B1(n111057), .B2(n105553), .A(n95072), .ZN(
        \DLX_Datapath/RegisterFile/N26219 ) );
  AOI22_X1 U81251 ( .A1(n105549), .A2(n81265), .B1(n105546), .B2(n107199), 
        .ZN(n95072) );
  AOI21_X1 U81252 ( .B1(n94932), .B2(n94398), .A(n105554), .ZN(n95041) );
  NOR2_X1 U81253 ( .A1(n95073), .A2(n105554), .ZN(n95040) );
  NAND2_X1 U81254 ( .A1(n94933), .A2(n94399), .ZN(n95038) );
  OAI21_X1 U81255 ( .B1(n107371), .B2(n105544), .A(n95075), .ZN(
        \DLX_Datapath/RegisterFile/N26218 ) );
  AOI22_X1 U81256 ( .A1(n105542), .A2(n94559), .B1(n105539), .B2(n70405), .ZN(
        n95075) );
  OAI21_X1 U81257 ( .B1(n107373), .B2(n105543), .A(n95078), .ZN(
        \DLX_Datapath/RegisterFile/N26217 ) );
  AOI22_X1 U81258 ( .A1(n105541), .A2(n94562), .B1(n105538), .B2(n70547), .ZN(
        n95078) );
  OAI21_X1 U81259 ( .B1(n106832), .B2(n105544), .A(n95079), .ZN(
        \DLX_Datapath/RegisterFile/N26216 ) );
  AOI22_X1 U81260 ( .A1(n105542), .A2(n94564), .B1(n105539), .B2(n69463), .ZN(
        n95079) );
  OAI21_X1 U81261 ( .B1(n107376), .B2(n105543), .A(n95080), .ZN(
        \DLX_Datapath/RegisterFile/N26215 ) );
  AOI22_X1 U81262 ( .A1(n105541), .A2(n94566), .B1(n105538), .B2(n70261), .ZN(
        n95080) );
  OAI21_X1 U81263 ( .B1(n107378), .B2(n105544), .A(n95081), .ZN(
        \DLX_Datapath/RegisterFile/N26214 ) );
  AOI22_X1 U81264 ( .A1(n105542), .A2(n94568), .B1(n105539), .B2(n74107), .ZN(
        n95081) );
  OAI21_X1 U81265 ( .B1(n107380), .B2(n105543), .A(n95082), .ZN(
        \DLX_Datapath/RegisterFile/N26213 ) );
  AOI22_X1 U81266 ( .A1(n105541), .A2(n94570), .B1(n105538), .B2(n70694), .ZN(
        n95082) );
  OAI21_X1 U81267 ( .B1(n107382), .B2(n105544), .A(n95083), .ZN(
        \DLX_Datapath/RegisterFile/N26212 ) );
  AOI22_X1 U81268 ( .A1(n105542), .A2(n94572), .B1(n105539), .B2(n74248), .ZN(
        n95083) );
  OAI21_X1 U81269 ( .B1(n107384), .B2(n105543), .A(n95084), .ZN(
        \DLX_Datapath/RegisterFile/N26211 ) );
  AOI22_X1 U81270 ( .A1(n105541), .A2(n94574), .B1(n105538), .B2(n74388), .ZN(
        n95084) );
  OAI21_X1 U81271 ( .B1(n107386), .B2(n105544), .A(n95085), .ZN(
        \DLX_Datapath/RegisterFile/N26210 ) );
  AOI22_X1 U81272 ( .A1(n105540), .A2(n94576), .B1(n105537), .B2(n73824), .ZN(
        n95085) );
  OAI21_X1 U81273 ( .B1(n107388), .B2(n105544), .A(n95086), .ZN(
        \DLX_Datapath/RegisterFile/N26209 ) );
  AOI22_X1 U81274 ( .A1(n105540), .A2(n94578), .B1(n105537), .B2(n73528), .ZN(
        n95086) );
  OAI21_X1 U81275 ( .B1(n107390), .B2(n105544), .A(n95087), .ZN(
        \DLX_Datapath/RegisterFile/N26208 ) );
  AOI22_X1 U81276 ( .A1(n105540), .A2(n94580), .B1(n105537), .B2(n73965), .ZN(
        n95087) );
  OAI21_X1 U81277 ( .B1(n107392), .B2(n105544), .A(n95088), .ZN(
        \DLX_Datapath/RegisterFile/N26207 ) );
  AOI22_X1 U81278 ( .A1(n105540), .A2(n94582), .B1(n105537), .B2(n73677), .ZN(
        n95088) );
  OAI21_X1 U81279 ( .B1(n107394), .B2(n105544), .A(n95089), .ZN(
        \DLX_Datapath/RegisterFile/N26206 ) );
  AOI22_X1 U81280 ( .A1(n105540), .A2(n94584), .B1(n105537), .B2(n73239), .ZN(
        n95089) );
  OAI21_X1 U81281 ( .B1(n107396), .B2(n105544), .A(n95090), .ZN(
        \DLX_Datapath/RegisterFile/N26205 ) );
  AOI22_X1 U81282 ( .A1(n105540), .A2(n94586), .B1(n105537), .B2(n73381), .ZN(
        n95090) );
  OAI21_X1 U81283 ( .B1(n107398), .B2(n105544), .A(n95091), .ZN(
        \DLX_Datapath/RegisterFile/N26204 ) );
  AOI22_X1 U81284 ( .A1(n105540), .A2(n94588), .B1(n105537), .B2(n73097), .ZN(
        n95091) );
  OAI21_X1 U81285 ( .B1(n107400), .B2(n105544), .A(n95092), .ZN(
        \DLX_Datapath/RegisterFile/N26203 ) );
  AOI22_X1 U81286 ( .A1(n105540), .A2(n94590), .B1(n105537), .B2(n72947), .ZN(
        n95092) );
  OAI21_X1 U81287 ( .B1(n107402), .B2(n105544), .A(n95093), .ZN(
        \DLX_Datapath/RegisterFile/N26202 ) );
  AOI22_X1 U81288 ( .A1(n105540), .A2(n94592), .B1(n105537), .B2(n70843), .ZN(
        n95093) );
  OAI21_X1 U81289 ( .B1(n107404), .B2(n105544), .A(n95094), .ZN(
        \DLX_Datapath/RegisterFile/N26201 ) );
  AOI22_X1 U81290 ( .A1(n105540), .A2(n94594), .B1(n105537), .B2(n71002), .ZN(
        n95094) );
  OAI21_X1 U81291 ( .B1(n107406), .B2(n105544), .A(n95095), .ZN(
        \DLX_Datapath/RegisterFile/N26200 ) );
  AOI22_X1 U81292 ( .A1(n105540), .A2(n94596), .B1(n105537), .B2(n71147), .ZN(
        n95095) );
  OAI21_X1 U81293 ( .B1(n107408), .B2(n105544), .A(n95096), .ZN(
        \DLX_Datapath/RegisterFile/N26199 ) );
  AOI22_X1 U81294 ( .A1(n105541), .A2(n94598), .B1(n105538), .B2(n70108), .ZN(
        n95096) );
  OAI21_X1 U81295 ( .B1(n107410), .B2(n105543), .A(n95097), .ZN(
        \DLX_Datapath/RegisterFile/N26198 ) );
  AOI22_X1 U81296 ( .A1(n105542), .A2(n94600), .B1(n105539), .B2(n72637), .ZN(
        n95097) );
  OAI21_X1 U81297 ( .B1(n107412), .B2(n105543), .A(n95098), .ZN(
        \DLX_Datapath/RegisterFile/N26197 ) );
  AOI22_X1 U81298 ( .A1(n105541), .A2(n94602), .B1(n105538), .B2(n71296), .ZN(
        n95098) );
  OAI21_X1 U81299 ( .B1(n107367), .B2(n105543), .A(n95099), .ZN(
        \DLX_Datapath/RegisterFile/N26196 ) );
  AOI22_X1 U81300 ( .A1(n105542), .A2(n94604), .B1(n105539), .B2(n72779), .ZN(
        n95099) );
  OAI21_X1 U81301 ( .B1(n107369), .B2(n105543), .A(n95100), .ZN(
        \DLX_Datapath/RegisterFile/N26195 ) );
  AOI22_X1 U81302 ( .A1(n105541), .A2(n94606), .B1(n105538), .B2(n72489), .ZN(
        n95100) );
  OAI21_X1 U81303 ( .B1(n108974), .B2(n105543), .A(n95101), .ZN(
        \DLX_Datapath/RegisterFile/N26194 ) );
  AOI22_X1 U81304 ( .A1(n105541), .A2(n94608), .B1(n105538), .B2(n71889), .ZN(
        n95101) );
  OAI21_X1 U81305 ( .B1(n111063), .B2(n105543), .A(n95102), .ZN(
        \DLX_Datapath/RegisterFile/N26193 ) );
  AOI22_X1 U81306 ( .A1(n105542), .A2(n94610), .B1(n105539), .B2(n72338), .ZN(
        n95102) );
  OAI21_X1 U81307 ( .B1(n111062), .B2(n105543), .A(n95103), .ZN(
        \DLX_Datapath/RegisterFile/N26192 ) );
  AOI22_X1 U81308 ( .A1(n105541), .A2(n94612), .B1(n105538), .B2(n72187), .ZN(
        n95103) );
  OAI21_X1 U81309 ( .B1(n111061), .B2(n105543), .A(n95104), .ZN(
        \DLX_Datapath/RegisterFile/N26191 ) );
  AOI22_X1 U81310 ( .A1(n105542), .A2(n94614), .B1(n105539), .B2(n72043), .ZN(
        n95104) );
  OAI21_X1 U81311 ( .B1(n111060), .B2(n105543), .A(n95105), .ZN(
        \DLX_Datapath/RegisterFile/N26190 ) );
  AOI22_X1 U81312 ( .A1(n105541), .A2(n94616), .B1(n105538), .B2(n71445), .ZN(
        n95105) );
  OAI21_X1 U81313 ( .B1(n111059), .B2(n105543), .A(n95106), .ZN(
        \DLX_Datapath/RegisterFile/N26189 ) );
  AOI22_X1 U81314 ( .A1(n105542), .A2(n94618), .B1(n105539), .B2(n71740), .ZN(
        n95106) );
  OAI21_X1 U81315 ( .B1(n111058), .B2(n105543), .A(n95107), .ZN(
        \DLX_Datapath/RegisterFile/N26188 ) );
  AOI22_X1 U81316 ( .A1(n105541), .A2(n94620), .B1(n105538), .B2(n71596), .ZN(
        n95107) );
  OAI21_X1 U81317 ( .B1(n111057), .B2(n105543), .A(n95108), .ZN(
        \DLX_Datapath/RegisterFile/N26187 ) );
  AOI22_X1 U81318 ( .A1(n105542), .A2(n94622), .B1(n105539), .B2(n69464), .ZN(
        n95108) );
  NOR2_X1 U81320 ( .A1(n95073), .A2(n105545), .ZN(n95076) );
  OAI21_X1 U81322 ( .B1(n107384), .B2(n105950), .A(n95110), .ZN(
        \DLX_Datapath/RegisterFile/N26179 ) );
  AOI22_X1 U81323 ( .A1(n74387), .A2(n105948), .B1(n104953), .B2(n81632), .ZN(
        n95110) );
  OAI21_X1 U81324 ( .B1(n107386), .B2(n105950), .A(n95111), .ZN(
        \DLX_Datapath/RegisterFile/N26178 ) );
  AOI22_X1 U81325 ( .A1(n73823), .A2(n105948), .B1(n104953), .B2(n81414), .ZN(
        n95111) );
  OAI21_X1 U81326 ( .B1(n107390), .B2(n105950), .A(n95112), .ZN(
        \DLX_Datapath/RegisterFile/N26176 ) );
  AOI22_X1 U81327 ( .A1(n73964), .A2(n105948), .B1(n104955), .B2(n81386), .ZN(
        n95112) );
  OAI21_X1 U81328 ( .B1(n107398), .B2(n105950), .A(n95113), .ZN(
        \DLX_Datapath/RegisterFile/N26172 ) );
  AOI22_X1 U81329 ( .A1(n73096), .A2(n105948), .B1(n104954), .B2(n81402), .ZN(
        n95113) );
  OAI21_X1 U81330 ( .B1(n107400), .B2(n105950), .A(n95114), .ZN(
        \DLX_Datapath/RegisterFile/N26171 ) );
  AOI22_X1 U81331 ( .A1(n72946), .A2(n105948), .B1(n104954), .B2(n81400), .ZN(
        n95114) );
  OAI21_X1 U81332 ( .B1(n107402), .B2(n105950), .A(n95115), .ZN(
        \DLX_Datapath/RegisterFile/N26170 ) );
  AOI22_X1 U81333 ( .A1(n70842), .A2(n105948), .B1(n104953), .B2(n81332), .ZN(
        n95115) );
  OAI21_X1 U81334 ( .B1(n107404), .B2(n105950), .A(n95116), .ZN(
        \DLX_Datapath/RegisterFile/N26169 ) );
  AOI22_X1 U81335 ( .A1(n71001), .A2(n105948), .B1(n104953), .B2(n81373), .ZN(
        n95116) );
  OAI21_X1 U81336 ( .B1(n107406), .B2(n105950), .A(n95117), .ZN(
        \DLX_Datapath/RegisterFile/N26168 ) );
  AOI22_X1 U81337 ( .A1(n71146), .A2(n105948), .B1(n104955), .B2(n81322), .ZN(
        n95117) );
  OAI21_X1 U81338 ( .B1(n107408), .B2(n105950), .A(n95118), .ZN(
        \DLX_Datapath/RegisterFile/N26167 ) );
  AOI22_X1 U81339 ( .A1(n70107), .A2(n105947), .B1(n104954), .B2(n81506), .ZN(
        n95118) );
  OAI21_X1 U81340 ( .B1(n107410), .B2(n105949), .A(n95119), .ZN(
        \DLX_Datapath/RegisterFile/N26166 ) );
  AOI22_X1 U81341 ( .A1(n72636), .A2(n105946), .B1(n104955), .B2(n81313), .ZN(
        n95119) );
  OAI21_X1 U81342 ( .B1(n107412), .B2(n105949), .A(n95120), .ZN(
        \DLX_Datapath/RegisterFile/N26165 ) );
  AOI22_X1 U81343 ( .A1(n71295), .A2(n105947), .B1(n104953), .B2(n81330), .ZN(
        n95120) );
  OAI21_X1 U81344 ( .B1(n107367), .B2(n105949), .A(n95121), .ZN(
        \DLX_Datapath/RegisterFile/N26164 ) );
  AOI22_X1 U81345 ( .A1(n72778), .A2(n105946), .B1(n104955), .B2(n81425), .ZN(
        n95121) );
  OAI21_X1 U81346 ( .B1(n107369), .B2(n105949), .A(n95122), .ZN(
        \DLX_Datapath/RegisterFile/N26163 ) );
  AOI22_X1 U81347 ( .A1(n72488), .A2(n105947), .B1(n104954), .B2(n81396), .ZN(
        n95122) );
  OAI21_X1 U81348 ( .B1(n108974), .B2(n105949), .A(n95123), .ZN(
        \DLX_Datapath/RegisterFile/N26162 ) );
  AOI22_X1 U81349 ( .A1(n71888), .A2(n105946), .B1(n104954), .B2(n81590), .ZN(
        n95123) );
  OAI21_X1 U81350 ( .B1(n111063), .B2(n105949), .A(n95124), .ZN(
        \DLX_Datapath/RegisterFile/N26161 ) );
  AOI22_X1 U81351 ( .A1(n72337), .A2(n105947), .B1(n104953), .B2(n81423), .ZN(
        n95124) );
  OAI21_X1 U81352 ( .B1(n111062), .B2(n105949), .A(n95125), .ZN(
        \DLX_Datapath/RegisterFile/N26160 ) );
  AOI22_X1 U81353 ( .A1(n72186), .A2(n105946), .B1(n104953), .B2(n81511), .ZN(
        n95125) );
  OAI21_X1 U81354 ( .B1(n111061), .B2(n105949), .A(n95126), .ZN(
        \DLX_Datapath/RegisterFile/N26159 ) );
  AOI22_X1 U81355 ( .A1(n72042), .A2(n105947), .B1(n104955), .B2(n81503), .ZN(
        n95126) );
  OAI21_X1 U81356 ( .B1(n111060), .B2(n105949), .A(n95127), .ZN(
        \DLX_Datapath/RegisterFile/N26158 ) );
  AOI22_X1 U81357 ( .A1(n71444), .A2(n105946), .B1(n104955), .B2(n81417), .ZN(
        n95127) );
  OAI21_X1 U81358 ( .B1(n111059), .B2(n105949), .A(n95128), .ZN(
        \DLX_Datapath/RegisterFile/N26157 ) );
  AOI22_X1 U81359 ( .A1(n71739), .A2(n105947), .B1(n104953), .B2(n81500), .ZN(
        n95128) );
  OAI21_X1 U81360 ( .B1(n111058), .B2(n105949), .A(n95129), .ZN(
        \DLX_Datapath/RegisterFile/N26156 ) );
  AOI22_X1 U81361 ( .A1(n71595), .A2(n105946), .B1(n104954), .B2(n81335), .ZN(
        n95129) );
  OAI21_X1 U81362 ( .B1(n111057), .B2(n105949), .A(n95130), .ZN(
        \DLX_Datapath/RegisterFile/N26155 ) );
  AOI22_X1 U81363 ( .A1(n69466), .A2(n105947), .B1(n104954), .B2(n81327), .ZN(
        n95130) );
  NOR2_X1 U81364 ( .A1(n95073), .A2(n105951), .ZN(n81691) );
  NOR2_X1 U81365 ( .A1(n95109), .A2(n105951), .ZN(n81690) );
  AOI21_X1 U81366 ( .B1(n105206), .B2(n95073), .A(n94663), .ZN(n95109) );
  OR2_X1 U81367 ( .A1(n94998), .A2(n95131), .ZN(n95073) );
  NAND2_X1 U81368 ( .A1(n104908), .A2(n95132), .ZN(n81688) );
  OAI21_X1 U81369 ( .B1(n107371), .B2(n105536), .A(n95134), .ZN(
        \DLX_Datapath/RegisterFile/N26154 ) );
  AOI22_X1 U81370 ( .A1(n105535), .A2(n94667), .B1(n105047), .B2(n107928), 
        .ZN(n95134) );
  OAI21_X1 U81371 ( .B1(n107373), .B2(n105536), .A(n95136), .ZN(
        \DLX_Datapath/RegisterFile/N26153 ) );
  AOI22_X1 U81372 ( .A1(n105534), .A2(n94670), .B1(n105047), .B2(n108024), 
        .ZN(n95136) );
  OAI21_X1 U81373 ( .B1(n106832), .B2(n105536), .A(n95137), .ZN(
        \DLX_Datapath/RegisterFile/N26152 ) );
  AOI22_X1 U81374 ( .A1(n105535), .A2(n94672), .B1(n105181), .B2(n107200), 
        .ZN(n95137) );
  OAI21_X1 U81375 ( .B1(n107376), .B2(n105536), .A(n95138), .ZN(
        \DLX_Datapath/RegisterFile/N26151 ) );
  AOI22_X1 U81376 ( .A1(n105534), .A2(n94674), .B1(n105047), .B2(n107833), 
        .ZN(n95138) );
  OAI21_X1 U81377 ( .B1(n107378), .B2(n105536), .A(n95139), .ZN(
        \DLX_Datapath/RegisterFile/N26150 ) );
  AOI22_X1 U81378 ( .A1(n105535), .A2(n94676), .B1(n105047), .B2(n110728), 
        .ZN(n95139) );
  OAI21_X1 U81379 ( .B1(n107380), .B2(n105536), .A(n95140), .ZN(
        \DLX_Datapath/RegisterFile/N26149 ) );
  AOI22_X1 U81380 ( .A1(n105534), .A2(n94678), .B1(n105046), .B2(n108133), 
        .ZN(n95140) );
  OAI21_X1 U81381 ( .B1(n107382), .B2(n105536), .A(n95141), .ZN(
        \DLX_Datapath/RegisterFile/N26148 ) );
  AOI22_X1 U81382 ( .A1(n105535), .A2(n94680), .B1(n105047), .B2(n110831), 
        .ZN(n95141) );
  OAI21_X1 U81383 ( .B1(n107384), .B2(n105536), .A(n95142), .ZN(
        \DLX_Datapath/RegisterFile/N26147 ) );
  AOI22_X1 U81384 ( .A1(n105534), .A2(n94682), .B1(n105181), .B2(n110932), 
        .ZN(n95142) );
  OAI21_X1 U81385 ( .B1(n107386), .B2(n105536), .A(n95143), .ZN(
        \DLX_Datapath/RegisterFile/N26146 ) );
  AOI22_X1 U81386 ( .A1(n105534), .A2(n94684), .B1(n105047), .B2(n110525), 
        .ZN(n95143) );
  OAI21_X1 U81387 ( .B1(n107388), .B2(n105536), .A(n95144), .ZN(
        \DLX_Datapath/RegisterFile/N26145 ) );
  AOI22_X1 U81388 ( .A1(n105535), .A2(n94686), .B1(n105181), .B2(n110310), 
        .ZN(n95144) );
  OAI21_X1 U81389 ( .B1(n107390), .B2(n105536), .A(n95145), .ZN(
        \DLX_Datapath/RegisterFile/N26144 ) );
  AOI22_X1 U81390 ( .A1(n105533), .A2(n94688), .B1(n105180), .B2(n110630), 
        .ZN(n95145) );
  OAI21_X1 U81391 ( .B1(n107392), .B2(n105536), .A(n95146), .ZN(
        \DLX_Datapath/RegisterFile/N26143 ) );
  AOI22_X1 U81392 ( .A1(n105533), .A2(n94690), .B1(n105180), .B2(n110419), 
        .ZN(n95146) );
  OAI21_X1 U81393 ( .B1(n107394), .B2(n105536), .A(n95147), .ZN(
        \DLX_Datapath/RegisterFile/N26142 ) );
  AOI22_X1 U81394 ( .A1(n105533), .A2(n94692), .B1(n105046), .B2(n110097), 
        .ZN(n95147) );
  OAI21_X1 U81395 ( .B1(n107396), .B2(n105536), .A(n95148), .ZN(
        \DLX_Datapath/RegisterFile/N26141 ) );
  AOI22_X1 U81396 ( .A1(n105533), .A2(n94694), .B1(n105047), .B2(n110204), 
        .ZN(n95148) );
  OAI21_X1 U81397 ( .B1(n107398), .B2(n105536), .A(n95149), .ZN(
        \DLX_Datapath/RegisterFile/N26140 ) );
  AOI22_X1 U81398 ( .A1(n105533), .A2(n94696), .B1(n105047), .B2(n109989), 
        .ZN(n95149) );
  OAI21_X1 U81399 ( .B1(n107400), .B2(n105536), .A(n95150), .ZN(
        \DLX_Datapath/RegisterFile/N26139 ) );
  AOI22_X1 U81400 ( .A1(n105533), .A2(n94698), .B1(n105180), .B2(n109872), 
        .ZN(n95150) );
  OAI21_X1 U81401 ( .B1(n107402), .B2(n105536), .A(n95151), .ZN(
        \DLX_Datapath/RegisterFile/N26138 ) );
  AOI22_X1 U81402 ( .A1(n105533), .A2(n94700), .B1(n105180), .B2(n108246), 
        .ZN(n95151) );
  OAI21_X1 U81403 ( .B1(n107404), .B2(n105536), .A(n95152), .ZN(
        \DLX_Datapath/RegisterFile/N26137 ) );
  AOI22_X1 U81404 ( .A1(n105533), .A2(n94702), .B1(n105181), .B2(n108369), 
        .ZN(n95152) );
  OAI21_X1 U81405 ( .B1(n107406), .B2(n105536), .A(n95153), .ZN(
        \DLX_Datapath/RegisterFile/N26136 ) );
  AOI22_X1 U81406 ( .A1(n105533), .A2(n94704), .B1(n105181), .B2(n108480), 
        .ZN(n95153) );
  OAI21_X1 U81407 ( .B1(n107408), .B2(n105536), .A(n95154), .ZN(
        \DLX_Datapath/RegisterFile/N26135 ) );
  AOI22_X1 U81408 ( .A1(n105533), .A2(n94706), .B1(n105181), .B2(n107717), 
        .ZN(n95154) );
  OAI21_X1 U81409 ( .B1(n107410), .B2(n105536), .A(n95155), .ZN(
        \DLX_Datapath/RegisterFile/N26134 ) );
  AOI22_X1 U81410 ( .A1(n105533), .A2(n94708), .B1(n105180), .B2(n109632), 
        .ZN(n95155) );
  OAI21_X1 U81411 ( .B1(n107412), .B2(n105536), .A(n95156), .ZN(
        \DLX_Datapath/RegisterFile/N26133 ) );
  AOI22_X1 U81412 ( .A1(n105534), .A2(n94710), .B1(n105046), .B2(n108594), 
        .ZN(n95156) );
  OAI21_X1 U81413 ( .B1(n107367), .B2(n105536), .A(n95157), .ZN(
        \DLX_Datapath/RegisterFile/N26132 ) );
  AOI22_X1 U81414 ( .A1(n105535), .A2(n94712), .B1(n105181), .B2(n109739), 
        .ZN(n95157) );
  OAI21_X1 U81415 ( .B1(n107369), .B2(n105536), .A(n95158), .ZN(
        \DLX_Datapath/RegisterFile/N26131 ) );
  AOI22_X1 U81416 ( .A1(n105534), .A2(n94714), .B1(n105047), .B2(n109524), 
        .ZN(n95158) );
  OAI21_X1 U81417 ( .B1(n108974), .B2(n105536), .A(n95159), .ZN(
        \DLX_Datapath/RegisterFile/N26130 ) );
  AOI22_X1 U81418 ( .A1(n105534), .A2(n81259), .B1(n105046), .B2(n109062), 
        .ZN(n95159) );
  OAI21_X1 U81419 ( .B1(n111063), .B2(n105536), .A(n95160), .ZN(
        \DLX_Datapath/RegisterFile/N26129 ) );
  AOI22_X1 U81420 ( .A1(n105535), .A2(n94717), .B1(n105181), .B2(n109409), 
        .ZN(n95160) );
  OAI21_X1 U81421 ( .B1(n111062), .B2(n105536), .A(n95161), .ZN(
        \DLX_Datapath/RegisterFile/N26128 ) );
  AOI22_X1 U81422 ( .A1(n105534), .A2(n94719), .B1(n105047), .B2(n109290), 
        .ZN(n95161) );
  OAI21_X1 U81423 ( .B1(n111061), .B2(n105536), .A(n95162), .ZN(
        \DLX_Datapath/RegisterFile/N26127 ) );
  AOI22_X1 U81424 ( .A1(n105535), .A2(n94721), .B1(n105181), .B2(n109182), 
        .ZN(n95162) );
  OAI21_X1 U81425 ( .B1(n111060), .B2(n105536), .A(n95163), .ZN(
        \DLX_Datapath/RegisterFile/N26126 ) );
  AOI22_X1 U81426 ( .A1(n105534), .A2(n94723), .B1(n105046), .B2(n108717), 
        .ZN(n95163) );
  OAI21_X1 U81427 ( .B1(n111059), .B2(n105536), .A(n95164), .ZN(
        \DLX_Datapath/RegisterFile/N26125 ) );
  AOI22_X1 U81428 ( .A1(n105535), .A2(n94725), .B1(n105047), .B2(n108945), 
        .ZN(n95164) );
  OAI21_X1 U81429 ( .B1(n111058), .B2(n105536), .A(n95165), .ZN(
        \DLX_Datapath/RegisterFile/N26124 ) );
  AOI22_X1 U81430 ( .A1(n105534), .A2(n94727), .B1(n105181), .B2(n108833), 
        .ZN(n95165) );
  OAI21_X1 U81431 ( .B1(n111057), .B2(n105536), .A(n95166), .ZN(
        \DLX_Datapath/RegisterFile/N26123 ) );
  AOI22_X1 U81432 ( .A1(n105535), .A2(n94729), .B1(n105181), .B2(n107201), 
        .ZN(n95166) );
  OAI21_X1 U81433 ( .B1(n95168), .B2(n94663), .A(n95133), .ZN(n95167) );
  AOI21_X1 U81434 ( .B1(n95036), .B2(n111023), .A(n94366), .ZN(n95168) );
  NAND2_X1 U81436 ( .A1(n95133), .A2(n111023), .ZN(n95169) );
  NAND2_X1 U81437 ( .A1(n94933), .A2(n94505), .ZN(n95133) );
  AND2_X2 U81438 ( .A1(n105135), .A2(n94093), .ZN(n94933) );
  OAI21_X1 U81439 ( .B1(n107371), .B2(n105531), .A(n95172), .ZN(
        \DLX_Datapath/RegisterFile/N26122 ) );
  AOI22_X1 U81440 ( .A1(n105529), .A2(n81360), .B1(n105526), .B2(n70402), .ZN(
        n95172) );
  OAI21_X1 U81441 ( .B1(n107373), .B2(n105530), .A(n95175), .ZN(
        \DLX_Datapath/RegisterFile/N26121 ) );
  AOI22_X1 U81442 ( .A1(n105529), .A2(n94511), .B1(n105526), .B2(n70544), .ZN(
        n95175) );
  OAI21_X1 U81443 ( .B1(n106832), .B2(n105531), .A(n95176), .ZN(
        \DLX_Datapath/RegisterFile/N26120 ) );
  AOI22_X1 U81444 ( .A1(n105529), .A2(n81539), .B1(n105526), .B2(n69469), .ZN(
        n95176) );
  OAI21_X1 U81445 ( .B1(n107376), .B2(n105530), .A(n95177), .ZN(
        \DLX_Datapath/RegisterFile/N26119 ) );
  AOI22_X1 U81446 ( .A1(n105529), .A2(n81301), .B1(n105526), .B2(n70258), .ZN(
        n95177) );
  OAI21_X1 U81447 ( .B1(n107378), .B2(n105531), .A(n95178), .ZN(
        \DLX_Datapath/RegisterFile/N26118 ) );
  AOI22_X1 U81448 ( .A1(n105529), .A2(n81308), .B1(n105526), .B2(n74104), .ZN(
        n95178) );
  OAI21_X1 U81449 ( .B1(n107380), .B2(n105530), .A(n95179), .ZN(
        \DLX_Datapath/RegisterFile/N26117 ) );
  AOI22_X1 U81450 ( .A1(n105529), .A2(n94516), .B1(n105526), .B2(n70691), .ZN(
        n95179) );
  OAI21_X1 U81451 ( .B1(n107382), .B2(n105531), .A(n95180), .ZN(
        \DLX_Datapath/RegisterFile/N26116 ) );
  AOI22_X1 U81452 ( .A1(n105529), .A2(n81272), .B1(n105526), .B2(n74245), .ZN(
        n95180) );
  OAI21_X1 U81453 ( .B1(n107384), .B2(n105530), .A(n95181), .ZN(
        \DLX_Datapath/RegisterFile/N26115 ) );
  AOI22_X1 U81454 ( .A1(n105529), .A2(n94519), .B1(n105526), .B2(n74385), .ZN(
        n95181) );
  OAI21_X1 U81455 ( .B1(n107386), .B2(n105531), .A(n95182), .ZN(
        \DLX_Datapath/RegisterFile/N26114 ) );
  AOI22_X1 U81456 ( .A1(n105528), .A2(n80192), .B1(n105525), .B2(n73821), .ZN(
        n95182) );
  OAI21_X1 U81457 ( .B1(n107388), .B2(n105531), .A(n95183), .ZN(
        \DLX_Datapath/RegisterFile/N26113 ) );
  AOI22_X1 U81458 ( .A1(n105528), .A2(n81474), .B1(n105525), .B2(n73525), .ZN(
        n95183) );
  OAI21_X1 U81459 ( .B1(n107390), .B2(n105531), .A(n95184), .ZN(
        \DLX_Datapath/RegisterFile/N26112 ) );
  AOI22_X1 U81460 ( .A1(n105528), .A2(n94523), .B1(n105525), .B2(n73962), .ZN(
        n95184) );
  OAI21_X1 U81461 ( .B1(n107392), .B2(n105531), .A(n95185), .ZN(
        \DLX_Datapath/RegisterFile/N26111 ) );
  AOI22_X1 U81462 ( .A1(n105528), .A2(n106060), .B1(n105525), .B2(n73674), 
        .ZN(n95185) );
  OAI21_X1 U81463 ( .B1(n107394), .B2(n105531), .A(n95186), .ZN(
        \DLX_Datapath/RegisterFile/N26110 ) );
  AOI22_X1 U81464 ( .A1(n105528), .A2(n81347), .B1(n105525), .B2(n73236), .ZN(
        n95186) );
  OAI21_X1 U81465 ( .B1(n107396), .B2(n105531), .A(n95187), .ZN(
        \DLX_Datapath/RegisterFile/N26109 ) );
  AOI22_X1 U81466 ( .A1(n105528), .A2(n94527), .B1(n105525), .B2(n73378), .ZN(
        n95187) );
  OAI21_X1 U81467 ( .B1(n107398), .B2(n105531), .A(n95188), .ZN(
        \DLX_Datapath/RegisterFile/N26108 ) );
  AOI22_X1 U81468 ( .A1(n105528), .A2(n81297), .B1(n105525), .B2(n73094), .ZN(
        n95188) );
  OAI21_X1 U81469 ( .B1(n107400), .B2(n105531), .A(n95189), .ZN(
        \DLX_Datapath/RegisterFile/N26107 ) );
  AOI22_X1 U81470 ( .A1(n105528), .A2(n94530), .B1(n105525), .B2(n72944), .ZN(
        n95189) );
  OAI21_X1 U81471 ( .B1(n107402), .B2(n105531), .A(n95190), .ZN(
        \DLX_Datapath/RegisterFile/N26106 ) );
  AOI22_X1 U81472 ( .A1(n105528), .A2(n81286), .B1(n105525), .B2(n70840), .ZN(
        n95190) );
  OAI21_X1 U81473 ( .B1(n107404), .B2(n105531), .A(n95191), .ZN(
        \DLX_Datapath/RegisterFile/N26105 ) );
  AOI22_X1 U81474 ( .A1(n105528), .A2(n106167), .B1(n105525), .B2(n70999), 
        .ZN(n95191) );
  OAI21_X1 U81475 ( .B1(n107406), .B2(n105531), .A(n95192), .ZN(
        \DLX_Datapath/RegisterFile/N26104 ) );
  AOI22_X1 U81476 ( .A1(n105528), .A2(n81283), .B1(n105525), .B2(n71144), .ZN(
        n95192) );
  OAI21_X1 U81477 ( .B1(n107408), .B2(n105531), .A(n95193), .ZN(
        \DLX_Datapath/RegisterFile/N26103 ) );
  AOI22_X1 U81478 ( .A1(n105528), .A2(n81453), .B1(n105525), .B2(n70105), .ZN(
        n95193) );
  OAI21_X1 U81479 ( .B1(n107410), .B2(n105530), .A(n95194), .ZN(
        \DLX_Datapath/RegisterFile/N26102 ) );
  AOI22_X1 U81480 ( .A1(n105527), .A2(n105626), .B1(n105524), .B2(n72634), 
        .ZN(n95194) );
  OAI21_X1 U81481 ( .B1(n107412), .B2(n105530), .A(n95195), .ZN(
        \DLX_Datapath/RegisterFile/N26101 ) );
  AOI22_X1 U81482 ( .A1(n105527), .A2(n106240), .B1(n105524), .B2(n71293), 
        .ZN(n95195) );
  OAI21_X1 U81483 ( .B1(n107367), .B2(n105530), .A(n95196), .ZN(
        \DLX_Datapath/RegisterFile/N26100 ) );
  AOI22_X1 U81484 ( .A1(n105527), .A2(n81351), .B1(n105524), .B2(n72776), .ZN(
        n95196) );
  OAI21_X1 U81485 ( .B1(n107369), .B2(n105530), .A(n95197), .ZN(
        \DLX_Datapath/RegisterFile/N26099 ) );
  AOI22_X1 U81486 ( .A1(n105527), .A2(n106019), .B1(n105524), .B2(n72486), 
        .ZN(n95197) );
  OAI21_X1 U81487 ( .B1(n108974), .B2(n105530), .A(n95198), .ZN(
        \DLX_Datapath/RegisterFile/N26098 ) );
  AOI22_X1 U81488 ( .A1(n105527), .A2(n94541), .B1(n105524), .B2(n71886), .ZN(
        n95198) );
  OAI21_X1 U81489 ( .B1(n111063), .B2(n105530), .A(n95199), .ZN(
        \DLX_Datapath/RegisterFile/N26097 ) );
  AOI22_X1 U81490 ( .A1(n105527), .A2(n81269), .B1(n105524), .B2(n72335), .ZN(
        n95199) );
  OAI21_X1 U81491 ( .B1(n111062), .B2(n105530), .A(n95200), .ZN(
        \DLX_Datapath/RegisterFile/N26096 ) );
  AOI22_X1 U81492 ( .A1(n105527), .A2(n105623), .B1(n105524), .B2(n72184), 
        .ZN(n95200) );
  OAI21_X1 U81493 ( .B1(n111061), .B2(n105530), .A(n95201), .ZN(
        \DLX_Datapath/RegisterFile/N26095 ) );
  AOI22_X1 U81494 ( .A1(n105527), .A2(n105622), .B1(n105524), .B2(n72040), 
        .ZN(n95201) );
  OAI21_X1 U81495 ( .B1(n111060), .B2(n105530), .A(n95202), .ZN(
        \DLX_Datapath/RegisterFile/N26094 ) );
  AOI22_X1 U81496 ( .A1(n105527), .A2(n105621), .B1(n105524), .B2(n71442), 
        .ZN(n95202) );
  OAI21_X1 U81497 ( .B1(n111059), .B2(n105530), .A(n95203), .ZN(
        \DLX_Datapath/RegisterFile/N26093 ) );
  AOI22_X1 U81498 ( .A1(n105527), .A2(n105911), .B1(n105524), .B2(n71737), 
        .ZN(n95203) );
  OAI21_X1 U81499 ( .B1(n111058), .B2(n105530), .A(n95204), .ZN(
        \DLX_Datapath/RegisterFile/N26092 ) );
  AOI22_X1 U81500 ( .A1(n105527), .A2(n80188), .B1(n105524), .B2(n71593), .ZN(
        n95204) );
  OAI21_X1 U81501 ( .B1(n111057), .B2(n105530), .A(n95205), .ZN(
        \DLX_Datapath/RegisterFile/N26091 ) );
  AOI22_X1 U81502 ( .A1(n105527), .A2(n81265), .B1(n105524), .B2(n69470), .ZN(
        n95205) );
  AOI21_X1 U81503 ( .B1(n94932), .B2(n94554), .A(n105532), .ZN(n95174) );
  NOR2_X1 U81504 ( .A1(n95206), .A2(n105532), .ZN(n95173) );
  NAND2_X1 U81505 ( .A1(n105135), .A2(n94555), .ZN(n95171) );
  OAI21_X1 U81506 ( .B1(n107371), .B2(n105522), .A(n95208), .ZN(
        \DLX_Datapath/RegisterFile/N26090 ) );
  AOI22_X1 U81507 ( .A1(n105520), .A2(n107927), .B1(n105517), .B2(n94559), 
        .ZN(n95208) );
  OAI21_X1 U81508 ( .B1(n107373), .B2(n105521), .A(n95211), .ZN(
        \DLX_Datapath/RegisterFile/N26089 ) );
  AOI22_X1 U81509 ( .A1(n105520), .A2(n108023), .B1(n105517), .B2(n94562), 
        .ZN(n95211) );
  OAI21_X1 U81510 ( .B1(n106832), .B2(n105522), .A(n95212), .ZN(
        \DLX_Datapath/RegisterFile/N26088 ) );
  AOI22_X1 U81511 ( .A1(n105520), .A2(n107202), .B1(n105517), .B2(n94564), 
        .ZN(n95212) );
  OAI21_X1 U81512 ( .B1(n107376), .B2(n105521), .A(n95213), .ZN(
        \DLX_Datapath/RegisterFile/N26087 ) );
  AOI22_X1 U81513 ( .A1(n105520), .A2(n107831), .B1(n105517), .B2(n94566), 
        .ZN(n95213) );
  OAI21_X1 U81514 ( .B1(n107378), .B2(n105522), .A(n95214), .ZN(
        \DLX_Datapath/RegisterFile/N26086 ) );
  AOI22_X1 U81515 ( .A1(n105520), .A2(n110727), .B1(n105517), .B2(n94568), 
        .ZN(n95214) );
  OAI21_X1 U81516 ( .B1(n107380), .B2(n105521), .A(n95215), .ZN(
        \DLX_Datapath/RegisterFile/N26085 ) );
  AOI22_X1 U81517 ( .A1(n105520), .A2(n108131), .B1(n105517), .B2(n94570), 
        .ZN(n95215) );
  OAI21_X1 U81518 ( .B1(n107382), .B2(n105522), .A(n95216), .ZN(
        \DLX_Datapath/RegisterFile/N26084 ) );
  AOI22_X1 U81519 ( .A1(n105520), .A2(n110830), .B1(n105517), .B2(n94572), 
        .ZN(n95216) );
  OAI21_X1 U81520 ( .B1(n107384), .B2(n105521), .A(n95217), .ZN(
        \DLX_Datapath/RegisterFile/N26083 ) );
  AOI22_X1 U81521 ( .A1(n105520), .A2(n110931), .B1(n105517), .B2(n94574), 
        .ZN(n95217) );
  OAI21_X1 U81522 ( .B1(n107386), .B2(n105522), .A(n95218), .ZN(
        \DLX_Datapath/RegisterFile/N26082 ) );
  AOI22_X1 U81523 ( .A1(n105519), .A2(n110524), .B1(n105516), .B2(n94576), 
        .ZN(n95218) );
  OAI21_X1 U81524 ( .B1(n107388), .B2(n105522), .A(n95219), .ZN(
        \DLX_Datapath/RegisterFile/N26081 ) );
  AOI22_X1 U81525 ( .A1(n105519), .A2(n110309), .B1(n105516), .B2(n94578), 
        .ZN(n95219) );
  OAI21_X1 U81526 ( .B1(n107390), .B2(n105522), .A(n95220), .ZN(
        \DLX_Datapath/RegisterFile/N26080 ) );
  AOI22_X1 U81527 ( .A1(n105519), .A2(n110629), .B1(n105516), .B2(n94580), 
        .ZN(n95220) );
  OAI21_X1 U81528 ( .B1(n107392), .B2(n105522), .A(n95221), .ZN(
        \DLX_Datapath/RegisterFile/N26079 ) );
  AOI22_X1 U81529 ( .A1(n105519), .A2(n110418), .B1(n105516), .B2(n94582), 
        .ZN(n95221) );
  OAI21_X1 U81530 ( .B1(n107394), .B2(n105522), .A(n95222), .ZN(
        \DLX_Datapath/RegisterFile/N26078 ) );
  AOI22_X1 U81531 ( .A1(n105519), .A2(n110096), .B1(n105516), .B2(n94584), 
        .ZN(n95222) );
  OAI21_X1 U81532 ( .B1(n107396), .B2(n105522), .A(n95223), .ZN(
        \DLX_Datapath/RegisterFile/N26077 ) );
  AOI22_X1 U81533 ( .A1(n105519), .A2(n110203), .B1(n105516), .B2(n94586), 
        .ZN(n95223) );
  OAI21_X1 U81534 ( .B1(n107398), .B2(n105522), .A(n95224), .ZN(
        \DLX_Datapath/RegisterFile/N26076 ) );
  AOI22_X1 U81535 ( .A1(n105519), .A2(n109988), .B1(n105516), .B2(n94588), 
        .ZN(n95224) );
  OAI21_X1 U81536 ( .B1(n107400), .B2(n105522), .A(n95225), .ZN(
        \DLX_Datapath/RegisterFile/N26075 ) );
  AOI22_X1 U81537 ( .A1(n105519), .A2(n109871), .B1(n105516), .B2(n94590), 
        .ZN(n95225) );
  OAI21_X1 U81538 ( .B1(n107402), .B2(n105522), .A(n95226), .ZN(
        \DLX_Datapath/RegisterFile/N26074 ) );
  AOI22_X1 U81539 ( .A1(n105519), .A2(n108245), .B1(n105516), .B2(n94592), 
        .ZN(n95226) );
  OAI21_X1 U81540 ( .B1(n107404), .B2(n105522), .A(n95227), .ZN(
        \DLX_Datapath/RegisterFile/N26073 ) );
  AOI22_X1 U81541 ( .A1(n105519), .A2(n108368), .B1(n105516), .B2(n94594), 
        .ZN(n95227) );
  OAI21_X1 U81542 ( .B1(n107406), .B2(n105522), .A(n95228), .ZN(
        \DLX_Datapath/RegisterFile/N26072 ) );
  AOI22_X1 U81543 ( .A1(n105519), .A2(n108479), .B1(n105516), .B2(n94596), 
        .ZN(n95228) );
  OAI21_X1 U81544 ( .B1(n107408), .B2(n105522), .A(n95229), .ZN(
        \DLX_Datapath/RegisterFile/N26071 ) );
  AOI22_X1 U81545 ( .A1(n105519), .A2(n107716), .B1(n105516), .B2(n94598), 
        .ZN(n95229) );
  OAI21_X1 U81546 ( .B1(n107410), .B2(n105521), .A(n95230), .ZN(
        \DLX_Datapath/RegisterFile/N26070 ) );
  AOI22_X1 U81547 ( .A1(n105518), .A2(n109631), .B1(n105515), .B2(n94600), 
        .ZN(n95230) );
  OAI21_X1 U81548 ( .B1(n107412), .B2(n105521), .A(n95231), .ZN(
        \DLX_Datapath/RegisterFile/N26069 ) );
  AOI22_X1 U81549 ( .A1(n105518), .A2(n108593), .B1(n105515), .B2(n94602), 
        .ZN(n95231) );
  OAI21_X1 U81550 ( .B1(n107367), .B2(n105521), .A(n95232), .ZN(
        \DLX_Datapath/RegisterFile/N26068 ) );
  AOI22_X1 U81551 ( .A1(n105518), .A2(n109738), .B1(n105515), .B2(n94604), 
        .ZN(n95232) );
  OAI21_X1 U81552 ( .B1(n107369), .B2(n105521), .A(n95233), .ZN(
        \DLX_Datapath/RegisterFile/N26067 ) );
  AOI22_X1 U81553 ( .A1(n105518), .A2(n109523), .B1(n105515), .B2(n94606), 
        .ZN(n95233) );
  OAI21_X1 U81554 ( .B1(n108974), .B2(n105521), .A(n95234), .ZN(
        \DLX_Datapath/RegisterFile/N26066 ) );
  AOI22_X1 U81555 ( .A1(n105518), .A2(n109061), .B1(n105515), .B2(n94608), 
        .ZN(n95234) );
  OAI21_X1 U81556 ( .B1(n111063), .B2(n105521), .A(n95235), .ZN(
        \DLX_Datapath/RegisterFile/N26065 ) );
  AOI22_X1 U81557 ( .A1(n105518), .A2(n109408), .B1(n105515), .B2(n94610), 
        .ZN(n95235) );
  OAI21_X1 U81558 ( .B1(n111062), .B2(n105521), .A(n95236), .ZN(
        \DLX_Datapath/RegisterFile/N26064 ) );
  AOI22_X1 U81559 ( .A1(n105518), .A2(n109289), .B1(n105515), .B2(n94612), 
        .ZN(n95236) );
  OAI21_X1 U81560 ( .B1(n111061), .B2(n105521), .A(n95237), .ZN(
        \DLX_Datapath/RegisterFile/N26063 ) );
  AOI22_X1 U81561 ( .A1(n105518), .A2(n109181), .B1(n105515), .B2(n94614), 
        .ZN(n95237) );
  OAI21_X1 U81562 ( .B1(n111060), .B2(n105521), .A(n95238), .ZN(
        \DLX_Datapath/RegisterFile/N26062 ) );
  AOI22_X1 U81563 ( .A1(n105518), .A2(n108716), .B1(n105515), .B2(n94616), 
        .ZN(n95238) );
  OAI21_X1 U81564 ( .B1(n111059), .B2(n105521), .A(n95239), .ZN(
        \DLX_Datapath/RegisterFile/N26061 ) );
  AOI22_X1 U81565 ( .A1(n105518), .A2(n108944), .B1(n105515), .B2(n94618), 
        .ZN(n95239) );
  OAI21_X1 U81566 ( .B1(n111058), .B2(n105521), .A(n95240), .ZN(
        \DLX_Datapath/RegisterFile/N26060 ) );
  AOI22_X1 U81567 ( .A1(n105518), .A2(n108832), .B1(n105515), .B2(n94620), 
        .ZN(n95240) );
  OAI21_X1 U81568 ( .B1(n111057), .B2(n105521), .A(n95241), .ZN(
        \DLX_Datapath/RegisterFile/N26059 ) );
  AOI22_X1 U81569 ( .A1(n105518), .A2(n107203), .B1(n105515), .B2(n94622), 
        .ZN(n95241) );
  NOR2_X1 U81570 ( .A1(n95206), .A2(n105523), .ZN(n95210) );
  NOR2_X1 U81571 ( .A1(n95242), .A2(n105523), .ZN(n95209) );
  NAND2_X1 U81572 ( .A1(n105135), .A2(n94625), .ZN(n95207) );
  OAI21_X1 U81573 ( .B1(n107371), .B2(n105962), .A(n95243), .ZN(
        \DLX_Datapath/RegisterFile/N26058 ) );
  AOI22_X1 U81574 ( .A1(n105959), .A2(n81521), .B1(n105956), .B2(n107926), 
        .ZN(n95243) );
  OAI21_X1 U81575 ( .B1(n107373), .B2(n105962), .A(n95244), .ZN(
        \DLX_Datapath/RegisterFile/N26057 ) );
  AOI22_X1 U81576 ( .A1(n105959), .A2(n81653), .B1(n105956), .B2(n108022), 
        .ZN(n95244) );
  OAI21_X1 U81577 ( .B1(n106832), .B2(n105962), .A(n95245), .ZN(
        \DLX_Datapath/RegisterFile/N26056 ) );
  AOI22_X1 U81578 ( .A1(n105959), .A2(n81380), .B1(n105956), .B2(n107204), 
        .ZN(n95245) );
  OAI21_X1 U81579 ( .B1(n107376), .B2(n105962), .A(n95246), .ZN(
        \DLX_Datapath/RegisterFile/N26055 ) );
  AOI22_X1 U81580 ( .A1(n105959), .A2(n81377), .B1(n105956), .B2(n107830), 
        .ZN(n95246) );
  OAI21_X1 U81581 ( .B1(n107378), .B2(n105962), .A(n95247), .ZN(
        \DLX_Datapath/RegisterFile/N26054 ) );
  AOI22_X1 U81582 ( .A1(n105959), .A2(n81428), .B1(n105956), .B2(n110726), 
        .ZN(n95247) );
  OAI21_X1 U81583 ( .B1(n107380), .B2(n105962), .A(n95248), .ZN(
        \DLX_Datapath/RegisterFile/N26053 ) );
  AOI22_X1 U81584 ( .A1(n105959), .A2(n81410), .B1(n105956), .B2(n108130), 
        .ZN(n95248) );
  OAI21_X1 U81585 ( .B1(n107382), .B2(n105962), .A(n95249), .ZN(
        \DLX_Datapath/RegisterFile/N26052 ) );
  AOI22_X1 U81586 ( .A1(n81700), .A2(n105958), .B1(n105956), .B2(n110829), 
        .ZN(n95249) );
  OAI21_X1 U81587 ( .B1(n107384), .B2(n105962), .A(n95250), .ZN(
        \DLX_Datapath/RegisterFile/N26051 ) );
  AOI22_X1 U81588 ( .A1(n105959), .A2(n81632), .B1(n105956), .B2(n110930), 
        .ZN(n95250) );
  OAI21_X1 U81589 ( .B1(n107386), .B2(n105962), .A(n95251), .ZN(
        \DLX_Datapath/RegisterFile/N26050 ) );
  AOI22_X1 U81590 ( .A1(n105959), .A2(n81414), .B1(n105956), .B2(n110523), 
        .ZN(n95251) );
  OAI21_X1 U81591 ( .B1(n107388), .B2(n105961), .A(n95252), .ZN(
        \DLX_Datapath/RegisterFile/N26049 ) );
  AOI22_X1 U81592 ( .A1(n105959), .A2(n81317), .B1(n105955), .B2(n110308), 
        .ZN(n95252) );
  OAI21_X1 U81593 ( .B1(n107390), .B2(n105961), .A(n95253), .ZN(
        \DLX_Datapath/RegisterFile/N26048 ) );
  AOI22_X1 U81594 ( .A1(n105959), .A2(n81386), .B1(n105955), .B2(n110628), 
        .ZN(n95253) );
  OAI21_X1 U81595 ( .B1(n107392), .B2(n105961), .A(n95254), .ZN(
        \DLX_Datapath/RegisterFile/N26047 ) );
  AOI22_X1 U81596 ( .A1(n105959), .A2(n81320), .B1(n105955), .B2(n110417), 
        .ZN(n95254) );
  OAI21_X1 U81597 ( .B1(n107394), .B2(n105961), .A(n95255), .ZN(
        \DLX_Datapath/RegisterFile/N26046 ) );
  AOI22_X1 U81598 ( .A1(n105960), .A2(n81604), .B1(n105955), .B2(n110095), 
        .ZN(n95255) );
  OAI21_X1 U81599 ( .B1(n107396), .B2(n105961), .A(n95256), .ZN(
        \DLX_Datapath/RegisterFile/N26045 ) );
  AOI22_X1 U81600 ( .A1(n105960), .A2(n81405), .B1(n105955), .B2(n110202), 
        .ZN(n95256) );
  OAI21_X1 U81601 ( .B1(n107398), .B2(n105961), .A(n95257), .ZN(
        \DLX_Datapath/RegisterFile/N26044 ) );
  AOI22_X1 U81602 ( .A1(n105960), .A2(n81402), .B1(n105955), .B2(n109987), 
        .ZN(n95257) );
  OAI21_X1 U81603 ( .B1(n107400), .B2(n105961), .A(n95258), .ZN(
        \DLX_Datapath/RegisterFile/N26043 ) );
  AOI22_X1 U81604 ( .A1(n105960), .A2(n81400), .B1(n105955), .B2(n109870), 
        .ZN(n95258) );
  OAI21_X1 U81605 ( .B1(n107410), .B2(n105961), .A(n95259), .ZN(
        \DLX_Datapath/RegisterFile/N26038 ) );
  AOI22_X1 U81606 ( .A1(n105960), .A2(n81313), .B1(n105955), .B2(n109630), 
        .ZN(n95259) );
  OAI21_X1 U81607 ( .B1(n107367), .B2(n105961), .A(n95260), .ZN(
        \DLX_Datapath/RegisterFile/N26036 ) );
  AOI22_X1 U81608 ( .A1(n105960), .A2(n81425), .B1(n105955), .B2(n109737), 
        .ZN(n95260) );
  OAI21_X1 U81609 ( .B1(n108974), .B2(n105961), .A(n95261), .ZN(
        \DLX_Datapath/RegisterFile/N26034 ) );
  AOI22_X1 U81610 ( .A1(n105960), .A2(n81590), .B1(n105955), .B2(n109060), 
        .ZN(n95261) );
  OAI21_X1 U81611 ( .B1(n111063), .B2(n105961), .A(n95262), .ZN(
        \DLX_Datapath/RegisterFile/N26033 ) );
  AOI22_X1 U81612 ( .A1(n105960), .A2(n81423), .B1(n105955), .B2(n109407), 
        .ZN(n95262) );
  OAI21_X1 U81613 ( .B1(n111061), .B2(n105961), .A(n95263), .ZN(
        \DLX_Datapath/RegisterFile/N26031 ) );
  AOI22_X1 U81614 ( .A1(n105958), .A2(n81503), .B1(n105955), .B2(n109180), 
        .ZN(n95263) );
  NOR2_X1 U81615 ( .A1(n95242), .A2(n105963), .ZN(n81669) );
  AOI21_X1 U81616 ( .B1(n105206), .B2(n95206), .A(n94663), .ZN(n95242) );
  NOR2_X1 U81617 ( .A1(n95206), .A2(n105963), .ZN(n81668) );
  OR2_X1 U81618 ( .A1(n94998), .A2(n86230), .ZN(n95206) );
  NAND2_X1 U81619 ( .A1(n105135), .A2(n94664), .ZN(n81666) );
  OAI21_X1 U81620 ( .B1(n107371), .B2(n105514), .A(n95265), .ZN(
        \DLX_Datapath/RegisterFile/N26026 ) );
  AOI22_X1 U81621 ( .A1(n95266), .A2(n94667), .B1(n105179), .B2(n107925), .ZN(
        n95265) );
  OAI21_X1 U81622 ( .B1(n107373), .B2(n105514), .A(n95267), .ZN(
        \DLX_Datapath/RegisterFile/N26025 ) );
  AOI22_X1 U81623 ( .A1(n104998), .A2(n94670), .B1(n106750), .B2(n108021), 
        .ZN(n95267) );
  OAI21_X1 U81624 ( .B1(n106832), .B2(n105514), .A(n95268), .ZN(
        \DLX_Datapath/RegisterFile/N26024 ) );
  AOI22_X1 U81625 ( .A1(n95266), .A2(n94672), .B1(n105179), .B2(n107206), .ZN(
        n95268) );
  OAI21_X1 U81626 ( .B1(n107376), .B2(n105514), .A(n95269), .ZN(
        \DLX_Datapath/RegisterFile/N26023 ) );
  AOI22_X1 U81627 ( .A1(n104999), .A2(n94674), .B1(n105178), .B2(n107829), 
        .ZN(n95269) );
  OAI21_X1 U81628 ( .B1(n107378), .B2(n105514), .A(n95270), .ZN(
        \DLX_Datapath/RegisterFile/N26022 ) );
  AOI22_X1 U81629 ( .A1(n104999), .A2(n94676), .B1(n105179), .B2(n110725), 
        .ZN(n95270) );
  OAI21_X1 U81630 ( .B1(n107380), .B2(n105514), .A(n95271), .ZN(
        \DLX_Datapath/RegisterFile/N26021 ) );
  AOI22_X1 U81631 ( .A1(n104998), .A2(n94678), .B1(n105178), .B2(n108129), 
        .ZN(n95271) );
  OAI21_X1 U81632 ( .B1(n107382), .B2(n105514), .A(n95272), .ZN(
        \DLX_Datapath/RegisterFile/N26020 ) );
  AOI22_X1 U81633 ( .A1(n104998), .A2(n94680), .B1(n105179), .B2(n110828), 
        .ZN(n95272) );
  OAI21_X1 U81634 ( .B1(n107384), .B2(n105514), .A(n95273), .ZN(
        \DLX_Datapath/RegisterFile/N26019 ) );
  AOI22_X1 U81635 ( .A1(n104999), .A2(n94682), .B1(n106750), .B2(n110929), 
        .ZN(n95273) );
  OAI21_X1 U81636 ( .B1(n107386), .B2(n105514), .A(n95274), .ZN(
        \DLX_Datapath/RegisterFile/N26018 ) );
  AOI22_X1 U81637 ( .A1(n104998), .A2(n94684), .B1(n106750), .B2(n110522), 
        .ZN(n95274) );
  OAI21_X1 U81638 ( .B1(n107388), .B2(n105514), .A(n95275), .ZN(
        \DLX_Datapath/RegisterFile/N26017 ) );
  AOI22_X1 U81639 ( .A1(n104999), .A2(n94686), .B1(n105179), .B2(n110307), 
        .ZN(n95275) );
  OAI21_X1 U81640 ( .B1(n107390), .B2(n105514), .A(n95276), .ZN(
        \DLX_Datapath/RegisterFile/N26016 ) );
  AOI22_X1 U81641 ( .A1(n95266), .A2(n94688), .B1(n105178), .B2(n110627), .ZN(
        n95276) );
  OAI21_X1 U81642 ( .B1(n107392), .B2(n105514), .A(n95277), .ZN(
        \DLX_Datapath/RegisterFile/N26015 ) );
  AOI22_X1 U81643 ( .A1(n104998), .A2(n94690), .B1(n105178), .B2(n110416), 
        .ZN(n95277) );
  OAI21_X1 U81644 ( .B1(n107394), .B2(n105514), .A(n95278), .ZN(
        \DLX_Datapath/RegisterFile/N26014 ) );
  AOI22_X1 U81645 ( .A1(n104999), .A2(n94692), .B1(n105178), .B2(n110094), 
        .ZN(n95278) );
  OAI21_X1 U81646 ( .B1(n107396), .B2(n105514), .A(n95279), .ZN(
        \DLX_Datapath/RegisterFile/N26013 ) );
  AOI22_X1 U81647 ( .A1(n104999), .A2(n94694), .B1(n105178), .B2(n110201), 
        .ZN(n95279) );
  OAI21_X1 U81648 ( .B1(n107398), .B2(n105514), .A(n95280), .ZN(
        \DLX_Datapath/RegisterFile/N26012 ) );
  AOI22_X1 U81649 ( .A1(n104998), .A2(n94696), .B1(n105178), .B2(n109986), 
        .ZN(n95280) );
  OAI21_X1 U81650 ( .B1(n107400), .B2(n105514), .A(n95281), .ZN(
        \DLX_Datapath/RegisterFile/N26011 ) );
  AOI22_X1 U81651 ( .A1(n95266), .A2(n94698), .B1(n105178), .B2(n109869), .ZN(
        n95281) );
  OAI21_X1 U81652 ( .B1(n107402), .B2(n105514), .A(n95282), .ZN(
        \DLX_Datapath/RegisterFile/N26010 ) );
  AOI22_X1 U81653 ( .A1(n104998), .A2(n94700), .B1(n105178), .B2(n108243), 
        .ZN(n95282) );
  OAI21_X1 U81654 ( .B1(n107404), .B2(n105514), .A(n95283), .ZN(
        \DLX_Datapath/RegisterFile/N26009 ) );
  AOI22_X1 U81655 ( .A1(n104999), .A2(n94702), .B1(n105178), .B2(n108366), 
        .ZN(n95283) );
  OAI21_X1 U81656 ( .B1(n107406), .B2(n105514), .A(n95284), .ZN(
        \DLX_Datapath/RegisterFile/N26008 ) );
  AOI22_X1 U81657 ( .A1(n104998), .A2(n94704), .B1(n105178), .B2(n108477), 
        .ZN(n95284) );
  OAI21_X1 U81658 ( .B1(n107408), .B2(n105514), .A(n95285), .ZN(
        \DLX_Datapath/RegisterFile/N26007 ) );
  AOI22_X1 U81659 ( .A1(n95266), .A2(n94706), .B1(n105178), .B2(n107714), .ZN(
        n95285) );
  OAI21_X1 U81660 ( .B1(n107410), .B2(n105514), .A(n95286), .ZN(
        \DLX_Datapath/RegisterFile/N26006 ) );
  AOI22_X1 U81661 ( .A1(n104998), .A2(n94708), .B1(n105178), .B2(n109629), 
        .ZN(n95286) );
  OAI21_X1 U81662 ( .B1(n107412), .B2(n105514), .A(n95287), .ZN(
        \DLX_Datapath/RegisterFile/N26005 ) );
  AOI22_X1 U81663 ( .A1(n95266), .A2(n94710), .B1(n106750), .B2(n108591), .ZN(
        n95287) );
  OAI21_X1 U81664 ( .B1(n107367), .B2(n105514), .A(n95288), .ZN(
        \DLX_Datapath/RegisterFile/N26004 ) );
  AOI22_X1 U81665 ( .A1(n104999), .A2(n94712), .B1(n105179), .B2(n109736), 
        .ZN(n95288) );
  OAI21_X1 U81666 ( .B1(n107369), .B2(n105514), .A(n95289), .ZN(
        \DLX_Datapath/RegisterFile/N26003 ) );
  AOI22_X1 U81667 ( .A1(n104998), .A2(n94714), .B1(n106750), .B2(n109521), 
        .ZN(n95289) );
  OAI21_X1 U81668 ( .B1(n108974), .B2(n105514), .A(n95290), .ZN(
        \DLX_Datapath/RegisterFile/N26002 ) );
  AOI22_X1 U81669 ( .A1(n104999), .A2(n81259), .B1(n105179), .B2(n109059), 
        .ZN(n95290) );
  OAI21_X1 U81670 ( .B1(n111063), .B2(n105514), .A(n95291), .ZN(
        \DLX_Datapath/RegisterFile/N26001 ) );
  AOI22_X1 U81671 ( .A1(n95266), .A2(n94717), .B1(n106750), .B2(n109406), .ZN(
        n95291) );
  OAI21_X1 U81672 ( .B1(n111062), .B2(n105514), .A(n95292), .ZN(
        \DLX_Datapath/RegisterFile/N26000 ) );
  AOI22_X1 U81673 ( .A1(n104998), .A2(n94719), .B1(n105179), .B2(n109287), 
        .ZN(n95292) );
  OAI21_X1 U81674 ( .B1(n111061), .B2(n105514), .A(n95293), .ZN(
        \DLX_Datapath/RegisterFile/N25999 ) );
  AOI22_X1 U81675 ( .A1(n104998), .A2(n94721), .B1(n105178), .B2(n109179), 
        .ZN(n95293) );
  OAI21_X1 U81676 ( .B1(n111060), .B2(n105514), .A(n95294), .ZN(
        \DLX_Datapath/RegisterFile/N25998 ) );
  AOI22_X1 U81677 ( .A1(n104998), .A2(n94723), .B1(n105179), .B2(n108714), 
        .ZN(n95294) );
  OAI21_X1 U81678 ( .B1(n111059), .B2(n105514), .A(n95295), .ZN(
        \DLX_Datapath/RegisterFile/N25997 ) );
  AOI22_X1 U81679 ( .A1(n104999), .A2(n94725), .B1(n105179), .B2(n108942), 
        .ZN(n95295) );
  OAI21_X1 U81680 ( .B1(n111058), .B2(n105514), .A(n95296), .ZN(
        \DLX_Datapath/RegisterFile/N25996 ) );
  AOI22_X1 U81681 ( .A1(n104998), .A2(n94727), .B1(n105179), .B2(n108830), 
        .ZN(n95296) );
  OAI21_X1 U81682 ( .B1(n111057), .B2(n105514), .A(n95297), .ZN(
        \DLX_Datapath/RegisterFile/N25995 ) );
  AOI22_X1 U81683 ( .A1(n104999), .A2(n94729), .B1(n106750), .B2(n107207), 
        .ZN(n95297) );
  OAI21_X1 U81684 ( .B1(n95299), .B2(n94663), .A(n95264), .ZN(n95298) );
  AOI21_X1 U81685 ( .B1(n95036), .B2(n111026), .A(n94366), .ZN(n95299) );
  NOR2_X1 U81686 ( .A1(n95300), .A2(n106748), .ZN(n95266) );
  NAND2_X1 U81687 ( .A1(n95264), .A2(n111026), .ZN(n95300) );
  NAND2_X1 U81688 ( .A1(n105135), .A2(n94734), .ZN(n95264) );
  OAI21_X1 U81689 ( .B1(n107371), .B2(n105912), .A(n95301), .ZN(
        \DLX_Datapath/RegisterFile/N25994 ) );
  AOI22_X1 U81690 ( .A1(n105909), .A2(n81360), .B1(n105907), .B2(n107924), 
        .ZN(n95301) );
  OAI21_X1 U81691 ( .B1(n107373), .B2(n105913), .A(n95302), .ZN(
        \DLX_Datapath/RegisterFile/N25993 ) );
  AOI22_X1 U81692 ( .A1(n94511), .A2(n105908), .B1(n105907), .B2(n108020), 
        .ZN(n95302) );
  OAI21_X1 U81693 ( .B1(n106832), .B2(n105912), .A(n95303), .ZN(
        \DLX_Datapath/RegisterFile/N25992 ) );
  AOI22_X1 U81694 ( .A1(n105909), .A2(n81539), .B1(n105907), .B2(n107208), 
        .ZN(n95303) );
  OAI21_X1 U81695 ( .B1(n107376), .B2(n105913), .A(n95304), .ZN(
        \DLX_Datapath/RegisterFile/N25991 ) );
  AOI22_X1 U81696 ( .A1(n105909), .A2(n81301), .B1(n105907), .B2(n107828), 
        .ZN(n95304) );
  OAI21_X1 U81697 ( .B1(n107378), .B2(n105912), .A(n95305), .ZN(
        \DLX_Datapath/RegisterFile/N25990 ) );
  AOI22_X1 U81698 ( .A1(n105909), .A2(n81308), .B1(n105907), .B2(n110724), 
        .ZN(n95305) );
  OAI21_X1 U81699 ( .B1(n107380), .B2(n105913), .A(n95306), .ZN(
        \DLX_Datapath/RegisterFile/N25989 ) );
  AOI22_X1 U81700 ( .A1(n94516), .A2(n105908), .B1(n105907), .B2(n108128), 
        .ZN(n95306) );
  OAI21_X1 U81701 ( .B1(n107382), .B2(n105913), .A(n95307), .ZN(
        \DLX_Datapath/RegisterFile/N25988 ) );
  AOI22_X1 U81702 ( .A1(n105909), .A2(n81272), .B1(n105906), .B2(n110827), 
        .ZN(n95307) );
  OAI21_X1 U81703 ( .B1(n107384), .B2(n105913), .A(n95308), .ZN(
        \DLX_Datapath/RegisterFile/N25987 ) );
  AOI22_X1 U81704 ( .A1(n94519), .A2(n105908), .B1(n105906), .B2(n110928), 
        .ZN(n95308) );
  OAI21_X1 U81705 ( .B1(n107386), .B2(n105913), .A(n95309), .ZN(
        \DLX_Datapath/RegisterFile/N25986 ) );
  AOI22_X1 U81706 ( .A1(n105909), .A2(n80192), .B1(n105906), .B2(n110521), 
        .ZN(n95309) );
  OAI21_X1 U81707 ( .B1(n107388), .B2(n105913), .A(n95310), .ZN(
        \DLX_Datapath/RegisterFile/N25985 ) );
  AOI22_X1 U81708 ( .A1(n105909), .A2(n81474), .B1(n105906), .B2(n110306), 
        .ZN(n95310) );
  OAI21_X1 U81709 ( .B1(n107390), .B2(n105913), .A(n95311), .ZN(
        \DLX_Datapath/RegisterFile/N25984 ) );
  AOI22_X1 U81710 ( .A1(n94523), .A2(n105908), .B1(n105906), .B2(n110626), 
        .ZN(n95311) );
  OAI21_X1 U81711 ( .B1(n107392), .B2(n105913), .A(n95312), .ZN(
        \DLX_Datapath/RegisterFile/N25983 ) );
  AOI22_X1 U81712 ( .A1(n105909), .A2(n106060), .B1(n105906), .B2(n110415), 
        .ZN(n95312) );
  OAI21_X1 U81713 ( .B1(n107394), .B2(n105913), .A(n95313), .ZN(
        \DLX_Datapath/RegisterFile/N25982 ) );
  AOI22_X1 U81714 ( .A1(n105909), .A2(n81347), .B1(n105906), .B2(n110093), 
        .ZN(n95313) );
  OAI21_X1 U81715 ( .B1(n107396), .B2(n105913), .A(n95314), .ZN(
        \DLX_Datapath/RegisterFile/N25981 ) );
  AOI22_X1 U81716 ( .A1(n94527), .A2(n105908), .B1(n105906), .B2(n110200), 
        .ZN(n95314) );
  OAI21_X1 U81717 ( .B1(n107398), .B2(n105913), .A(n95315), .ZN(
        \DLX_Datapath/RegisterFile/N25980 ) );
  AOI22_X1 U81718 ( .A1(n105909), .A2(n81297), .B1(n105906), .B2(n109985), 
        .ZN(n95315) );
  OAI21_X1 U81719 ( .B1(n107400), .B2(n105913), .A(n95316), .ZN(
        \DLX_Datapath/RegisterFile/N25979 ) );
  AOI22_X1 U81720 ( .A1(n94530), .A2(n105908), .B1(n105906), .B2(n109868), 
        .ZN(n95316) );
  OAI21_X1 U81721 ( .B1(n107402), .B2(n105913), .A(n95317), .ZN(
        \DLX_Datapath/RegisterFile/N25978 ) );
  AOI22_X1 U81722 ( .A1(n105910), .A2(n81286), .B1(n105906), .B2(n108242), 
        .ZN(n95317) );
  OAI21_X1 U81723 ( .B1(n107404), .B2(n105913), .A(n95318), .ZN(
        \DLX_Datapath/RegisterFile/N25977 ) );
  AOI22_X1 U81724 ( .A1(n105910), .A2(n106167), .B1(n105906), .B2(n108365), 
        .ZN(n95318) );
  OAI21_X1 U81725 ( .B1(n107406), .B2(n105912), .A(n95319), .ZN(
        \DLX_Datapath/RegisterFile/N25976 ) );
  AOI22_X1 U81726 ( .A1(n105910), .A2(n81283), .B1(n105905), .B2(n108476), 
        .ZN(n95319) );
  OAI21_X1 U81727 ( .B1(n107408), .B2(n105912), .A(n95320), .ZN(
        \DLX_Datapath/RegisterFile/N25975 ) );
  AOI22_X1 U81728 ( .A1(n105910), .A2(n81453), .B1(n105905), .B2(n107713), 
        .ZN(n95320) );
  OAI21_X1 U81729 ( .B1(n107410), .B2(n105912), .A(n95321), .ZN(
        \DLX_Datapath/RegisterFile/N25974 ) );
  AOI22_X1 U81730 ( .A1(n105626), .A2(n105908), .B1(n105905), .B2(n109628), 
        .ZN(n95321) );
  OAI21_X1 U81731 ( .B1(n107412), .B2(n105912), .A(n95322), .ZN(
        \DLX_Datapath/RegisterFile/N25973 ) );
  AOI22_X1 U81732 ( .A1(n105910), .A2(n106240), .B1(n105905), .B2(n108590), 
        .ZN(n95322) );
  OAI21_X1 U81733 ( .B1(n107367), .B2(n105912), .A(n95323), .ZN(
        \DLX_Datapath/RegisterFile/N25972 ) );
  AOI22_X1 U81734 ( .A1(n105910), .A2(n81351), .B1(n105905), .B2(n109735), 
        .ZN(n95323) );
  OAI21_X1 U81735 ( .B1(n107369), .B2(n105912), .A(n95324), .ZN(
        \DLX_Datapath/RegisterFile/N25971 ) );
  AOI22_X1 U81736 ( .A1(n105910), .A2(n106019), .B1(n105905), .B2(n109520), 
        .ZN(n95324) );
  OAI21_X1 U81737 ( .B1(n108974), .B2(n105912), .A(n95325), .ZN(
        \DLX_Datapath/RegisterFile/N25970 ) );
  AOI22_X1 U81738 ( .A1(n94541), .A2(n105908), .B1(n105905), .B2(n109058), 
        .ZN(n95325) );
  OAI21_X1 U81739 ( .B1(n111062), .B2(n105912), .A(n95326), .ZN(
        \DLX_Datapath/RegisterFile/N25968 ) );
  AOI22_X1 U81740 ( .A1(n105623), .A2(n105908), .B1(n105905), .B2(n109286), 
        .ZN(n95326) );
  OAI21_X1 U81741 ( .B1(n111061), .B2(n105912), .A(n95327), .ZN(
        \DLX_Datapath/RegisterFile/N25967 ) );
  AOI22_X1 U81742 ( .A1(n105622), .A2(n105908), .B1(n105905), .B2(n109178), 
        .ZN(n95327) );
  OAI21_X1 U81743 ( .B1(n111060), .B2(n105912), .A(n95328), .ZN(
        \DLX_Datapath/RegisterFile/N25966 ) );
  AOI22_X1 U81744 ( .A1(n105621), .A2(n105908), .B1(n105905), .B2(n108713), 
        .ZN(n95328) );
  OAI21_X1 U81745 ( .B1(n111058), .B2(n105912), .A(n95329), .ZN(
        \DLX_Datapath/RegisterFile/N25964 ) );
  AOI22_X1 U81746 ( .A1(n105910), .A2(n80188), .B1(n105905), .B2(n108829), 
        .ZN(n95329) );
  OAI21_X1 U81747 ( .B1(n111057), .B2(n105912), .A(n95330), .ZN(
        \DLX_Datapath/RegisterFile/N25963 ) );
  AOI22_X1 U81748 ( .A1(n105909), .A2(n81265), .B1(n105905), .B2(n107209), 
        .ZN(n95330) );
  AOI21_X1 U81749 ( .B1(n94932), .B2(n94771), .A(n105914), .ZN(n81785) );
  NAND2_X1 U81750 ( .A1(n94998), .A2(n105205), .ZN(n94932) );
  NOR2_X1 U81751 ( .A1(n95331), .A2(n105914), .ZN(n81784) );
  NAND2_X1 U81752 ( .A1(n105135), .A2(n94772), .ZN(n81781) );
  OAI21_X1 U81753 ( .B1(n107371), .B2(n105512), .A(n95333), .ZN(
        \DLX_Datapath/RegisterFile/N25962 ) );
  AOI22_X1 U81754 ( .A1(n105510), .A2(n107923), .B1(n105507), .B2(n94559), 
        .ZN(n95333) );
  OAI21_X1 U81755 ( .B1(n107373), .B2(n105511), .A(n95336), .ZN(
        \DLX_Datapath/RegisterFile/N25961 ) );
  AOI22_X1 U81756 ( .A1(n105510), .A2(n108019), .B1(n105507), .B2(n94562), 
        .ZN(n95336) );
  OAI21_X1 U81757 ( .B1(n106832), .B2(n105512), .A(n95337), .ZN(
        \DLX_Datapath/RegisterFile/N25960 ) );
  AOI22_X1 U81758 ( .A1(n105510), .A2(n107210), .B1(n105507), .B2(n94564), 
        .ZN(n95337) );
  OAI21_X1 U81759 ( .B1(n107376), .B2(n105511), .A(n95338), .ZN(
        \DLX_Datapath/RegisterFile/N25959 ) );
  AOI22_X1 U81760 ( .A1(n105510), .A2(n107827), .B1(n105507), .B2(n94566), 
        .ZN(n95338) );
  OAI21_X1 U81761 ( .B1(n107378), .B2(n105512), .A(n95339), .ZN(
        \DLX_Datapath/RegisterFile/N25958 ) );
  AOI22_X1 U81762 ( .A1(n105510), .A2(n110723), .B1(n105507), .B2(n94568), 
        .ZN(n95339) );
  OAI21_X1 U81763 ( .B1(n107380), .B2(n105511), .A(n95340), .ZN(
        \DLX_Datapath/RegisterFile/N25957 ) );
  AOI22_X1 U81764 ( .A1(n105510), .A2(n108127), .B1(n105507), .B2(n94570), 
        .ZN(n95340) );
  OAI21_X1 U81765 ( .B1(n107382), .B2(n105512), .A(n95341), .ZN(
        \DLX_Datapath/RegisterFile/N25956 ) );
  AOI22_X1 U81766 ( .A1(n105510), .A2(n110826), .B1(n105507), .B2(n94572), 
        .ZN(n95341) );
  OAI21_X1 U81767 ( .B1(n107384), .B2(n105511), .A(n95342), .ZN(
        \DLX_Datapath/RegisterFile/N25955 ) );
  AOI22_X1 U81768 ( .A1(n105510), .A2(n110927), .B1(n105507), .B2(n94574), 
        .ZN(n95342) );
  OAI21_X1 U81769 ( .B1(n107386), .B2(n105512), .A(n95343), .ZN(
        \DLX_Datapath/RegisterFile/N25954 ) );
  AOI22_X1 U81770 ( .A1(n105509), .A2(n110520), .B1(n105506), .B2(n94576), 
        .ZN(n95343) );
  OAI21_X1 U81771 ( .B1(n107388), .B2(n105512), .A(n95344), .ZN(
        \DLX_Datapath/RegisterFile/N25953 ) );
  AOI22_X1 U81772 ( .A1(n105509), .A2(n110305), .B1(n105506), .B2(n94578), 
        .ZN(n95344) );
  OAI21_X1 U81773 ( .B1(n107390), .B2(n105512), .A(n95345), .ZN(
        \DLX_Datapath/RegisterFile/N25952 ) );
  AOI22_X1 U81774 ( .A1(n105509), .A2(n110625), .B1(n105506), .B2(n94580), 
        .ZN(n95345) );
  OAI21_X1 U81775 ( .B1(n107392), .B2(n105512), .A(n95346), .ZN(
        \DLX_Datapath/RegisterFile/N25951 ) );
  AOI22_X1 U81776 ( .A1(n105509), .A2(n110414), .B1(n105506), .B2(n94582), 
        .ZN(n95346) );
  OAI21_X1 U81777 ( .B1(n107394), .B2(n105512), .A(n95347), .ZN(
        \DLX_Datapath/RegisterFile/N25950 ) );
  AOI22_X1 U81778 ( .A1(n105509), .A2(n110092), .B1(n105506), .B2(n94584), 
        .ZN(n95347) );
  OAI21_X1 U81779 ( .B1(n107396), .B2(n105512), .A(n95348), .ZN(
        \DLX_Datapath/RegisterFile/N25949 ) );
  AOI22_X1 U81780 ( .A1(n105509), .A2(n110199), .B1(n105506), .B2(n94586), 
        .ZN(n95348) );
  OAI21_X1 U81781 ( .B1(n107398), .B2(n105512), .A(n95349), .ZN(
        \DLX_Datapath/RegisterFile/N25948 ) );
  AOI22_X1 U81782 ( .A1(n105509), .A2(n109984), .B1(n105506), .B2(n94588), 
        .ZN(n95349) );
  OAI21_X1 U81783 ( .B1(n107400), .B2(n105512), .A(n95350), .ZN(
        \DLX_Datapath/RegisterFile/N25947 ) );
  AOI22_X1 U81784 ( .A1(n105509), .A2(n109867), .B1(n105506), .B2(n94590), 
        .ZN(n95350) );
  OAI21_X1 U81785 ( .B1(n107402), .B2(n105512), .A(n95351), .ZN(
        \DLX_Datapath/RegisterFile/N25946 ) );
  AOI22_X1 U81786 ( .A1(n105509), .A2(n108241), .B1(n105506), .B2(n94592), 
        .ZN(n95351) );
  OAI21_X1 U81787 ( .B1(n107404), .B2(n105512), .A(n95352), .ZN(
        \DLX_Datapath/RegisterFile/N25945 ) );
  AOI22_X1 U81788 ( .A1(n105509), .A2(n108364), .B1(n105506), .B2(n94594), 
        .ZN(n95352) );
  OAI21_X1 U81789 ( .B1(n107406), .B2(n105512), .A(n95353), .ZN(
        \DLX_Datapath/RegisterFile/N25944 ) );
  AOI22_X1 U81790 ( .A1(n105509), .A2(n108475), .B1(n105506), .B2(n94596), 
        .ZN(n95353) );
  OAI21_X1 U81791 ( .B1(n107408), .B2(n105512), .A(n95354), .ZN(
        \DLX_Datapath/RegisterFile/N25943 ) );
  AOI22_X1 U81792 ( .A1(n105509), .A2(n107712), .B1(n105506), .B2(n94598), 
        .ZN(n95354) );
  OAI21_X1 U81793 ( .B1(n107410), .B2(n105511), .A(n95355), .ZN(
        \DLX_Datapath/RegisterFile/N25942 ) );
  AOI22_X1 U81794 ( .A1(n105508), .A2(n109627), .B1(n105505), .B2(n94600), 
        .ZN(n95355) );
  OAI21_X1 U81795 ( .B1(n107412), .B2(n105511), .A(n95356), .ZN(
        \DLX_Datapath/RegisterFile/N25941 ) );
  AOI22_X1 U81796 ( .A1(n105508), .A2(n108589), .B1(n105505), .B2(n94602), 
        .ZN(n95356) );
  OAI21_X1 U81797 ( .B1(n107367), .B2(n105511), .A(n95357), .ZN(
        \DLX_Datapath/RegisterFile/N25940 ) );
  AOI22_X1 U81798 ( .A1(n105508), .A2(n109734), .B1(n105505), .B2(n94604), 
        .ZN(n95357) );
  OAI21_X1 U81799 ( .B1(n107369), .B2(n105511), .A(n95358), .ZN(
        \DLX_Datapath/RegisterFile/N25939 ) );
  AOI22_X1 U81800 ( .A1(n105508), .A2(n109519), .B1(n105505), .B2(n94606), 
        .ZN(n95358) );
  OAI21_X1 U81801 ( .B1(n108974), .B2(n105511), .A(n95359), .ZN(
        \DLX_Datapath/RegisterFile/N25938 ) );
  AOI22_X1 U81802 ( .A1(n105508), .A2(n109057), .B1(n105505), .B2(n94608), 
        .ZN(n95359) );
  OAI21_X1 U81803 ( .B1(n111063), .B2(n105511), .A(n95360), .ZN(
        \DLX_Datapath/RegisterFile/N25937 ) );
  AOI22_X1 U81804 ( .A1(n105508), .A2(n109404), .B1(n105505), .B2(n94610), 
        .ZN(n95360) );
  OAI21_X1 U81805 ( .B1(n111062), .B2(n105511), .A(n95361), .ZN(
        \DLX_Datapath/RegisterFile/N25936 ) );
  AOI22_X1 U81806 ( .A1(n105508), .A2(n109285), .B1(n105505), .B2(n94612), 
        .ZN(n95361) );
  OAI21_X1 U81807 ( .B1(n111061), .B2(n105511), .A(n95362), .ZN(
        \DLX_Datapath/RegisterFile/N25935 ) );
  AOI22_X1 U81808 ( .A1(n105508), .A2(n109177), .B1(n105505), .B2(n94614), 
        .ZN(n95362) );
  OAI21_X1 U81809 ( .B1(n111060), .B2(n105511), .A(n95363), .ZN(
        \DLX_Datapath/RegisterFile/N25934 ) );
  AOI22_X1 U81810 ( .A1(n105508), .A2(n108712), .B1(n105505), .B2(n94616), 
        .ZN(n95363) );
  OAI21_X1 U81811 ( .B1(n111059), .B2(n105511), .A(n95364), .ZN(
        \DLX_Datapath/RegisterFile/N25933 ) );
  AOI22_X1 U81812 ( .A1(n105508), .A2(n108940), .B1(n105505), .B2(n94618), 
        .ZN(n95364) );
  OAI21_X1 U81813 ( .B1(n111058), .B2(n105511), .A(n95365), .ZN(
        \DLX_Datapath/RegisterFile/N25932 ) );
  AOI22_X1 U81814 ( .A1(n105508), .A2(n108828), .B1(n105505), .B2(n94620), 
        .ZN(n95365) );
  OAI21_X1 U81815 ( .B1(n111057), .B2(n105511), .A(n95366), .ZN(
        \DLX_Datapath/RegisterFile/N25931 ) );
  AOI22_X1 U81816 ( .A1(n105508), .A2(n107211), .B1(n105505), .B2(n94622), 
        .ZN(n95366) );
  NOR2_X1 U81817 ( .A1(n95331), .A2(n105513), .ZN(n95335) );
  NOR2_X1 U81818 ( .A1(n105513), .A2(n95367), .ZN(n95334) );
  NAND2_X1 U81819 ( .A1(n105135), .A2(n94810), .ZN(n95332) );
  OAI21_X1 U81820 ( .B1(n107378), .B2(n105943), .A(n95368), .ZN(
        \DLX_Datapath/RegisterFile/N25926 ) );
  AOI22_X1 U81821 ( .A1(n105940), .A2(n81428), .B1(n105937), .B2(n110722), 
        .ZN(n95368) );
  OAI21_X1 U81822 ( .B1(n107382), .B2(n105943), .A(n95369), .ZN(
        \DLX_Datapath/RegisterFile/N25924 ) );
  AOI22_X1 U81823 ( .A1(n105940), .A2(n81700), .B1(n105937), .B2(n110825), 
        .ZN(n95369) );
  OAI21_X1 U81824 ( .B1(n107386), .B2(n105943), .A(n95370), .ZN(
        \DLX_Datapath/RegisterFile/N25922 ) );
  AOI22_X1 U81825 ( .A1(n105940), .A2(n81414), .B1(n105937), .B2(n110519), 
        .ZN(n95370) );
  OAI21_X1 U81826 ( .B1(n107390), .B2(n105943), .A(n95371), .ZN(
        \DLX_Datapath/RegisterFile/N25920 ) );
  AOI22_X1 U81827 ( .A1(n105940), .A2(n81386), .B1(n105937), .B2(n110624), 
        .ZN(n95371) );
  OAI21_X1 U81828 ( .B1(n107392), .B2(n105943), .A(n95372), .ZN(
        \DLX_Datapath/RegisterFile/N25919 ) );
  AOI22_X1 U81829 ( .A1(n105940), .A2(n81320), .B1(n105937), .B2(n110413), 
        .ZN(n95372) );
  NOR2_X1 U81830 ( .A1(n95367), .A2(n105945), .ZN(n81706) );
  AOI21_X1 U81831 ( .B1(n105206), .B2(n95331), .A(n94663), .ZN(n95367) );
  NOR2_X1 U81832 ( .A1(n95331), .A2(n105945), .ZN(n81705) );
  OR2_X1 U81833 ( .A1(n94998), .A2(n94848), .ZN(n95331) );
  NAND2_X1 U81834 ( .A1(n95373), .A2(n94850), .ZN(n94998) );
  NOR2_X1 U81835 ( .A1(n94851), .A2(n107028), .ZN(n95373) );
  NAND2_X1 U81836 ( .A1(n105135), .A2(n94853), .ZN(n81703) );
  OAI21_X1 U81837 ( .B1(n107371), .B2(n105504), .A(n95375), .ZN(
        \DLX_Datapath/RegisterFile/N25898 ) );
  AOI22_X1 U81838 ( .A1(n104952), .A2(n94667), .B1(n105177), .B2(n70395), .ZN(
        n95375) );
  OAI21_X1 U81839 ( .B1(n107373), .B2(n105504), .A(n95377), .ZN(
        \DLX_Datapath/RegisterFile/N25897 ) );
  AOI22_X1 U81840 ( .A1(n104951), .A2(n94670), .B1(n106749), .B2(n70537), .ZN(
        n95377) );
  OAI21_X1 U81841 ( .B1(n106832), .B2(n105504), .A(n95378), .ZN(
        \DLX_Datapath/RegisterFile/N25896 ) );
  AOI22_X1 U81842 ( .A1(n104951), .A2(n94672), .B1(n105176), .B2(n69483), .ZN(
        n95378) );
  OAI21_X1 U81843 ( .B1(n107376), .B2(n105504), .A(n95379), .ZN(
        \DLX_Datapath/RegisterFile/N25895 ) );
  AOI22_X1 U81844 ( .A1(n104952), .A2(n94674), .B1(n106749), .B2(n70251), .ZN(
        n95379) );
  OAI21_X1 U81845 ( .B1(n107378), .B2(n105504), .A(n95380), .ZN(
        \DLX_Datapath/RegisterFile/N25894 ) );
  AOI22_X1 U81846 ( .A1(n104951), .A2(n94676), .B1(n104856), .B2(n74097), .ZN(
        n95380) );
  OAI21_X1 U81847 ( .B1(n107380), .B2(n105504), .A(n95381), .ZN(
        \DLX_Datapath/RegisterFile/N25893 ) );
  AOI22_X1 U81848 ( .A1(n104951), .A2(n94678), .B1(n106749), .B2(n70684), .ZN(
        n95381) );
  OAI21_X1 U81849 ( .B1(n107382), .B2(n105504), .A(n95382), .ZN(
        \DLX_Datapath/RegisterFile/N25892 ) );
  AOI22_X1 U81850 ( .A1(n104951), .A2(n94680), .B1(n106749), .B2(n74238), .ZN(
        n95382) );
  OAI21_X1 U81851 ( .B1(n107384), .B2(n105504), .A(n95383), .ZN(
        \DLX_Datapath/RegisterFile/N25891 ) );
  AOI22_X1 U81852 ( .A1(n104952), .A2(n94682), .B1(n106749), .B2(n74378), .ZN(
        n95383) );
  OAI21_X1 U81853 ( .B1(n107386), .B2(n105504), .A(n95384), .ZN(
        \DLX_Datapath/RegisterFile/N25890 ) );
  AOI22_X1 U81854 ( .A1(n104951), .A2(n94684), .B1(n104856), .B2(n73814), .ZN(
        n95384) );
  OAI21_X1 U81855 ( .B1(n107388), .B2(n105504), .A(n95385), .ZN(
        \DLX_Datapath/RegisterFile/N25889 ) );
  AOI22_X1 U81856 ( .A1(n104952), .A2(n94686), .B1(n104856), .B2(n73518), .ZN(
        n95385) );
  OAI21_X1 U81857 ( .B1(n107390), .B2(n105504), .A(n95386), .ZN(
        \DLX_Datapath/RegisterFile/N25888 ) );
  AOI22_X1 U81858 ( .A1(n95376), .A2(n94688), .B1(n105177), .B2(n73955), .ZN(
        n95386) );
  OAI21_X1 U81859 ( .B1(n107392), .B2(n105504), .A(n95387), .ZN(
        \DLX_Datapath/RegisterFile/N25887 ) );
  AOI22_X1 U81860 ( .A1(n104951), .A2(n94690), .B1(n105177), .B2(n73667), .ZN(
        n95387) );
  OAI21_X1 U81861 ( .B1(n107394), .B2(n105504), .A(n95388), .ZN(
        \DLX_Datapath/RegisterFile/N25886 ) );
  AOI22_X1 U81862 ( .A1(n104952), .A2(n94692), .B1(n105177), .B2(n73229), .ZN(
        n95388) );
  OAI21_X1 U81863 ( .B1(n107396), .B2(n105504), .A(n95389), .ZN(
        \DLX_Datapath/RegisterFile/N25885 ) );
  AOI22_X1 U81864 ( .A1(n104952), .A2(n94694), .B1(n105177), .B2(n73371), .ZN(
        n95389) );
  OAI21_X1 U81865 ( .B1(n107398), .B2(n105504), .A(n95390), .ZN(
        \DLX_Datapath/RegisterFile/N25884 ) );
  AOI22_X1 U81866 ( .A1(n95376), .A2(n94696), .B1(n105177), .B2(n73087), .ZN(
        n95390) );
  OAI21_X1 U81867 ( .B1(n107400), .B2(n105504), .A(n95391), .ZN(
        \DLX_Datapath/RegisterFile/N25883 ) );
  AOI22_X1 U81868 ( .A1(n95376), .A2(n94698), .B1(n105177), .B2(n72937), .ZN(
        n95391) );
  OAI21_X1 U81869 ( .B1(n107402), .B2(n105504), .A(n95392), .ZN(
        \DLX_Datapath/RegisterFile/N25882 ) );
  AOI22_X1 U81870 ( .A1(n104951), .A2(n94700), .B1(n105177), .B2(n70833), .ZN(
        n95392) );
  OAI21_X1 U81871 ( .B1(n107404), .B2(n105504), .A(n95393), .ZN(
        \DLX_Datapath/RegisterFile/N25881 ) );
  AOI22_X1 U81872 ( .A1(n104952), .A2(n94702), .B1(n104856), .B2(n70992), .ZN(
        n95393) );
  OAI21_X1 U81873 ( .B1(n107406), .B2(n105504), .A(n95394), .ZN(
        \DLX_Datapath/RegisterFile/N25880 ) );
  AOI22_X1 U81874 ( .A1(n104951), .A2(n94704), .B1(n105176), .B2(n71137), .ZN(
        n95394) );
  OAI21_X1 U81875 ( .B1(n107408), .B2(n105504), .A(n95395), .ZN(
        \DLX_Datapath/RegisterFile/N25879 ) );
  AOI22_X1 U81876 ( .A1(n95376), .A2(n94706), .B1(n106749), .B2(n70098), .ZN(
        n95395) );
  OAI21_X1 U81877 ( .B1(n107410), .B2(n105504), .A(n95396), .ZN(
        \DLX_Datapath/RegisterFile/N25878 ) );
  AOI22_X1 U81878 ( .A1(n104951), .A2(n94708), .B1(n105177), .B2(n72627), .ZN(
        n95396) );
  OAI21_X1 U81879 ( .B1(n107412), .B2(n105504), .A(n95397), .ZN(
        \DLX_Datapath/RegisterFile/N25877 ) );
  AOI22_X1 U81880 ( .A1(n95376), .A2(n94710), .B1(n106749), .B2(n71286), .ZN(
        n95397) );
  OAI21_X1 U81881 ( .B1(n107367), .B2(n105504), .A(n95398), .ZN(
        \DLX_Datapath/RegisterFile/N25876 ) );
  AOI22_X1 U81882 ( .A1(n104952), .A2(n94712), .B1(n105177), .B2(n72769), .ZN(
        n95398) );
  OAI21_X1 U81883 ( .B1(n107369), .B2(n105504), .A(n95399), .ZN(
        \DLX_Datapath/RegisterFile/N25875 ) );
  AOI22_X1 U81884 ( .A1(n104951), .A2(n94714), .B1(n106749), .B2(n72479), .ZN(
        n95399) );
  OAI21_X1 U81885 ( .B1(n108974), .B2(n105504), .A(n95400), .ZN(
        \DLX_Datapath/RegisterFile/N25874 ) );
  AOI22_X1 U81886 ( .A1(n104952), .A2(n81259), .B1(n105176), .B2(n71879), .ZN(
        n95400) );
  OAI21_X1 U81887 ( .B1(n111063), .B2(n105504), .A(n95401), .ZN(
        \DLX_Datapath/RegisterFile/N25873 ) );
  AOI22_X1 U81888 ( .A1(n95376), .A2(n94717), .B1(n105176), .B2(n72328), .ZN(
        n95401) );
  OAI21_X1 U81889 ( .B1(n111062), .B2(n105504), .A(n95402), .ZN(
        \DLX_Datapath/RegisterFile/N25872 ) );
  AOI22_X1 U81890 ( .A1(n95376), .A2(n94719), .B1(n105177), .B2(n72177), .ZN(
        n95402) );
  OAI21_X1 U81891 ( .B1(n111061), .B2(n105504), .A(n95403), .ZN(
        \DLX_Datapath/RegisterFile/N25871 ) );
  AOI22_X1 U81892 ( .A1(n104951), .A2(n94721), .B1(n106749), .B2(n72033), .ZN(
        n95403) );
  OAI21_X1 U81893 ( .B1(n111060), .B2(n105504), .A(n95404), .ZN(
        \DLX_Datapath/RegisterFile/N25870 ) );
  AOI22_X1 U81894 ( .A1(n104951), .A2(n94723), .B1(n106749), .B2(n71435), .ZN(
        n95404) );
  OAI21_X1 U81895 ( .B1(n111059), .B2(n105504), .A(n95405), .ZN(
        \DLX_Datapath/RegisterFile/N25869 ) );
  AOI22_X1 U81896 ( .A1(n104952), .A2(n94725), .B1(n106749), .B2(n71730), .ZN(
        n95405) );
  OAI21_X1 U81897 ( .B1(n111058), .B2(n105504), .A(n95406), .ZN(
        \DLX_Datapath/RegisterFile/N25868 ) );
  AOI22_X1 U81898 ( .A1(n104951), .A2(n94727), .B1(n104856), .B2(n71586), .ZN(
        n95406) );
  OAI21_X1 U81899 ( .B1(n111057), .B2(n105504), .A(n95407), .ZN(
        \DLX_Datapath/RegisterFile/N25867 ) );
  AOI22_X1 U81900 ( .A1(n104952), .A2(n94729), .B1(n105176), .B2(n69484), .ZN(
        n95407) );
  OAI21_X1 U81901 ( .B1(n95409), .B2(n94663), .A(n95374), .ZN(n95408) );
  AOI21_X1 U81902 ( .B1(n95036), .B2(n111024), .A(n94366), .ZN(n95409) );
  NOR2_X1 U81903 ( .A1(n95410), .A2(n106748), .ZN(n95376) );
  NOR2_X1 U81904 ( .A1(n95411), .A2(n106753), .ZN(n95036) );
  NAND2_X1 U81905 ( .A1(n95374), .A2(n111024), .ZN(n95410) );
  NAND2_X1 U81906 ( .A1(n105135), .A2(n94892), .ZN(n95374) );
  OAI21_X1 U81908 ( .B1(n106146), .B2(n105503), .A(n95414), .ZN(
        \DLX_Datapath/RegisterFile/N25866 ) );
  AOI22_X1 U81909 ( .A1(n104980), .A2(n70291), .B1(n104926), .B2(n81360), .ZN(
        n95414) );
  OAI21_X1 U81910 ( .B1(n105968), .B2(n105503), .A(n95417), .ZN(
        \DLX_Datapath/RegisterFile/N25865 ) );
  AOI22_X1 U81911 ( .A1(n104981), .A2(n70433), .B1(n104927), .B2(n94511), .ZN(
        n95417) );
  OAI21_X1 U81912 ( .B1(n106135), .B2(n105503), .A(n95418), .ZN(
        \DLX_Datapath/RegisterFile/N25864 ) );
  AOI22_X1 U81913 ( .A1(n104980), .A2(n69486), .B1(n104926), .B2(n81539), .ZN(
        n95418) );
  OAI21_X1 U81914 ( .B1(n106209), .B2(n105503), .A(n95419), .ZN(
        \DLX_Datapath/RegisterFile/N25863 ) );
  AOI22_X1 U81915 ( .A1(n104981), .A2(n70147), .B1(n104927), .B2(n81301), .ZN(
        n95419) );
  OAI21_X1 U81916 ( .B1(n81306), .B2(n105503), .A(n95420), .ZN(
        \DLX_Datapath/RegisterFile/N25862 ) );
  AOI22_X1 U81917 ( .A1(n104982), .A2(n73993), .B1(n104928), .B2(n81308), .ZN(
        n95420) );
  OAI21_X1 U81918 ( .B1(n81408), .B2(n105503), .A(n95421), .ZN(
        \DLX_Datapath/RegisterFile/N25861 ) );
  AOI22_X1 U81919 ( .A1(n104981), .A2(n70580), .B1(n104927), .B2(n94516), .ZN(
        n95421) );
  OAI21_X1 U81920 ( .B1(n106254), .B2(n105503), .A(n95422), .ZN(
        \DLX_Datapath/RegisterFile/N25860 ) );
  AOI22_X1 U81921 ( .A1(n104980), .A2(n74134), .B1(n104926), .B2(n81272), .ZN(
        n95422) );
  OAI21_X1 U81922 ( .B1(n105990), .B2(n105503), .A(n95423), .ZN(
        \DLX_Datapath/RegisterFile/N25859 ) );
  AOI22_X1 U81923 ( .A1(n104982), .A2(n74274), .B1(n104928), .B2(n94519), .ZN(
        n95423) );
  OAI21_X1 U81924 ( .B1(n106332), .B2(n105503), .A(n95424), .ZN(
        \DLX_Datapath/RegisterFile/N25858 ) );
  AOI22_X1 U81925 ( .A1(n104982), .A2(n73710), .B1(n104928), .B2(n80192), .ZN(
        n95424) );
  OAI21_X1 U81926 ( .B1(n81315), .B2(n105503), .A(n95425), .ZN(
        \DLX_Datapath/RegisterFile/N25857 ) );
  AOI22_X1 U81927 ( .A1(n104980), .A2(n73414), .B1(n104926), .B2(n81474), .ZN(
        n95425) );
  OAI21_X1 U81928 ( .B1(n106131), .B2(n105503), .A(n95426), .ZN(
        \DLX_Datapath/RegisterFile/N25856 ) );
  AOI22_X1 U81929 ( .A1(n104981), .A2(n73851), .B1(n104927), .B2(n94523), .ZN(
        n95426) );
  OAI21_X1 U81930 ( .B1(n81318), .B2(n105503), .A(n95427), .ZN(
        \DLX_Datapath/RegisterFile/N25855 ) );
  AOI22_X1 U81931 ( .A1(n104982), .A2(n73563), .B1(n104928), .B2(n106061), 
        .ZN(n95427) );
  OAI21_X1 U81932 ( .B1(n106164), .B2(n105503), .A(n95428), .ZN(
        \DLX_Datapath/RegisterFile/N25854 ) );
  AOI22_X1 U81933 ( .A1(n104982), .A2(n73125), .B1(n104927), .B2(n81347), .ZN(
        n95428) );
  OAI21_X1 U81934 ( .B1(n106104), .B2(n105503), .A(n95429), .ZN(
        \DLX_Datapath/RegisterFile/N25853 ) );
  AOI22_X1 U81935 ( .A1(n104980), .A2(n73267), .B1(n104928), .B2(n94527), .ZN(
        n95429) );
  OAI21_X1 U81936 ( .B1(n81294), .B2(n105503), .A(n95430), .ZN(
        \DLX_Datapath/RegisterFile/N25852 ) );
  AOI22_X1 U81937 ( .A1(n104980), .A2(n72983), .B1(n104926), .B2(n81297), .ZN(
        n95430) );
  OAI21_X1 U81938 ( .B1(n106108), .B2(n105503), .A(n95431), .ZN(
        \DLX_Datapath/RegisterFile/N25851 ) );
  AOI22_X1 U81939 ( .A1(n104981), .A2(n72833), .B1(n104926), .B2(n94530), .ZN(
        n95431) );
  OAI21_X1 U81940 ( .B1(n106230), .B2(n105503), .A(n95432), .ZN(
        \DLX_Datapath/RegisterFile/N25850 ) );
  AOI22_X1 U81941 ( .A1(n104982), .A2(n70729), .B1(n104928), .B2(n81286), .ZN(
        n95432) );
  OAI21_X1 U81942 ( .B1(n106171), .B2(n105503), .A(n95433), .ZN(
        \DLX_Datapath/RegisterFile/N25849 ) );
  AOI22_X1 U81943 ( .A1(n104981), .A2(n70888), .B1(n104928), .B2(n106169), 
        .ZN(n95433) );
  OAI21_X1 U81944 ( .B1(n81281), .B2(n105503), .A(n95434), .ZN(
        \DLX_Datapath/RegisterFile/N25848 ) );
  AOI22_X1 U81945 ( .A1(n104980), .A2(n71033), .B1(n104927), .B2(n81283), .ZN(
        n95434) );
  OAI21_X1 U81946 ( .B1(n106069), .B2(n105503), .A(n95435), .ZN(
        \DLX_Datapath/RegisterFile/N25847 ) );
  AOI22_X1 U81947 ( .A1(n104981), .A2(n69994), .B1(n104926), .B2(n81453), .ZN(
        n95435) );
  OAI21_X1 U81948 ( .B1(n81310), .B2(n105503), .A(n95436), .ZN(
        \DLX_Datapath/RegisterFile/N25846 ) );
  AOI22_X1 U81949 ( .A1(n104982), .A2(n72523), .B1(n104927), .B2(n94536), .ZN(
        n95436) );
  OAI21_X1 U81950 ( .B1(n106244), .B2(n95413), .A(n95437), .ZN(
        \DLX_Datapath/RegisterFile/N25845 ) );
  AOI22_X1 U81951 ( .A1(n104981), .A2(n71182), .B1(n104928), .B2(n106241), 
        .ZN(n95437) );
  OAI21_X1 U81952 ( .B1(n106157), .B2(n95413), .A(n95438), .ZN(
        \DLX_Datapath/RegisterFile/N25844 ) );
  AOI22_X1 U81953 ( .A1(n104982), .A2(n72665), .B1(n104927), .B2(n81351), .ZN(
        n95438) );
  OAI21_X1 U81954 ( .B1(n106114), .B2(n95413), .A(n95439), .ZN(
        \DLX_Datapath/RegisterFile/N25843 ) );
  AOI22_X1 U81955 ( .A1(n104982), .A2(n72375), .B1(n104926), .B2(n106020), 
        .ZN(n95439) );
  OAI21_X1 U81956 ( .B1(n81588), .B2(n105503), .A(n95440), .ZN(
        \DLX_Datapath/RegisterFile/N25842 ) );
  AOI22_X1 U81957 ( .A1(n104980), .A2(n71775), .B1(n104926), .B2(n94541), .ZN(
        n95440) );
  OAI21_X1 U81958 ( .B1(n106259), .B2(n95413), .A(n95441), .ZN(
        \DLX_Datapath/RegisterFile/N25841 ) );
  AOI22_X1 U81959 ( .A1(n104980), .A2(n72224), .B1(n104927), .B2(n81269), .ZN(
        n95441) );
  OAI21_X1 U81960 ( .B1(n106046), .B2(n95413), .A(n95442), .ZN(
        \DLX_Datapath/RegisterFile/N25840 ) );
  AOI22_X1 U81961 ( .A1(n104981), .A2(n72073), .B1(n104926), .B2(n105624), 
        .ZN(n95442) );
  OAI21_X1 U81962 ( .B1(n106048), .B2(n95413), .A(n95443), .ZN(
        \DLX_Datapath/RegisterFile/N25839 ) );
  AOI22_X1 U81963 ( .A1(n104982), .A2(n71929), .B1(n104927), .B2(n94546), .ZN(
        n95443) );
  OAI21_X1 U81964 ( .B1(n106096), .B2(n95413), .A(n95444), .ZN(
        \DLX_Datapath/RegisterFile/N25838 ) );
  AOI22_X1 U81965 ( .A1(n104981), .A2(n71331), .B1(n104927), .B2(n94548), .ZN(
        n95444) );
  OAI21_X1 U81966 ( .B1(n81498), .B2(n105503), .A(n95445), .ZN(
        \DLX_Datapath/RegisterFile/N25837 ) );
  AOI22_X1 U81967 ( .A1(n104980), .A2(n71626), .B1(n104928), .B2(n81783), .ZN(
        n95445) );
  OAI21_X1 U81968 ( .B1(n105220), .B2(n95413), .A(n95446), .ZN(
        \DLX_Datapath/RegisterFile/N25836 ) );
  AOI22_X1 U81969 ( .A1(n104980), .A2(n71482), .B1(n104928), .B2(n80188), .ZN(
        n95446) );
  OAI21_X1 U81970 ( .B1(n106266), .B2(n95413), .A(n95447), .ZN(
        \DLX_Datapath/RegisterFile/N25835 ) );
  AOI22_X1 U81971 ( .A1(n104981), .A2(n69591), .B1(n104926), .B2(n81265), .ZN(
        n95447) );
  AOI21_X1 U81973 ( .B1(n95450), .B2(n94258), .A(n95449), .ZN(n95415) );
  NOR2_X1 U81974 ( .A1(n95413), .A2(n105091), .ZN(n95449) );
  NAND2_X1 U81975 ( .A1(n105134), .A2(n94934), .ZN(n95413) );
  OAI21_X1 U81976 ( .B1(n106146), .B2(n105499), .A(n95454), .ZN(
        \DLX_Datapath/RegisterFile/N25834 ) );
  AOI22_X1 U81977 ( .A1(n105498), .A2(n94559), .B1(n104977), .B2(n107855), 
        .ZN(n95454) );
  OAI21_X1 U81978 ( .B1(n105969), .B2(n105499), .A(n95457), .ZN(
        \DLX_Datapath/RegisterFile/N25833 ) );
  AOI22_X1 U81979 ( .A1(n105497), .A2(n94562), .B1(n104978), .B2(n107952), 
        .ZN(n95457) );
  OAI21_X1 U81980 ( .B1(n81378), .B2(n105499), .A(n95458), .ZN(
        \DLX_Datapath/RegisterFile/N25832 ) );
  AOI22_X1 U81981 ( .A1(n105498), .A2(n94564), .B1(n104977), .B2(n107214), 
        .ZN(n95458) );
  OAI21_X1 U81982 ( .B1(n106211), .B2(n105499), .A(n95459), .ZN(
        \DLX_Datapath/RegisterFile/N25831 ) );
  AOI22_X1 U81983 ( .A1(n105497), .A2(n94566), .B1(n104979), .B2(n107752), 
        .ZN(n95459) );
  OAI21_X1 U81984 ( .B1(n81306), .B2(n105499), .A(n95460), .ZN(
        \DLX_Datapath/RegisterFile/N25830 ) );
  AOI22_X1 U81985 ( .A1(n105498), .A2(n94568), .B1(n104977), .B2(n110655), 
        .ZN(n95460) );
  OAI21_X1 U81986 ( .B1(n81408), .B2(n105499), .A(n95461), .ZN(
        \DLX_Datapath/RegisterFile/N25829 ) );
  AOI22_X1 U81987 ( .A1(n105497), .A2(n94570), .B1(n104978), .B2(n108054), 
        .ZN(n95461) );
  OAI21_X1 U81988 ( .B1(n106254), .B2(n105499), .A(n95462), .ZN(
        \DLX_Datapath/RegisterFile/N25828 ) );
  AOI22_X1 U81989 ( .A1(n105498), .A2(n94572), .B1(n104978), .B2(n110752), 
        .ZN(n95462) );
  OAI21_X1 U81990 ( .B1(n105990), .B2(n105499), .A(n95463), .ZN(
        \DLX_Datapath/RegisterFile/N25827 ) );
  AOI22_X1 U81991 ( .A1(n105497), .A2(n94574), .B1(n104979), .B2(n110853), 
        .ZN(n95463) );
  OAI21_X1 U81992 ( .B1(n106332), .B2(n105499), .A(n95464), .ZN(
        \DLX_Datapath/RegisterFile/N25826 ) );
  AOI22_X1 U81993 ( .A1(n105497), .A2(n94576), .B1(n104979), .B2(n110448), 
        .ZN(n95464) );
  OAI21_X1 U81994 ( .B1(n81315), .B2(n105499), .A(n95465), .ZN(
        \DLX_Datapath/RegisterFile/N25825 ) );
  AOI22_X1 U81995 ( .A1(n105496), .A2(n94578), .B1(n104977), .B2(n110231), 
        .ZN(n95465) );
  OAI21_X1 U81996 ( .B1(n106131), .B2(n105499), .A(n95466), .ZN(
        \DLX_Datapath/RegisterFile/N25824 ) );
  AOI22_X1 U81997 ( .A1(n105496), .A2(n94580), .B1(n104978), .B2(n110548), 
        .ZN(n95466) );
  OAI21_X1 U81998 ( .B1(n106185), .B2(n105499), .A(n95467), .ZN(
        \DLX_Datapath/RegisterFile/N25823 ) );
  AOI22_X1 U81999 ( .A1(n105496), .A2(n94582), .B1(n104979), .B2(n110339), 
        .ZN(n95467) );
  OAI21_X1 U82000 ( .B1(n106165), .B2(n105499), .A(n95468), .ZN(
        \DLX_Datapath/RegisterFile/N25822 ) );
  AOI22_X1 U82001 ( .A1(n105496), .A2(n94584), .B1(n104979), .B2(n110013), 
        .ZN(n95468) );
  OAI21_X1 U82002 ( .B1(n106103), .B2(n105499), .A(n95469), .ZN(
        \DLX_Datapath/RegisterFile/N25821 ) );
  AOI22_X1 U82003 ( .A1(n105496), .A2(n94586), .B1(n104977), .B2(n110121), 
        .ZN(n95469) );
  OAI21_X1 U82004 ( .B1(n81294), .B2(n105499), .A(n95470), .ZN(
        \DLX_Datapath/RegisterFile/N25820 ) );
  AOI22_X1 U82005 ( .A1(n105496), .A2(n94588), .B1(n104977), .B2(n109904), 
        .ZN(n95470) );
  OAI21_X1 U82006 ( .B1(n106111), .B2(n105499), .A(n95471), .ZN(
        \DLX_Datapath/RegisterFile/N25819 ) );
  AOI22_X1 U82007 ( .A1(n105496), .A2(n94590), .B1(n104978), .B2(n109786), 
        .ZN(n95471) );
  OAI21_X1 U82008 ( .B1(n106230), .B2(n105499), .A(n95472), .ZN(
        \DLX_Datapath/RegisterFile/N25818 ) );
  AOI22_X1 U82009 ( .A1(n105496), .A2(n94592), .B1(n104979), .B2(n108160), 
        .ZN(n95472) );
  OAI21_X1 U82010 ( .B1(n106170), .B2(n105499), .A(n95473), .ZN(
        \DLX_Datapath/RegisterFile/N25817 ) );
  AOI22_X1 U82011 ( .A1(n105496), .A2(n94594), .B1(n104978), .B2(n108283), 
        .ZN(n95473) );
  OAI21_X1 U82012 ( .B1(n106236), .B2(n105499), .A(n95474), .ZN(
        \DLX_Datapath/RegisterFile/N25816 ) );
  AOI22_X1 U82013 ( .A1(n105496), .A2(n94596), .B1(n104977), .B2(n108394), 
        .ZN(n95474) );
  OAI21_X1 U82014 ( .B1(n106071), .B2(n105499), .A(n95475), .ZN(
        \DLX_Datapath/RegisterFile/N25815 ) );
  AOI22_X1 U82015 ( .A1(n105496), .A2(n94598), .B1(n104978), .B2(n107632), 
        .ZN(n95475) );
  OAI21_X1 U82016 ( .B1(n81310), .B2(n105499), .A(n95476), .ZN(
        \DLX_Datapath/RegisterFile/N25814 ) );
  AOI22_X1 U82017 ( .A1(n105497), .A2(n94600), .B1(n104979), .B2(n109550), 
        .ZN(n95476) );
  OAI21_X1 U82018 ( .B1(n106244), .B2(n95453), .A(n95477), .ZN(
        \DLX_Datapath/RegisterFile/N25813 ) );
  AOI22_X1 U82019 ( .A1(n105497), .A2(n94602), .B1(n104978), .B2(n108511), 
        .ZN(n95477) );
  OAI21_X1 U82020 ( .B1(n106157), .B2(n95453), .A(n95478), .ZN(
        \DLX_Datapath/RegisterFile/N25812 ) );
  AOI22_X1 U82021 ( .A1(n105498), .A2(n94604), .B1(n104979), .B2(n109655), 
        .ZN(n95478) );
  OAI21_X1 U82022 ( .B1(n106113), .B2(n95453), .A(n95479), .ZN(
        \DLX_Datapath/RegisterFile/N25811 ) );
  AOI22_X1 U82023 ( .A1(n105497), .A2(n94606), .B1(n104979), .B2(n109439), 
        .ZN(n95479) );
  OAI21_X1 U82024 ( .B1(n81588), .B2(n105499), .A(n95480), .ZN(
        \DLX_Datapath/RegisterFile/N25810 ) );
  AOI22_X1 U82025 ( .A1(n105498), .A2(n94608), .B1(n104978), .B2(n108976), 
        .ZN(n95480) );
  OAI21_X1 U82026 ( .B1(n106259), .B2(n95453), .A(n95481), .ZN(
        \DLX_Datapath/RegisterFile/N25809 ) );
  AOI22_X1 U82027 ( .A1(n105498), .A2(n94610), .B1(n104977), .B2(n109324), 
        .ZN(n95481) );
  OAI21_X1 U82028 ( .B1(n106045), .B2(n95453), .A(n95482), .ZN(
        \DLX_Datapath/RegisterFile/N25808 ) );
  AOI22_X1 U82029 ( .A1(n105497), .A2(n94612), .B1(n104977), .B2(n109206), 
        .ZN(n95482) );
  OAI21_X1 U82030 ( .B1(n106050), .B2(n95453), .A(n95483), .ZN(
        \DLX_Datapath/RegisterFile/N25807 ) );
  AOI22_X1 U82031 ( .A1(n105498), .A2(n94614), .B1(n104978), .B2(n109098), 
        .ZN(n95483) );
  OAI21_X1 U82032 ( .B1(n106094), .B2(n95453), .A(n95484), .ZN(
        \DLX_Datapath/RegisterFile/N25806 ) );
  AOI22_X1 U82033 ( .A1(n105497), .A2(n94616), .B1(n104978), .B2(n108633), 
        .ZN(n95484) );
  OAI21_X1 U82034 ( .B1(n81498), .B2(n105499), .A(n95485), .ZN(
        \DLX_Datapath/RegisterFile/N25805 ) );
  AOI22_X1 U82035 ( .A1(n105498), .A2(n94618), .B1(n104979), .B2(n108860), 
        .ZN(n95485) );
  OAI21_X1 U82036 ( .B1(n105218), .B2(n95453), .A(n95486), .ZN(
        \DLX_Datapath/RegisterFile/N25804 ) );
  AOI22_X1 U82037 ( .A1(n105498), .A2(n94620), .B1(n104977), .B2(n108748), 
        .ZN(n95486) );
  OAI21_X1 U82038 ( .B1(n106266), .B2(n95453), .A(n95487), .ZN(
        \DLX_Datapath/RegisterFile/N25803 ) );
  AOI22_X1 U82039 ( .A1(n105497), .A2(n94622), .B1(n104977), .B2(n107288), 
        .ZN(n95487) );
  NOR2_X1 U82041 ( .A1(n95448), .A2(n95489), .ZN(n95455) );
  NOR2_X1 U82042 ( .A1(n95453), .A2(n105089), .ZN(n95489) );
  NAND2_X1 U82043 ( .A1(n94296), .A2(n105134), .ZN(n95453) );
  OAI21_X1 U82044 ( .B1(n106146), .B2(n81647), .A(n95490), .ZN(
        \DLX_Datapath/RegisterFile/N25802 ) );
  AOI22_X1 U82045 ( .A1(n104930), .A2(n107856), .B1(n105975), .B2(n81521), 
        .ZN(n95490) );
  OAI21_X1 U82046 ( .B1(n106136), .B2(n81647), .A(n95491), .ZN(
        \DLX_Datapath/RegisterFile/N25800 ) );
  AOI22_X1 U82047 ( .A1(n104931), .A2(n107215), .B1(n105974), .B2(n81380), 
        .ZN(n95491) );
  OAI21_X1 U82048 ( .B1(n106208), .B2(n81647), .A(n95492), .ZN(
        \DLX_Datapath/RegisterFile/N25799 ) );
  AOI22_X1 U82049 ( .A1(n104930), .A2(n107753), .B1(n105975), .B2(n81377), 
        .ZN(n95492) );
  OAI21_X1 U82050 ( .B1(n81306), .B2(n105976), .A(n95493), .ZN(
        \DLX_Datapath/RegisterFile/N25798 ) );
  AOI22_X1 U82051 ( .A1(n104931), .A2(n110656), .B1(n105975), .B2(n81428), 
        .ZN(n95493) );
  OAI21_X1 U82052 ( .B1(n81408), .B2(n81647), .A(n95494), .ZN(
        \DLX_Datapath/RegisterFile/N25797 ) );
  AOI22_X1 U82053 ( .A1(n104929), .A2(n108055), .B1(n105974), .B2(n81410), 
        .ZN(n95494) );
  OAI21_X1 U82054 ( .B1(n106254), .B2(n105976), .A(n95495), .ZN(
        \DLX_Datapath/RegisterFile/N25796 ) );
  AOI22_X1 U82055 ( .A1(n104929), .A2(n110753), .B1(n81700), .B2(n105973), 
        .ZN(n95495) );
  OAI21_X1 U82056 ( .B1(n81629), .B2(n105976), .A(n95496), .ZN(
        \DLX_Datapath/RegisterFile/N25795 ) );
  AOI22_X1 U82057 ( .A1(n104930), .A2(n110854), .B1(n105974), .B2(n81632), 
        .ZN(n95496) );
  OAI21_X1 U82058 ( .B1(n106330), .B2(n105976), .A(n95497), .ZN(
        \DLX_Datapath/RegisterFile/N25794 ) );
  AOI22_X1 U82059 ( .A1(n104931), .A2(n110449), .B1(n105975), .B2(n81414), 
        .ZN(n95497) );
  OAI21_X1 U82060 ( .B1(n81315), .B2(n105976), .A(n95498), .ZN(
        \DLX_Datapath/RegisterFile/N25793 ) );
  AOI22_X1 U82061 ( .A1(n104931), .A2(n111020), .B1(n105973), .B2(n81317), 
        .ZN(n95498) );
  OAI21_X1 U82062 ( .B1(n106128), .B2(n105976), .A(n95499), .ZN(
        \DLX_Datapath/RegisterFile/N25792 ) );
  AOI22_X1 U82063 ( .A1(n104929), .A2(n111018), .B1(n105973), .B2(n81386), 
        .ZN(n95499) );
  OAI21_X1 U82064 ( .B1(n106185), .B2(n105976), .A(n95500), .ZN(
        \DLX_Datapath/RegisterFile/N25791 ) );
  AOI22_X1 U82065 ( .A1(n104929), .A2(n111019), .B1(n105973), .B2(n81320), 
        .ZN(n95500) );
  OAI21_X1 U82066 ( .B1(n106164), .B2(n105976), .A(n95501), .ZN(
        \DLX_Datapath/RegisterFile/N25790 ) );
  AOI22_X1 U82067 ( .A1(n104930), .A2(n110014), .B1(n105973), .B2(n81604), 
        .ZN(n95501) );
  OAI21_X1 U82068 ( .B1(n106106), .B2(n105976), .A(n95502), .ZN(
        \DLX_Datapath/RegisterFile/N25789 ) );
  AOI22_X1 U82069 ( .A1(n104931), .A2(n111021), .B1(n105973), .B2(n81405), 
        .ZN(n95502) );
  OAI21_X1 U82070 ( .B1(n81294), .B2(n105976), .A(n95503), .ZN(
        \DLX_Datapath/RegisterFile/N25788 ) );
  AOI22_X1 U82071 ( .A1(n104930), .A2(n109905), .B1(n105973), .B2(n81402), 
        .ZN(n95503) );
  OAI21_X1 U82072 ( .B1(n106109), .B2(n105976), .A(n95504), .ZN(
        \DLX_Datapath/RegisterFile/N25787 ) );
  AOI22_X1 U82073 ( .A1(n104929), .A2(n109787), .B1(n105973), .B2(n81400), 
        .ZN(n95504) );
  OAI21_X1 U82074 ( .B1(n106170), .B2(n105976), .A(n95505), .ZN(
        \DLX_Datapath/RegisterFile/N25785 ) );
  AOI22_X1 U82075 ( .A1(n104930), .A2(n108284), .B1(n105973), .B2(n81373), 
        .ZN(n95505) );
  OAI21_X1 U82076 ( .B1(n81281), .B2(n105976), .A(n95506), .ZN(
        \DLX_Datapath/RegisterFile/N25784 ) );
  AOI22_X1 U82077 ( .A1(n104931), .A2(n108395), .B1(n105975), .B2(n81322), 
        .ZN(n95506) );
  OAI21_X1 U82078 ( .B1(n106072), .B2(n105976), .A(n95507), .ZN(
        \DLX_Datapath/RegisterFile/N25783 ) );
  AOI22_X1 U82079 ( .A1(n104930), .A2(n107633), .B1(n105974), .B2(n81506), 
        .ZN(n95507) );
  OAI21_X1 U82080 ( .B1(n81310), .B2(n105976), .A(n95508), .ZN(
        \DLX_Datapath/RegisterFile/N25782 ) );
  AOI22_X1 U82081 ( .A1(n104931), .A2(n109551), .B1(n105975), .B2(n81313), 
        .ZN(n95508) );
  OAI21_X1 U82082 ( .B1(n106159), .B2(n105976), .A(n95509), .ZN(
        \DLX_Datapath/RegisterFile/N25780 ) );
  AOI22_X1 U82083 ( .A1(n104929), .A2(n109656), .B1(n105974), .B2(n81425), 
        .ZN(n95509) );
  OAI21_X1 U82084 ( .B1(n106115), .B2(n105976), .A(n95510), .ZN(
        \DLX_Datapath/RegisterFile/N25779 ) );
  AOI22_X1 U82085 ( .A1(n104929), .A2(n109440), .B1(n105975), .B2(n81396), 
        .ZN(n95510) );
  OAI21_X1 U82086 ( .B1(n81588), .B2(n105976), .A(n95511), .ZN(
        \DLX_Datapath/RegisterFile/N25778 ) );
  AOI22_X1 U82087 ( .A1(n104930), .A2(n108977), .B1(n105974), .B2(n81590), 
        .ZN(n95511) );
  OAI21_X1 U82088 ( .B1(n106259), .B2(n105976), .A(n95512), .ZN(
        \DLX_Datapath/RegisterFile/N25777 ) );
  AOI22_X1 U82089 ( .A1(n104930), .A2(n109325), .B1(n105975), .B2(n81423), 
        .ZN(n95512) );
  OAI21_X1 U82090 ( .B1(n106044), .B2(n105976), .A(n95513), .ZN(
        \DLX_Datapath/RegisterFile/N25776 ) );
  AOI22_X1 U82091 ( .A1(n104931), .A2(n109207), .B1(n105974), .B2(n81511), 
        .ZN(n95513) );
  OAI21_X1 U82092 ( .B1(n106051), .B2(n105976), .A(n95514), .ZN(
        \DLX_Datapath/RegisterFile/N25775 ) );
  AOI22_X1 U82093 ( .A1(n104929), .A2(n109099), .B1(n105975), .B2(n81503), 
        .ZN(n95514) );
  OAI21_X1 U82094 ( .B1(n106266), .B2(n81647), .A(n95515), .ZN(
        \DLX_Datapath/RegisterFile/N25771 ) );
  AOI22_X1 U82095 ( .A1(n104931), .A2(n107289), .B1(n105974), .B2(n81327), 
        .ZN(n95515) );
  NOR2_X1 U82097 ( .A1(n95488), .A2(n95516), .ZN(n81649) );
  NOR2_X1 U82098 ( .A1(n81647), .A2(n105089), .ZN(n95516) );
  AOI21_X1 U82099 ( .B1(n105205), .B2(n95448), .A(n94663), .ZN(n95488) );
  OR2_X1 U82100 ( .A1(n95517), .A2(n94999), .ZN(n95448) );
  NAND2_X1 U82101 ( .A1(n105133), .A2(n94331), .ZN(n81647) );
  OAI21_X1 U82102 ( .B1(n106146), .B2(n105495), .A(n95519), .ZN(
        \DLX_Datapath/RegisterFile/N25770 ) );
  AOI22_X1 U82103 ( .A1(n104844), .A2(n94667), .B1(n105494), .B2(n107857), 
        .ZN(n95519) );
  OAI21_X1 U82104 ( .B1(n105968), .B2(n105495), .A(n95522), .ZN(
        \DLX_Datapath/RegisterFile/N25769 ) );
  AOI22_X1 U82105 ( .A1(n104844), .A2(n94670), .B1(n105493), .B2(n107954), 
        .ZN(n95522) );
  OAI21_X1 U82106 ( .B1(n106138), .B2(n105495), .A(n95523), .ZN(
        \DLX_Datapath/RegisterFile/N25768 ) );
  AOI22_X1 U82107 ( .A1(n104844), .A2(n94672), .B1(n95521), .B2(n107216), .ZN(
        n95523) );
  OAI21_X1 U82108 ( .B1(n81299), .B2(n105495), .A(n95524), .ZN(
        \DLX_Datapath/RegisterFile/N25767 ) );
  AOI22_X1 U82109 ( .A1(n104844), .A2(n94674), .B1(n95521), .B2(n107754), .ZN(
        n95524) );
  OAI21_X1 U82110 ( .B1(n81306), .B2(n105495), .A(n95525), .ZN(
        \DLX_Datapath/RegisterFile/N25766 ) );
  AOI22_X1 U82111 ( .A1(n104845), .A2(n94676), .B1(n95521), .B2(n110657), .ZN(
        n95525) );
  OAI21_X1 U82112 ( .B1(n81408), .B2(n105495), .A(n95526), .ZN(
        \DLX_Datapath/RegisterFile/N25765 ) );
  AOI22_X1 U82113 ( .A1(n104846), .A2(n94678), .B1(n95521), .B2(n108056), .ZN(
        n95526) );
  OAI21_X1 U82114 ( .B1(n106254), .B2(n105495), .A(n95527), .ZN(
        \DLX_Datapath/RegisterFile/N25764 ) );
  AOI22_X1 U82115 ( .A1(n104845), .A2(n94680), .B1(n95521), .B2(n110754), .ZN(
        n95527) );
  OAI21_X1 U82116 ( .B1(n81629), .B2(n105495), .A(n95528), .ZN(
        \DLX_Datapath/RegisterFile/N25763 ) );
  AOI22_X1 U82117 ( .A1(n104846), .A2(n94682), .B1(n95521), .B2(n110855), .ZN(
        n95528) );
  OAI21_X1 U82118 ( .B1(n106333), .B2(n105495), .A(n95529), .ZN(
        \DLX_Datapath/RegisterFile/N25762 ) );
  AOI22_X1 U82119 ( .A1(n104846), .A2(n94684), .B1(n105494), .B2(n110450), 
        .ZN(n95529) );
  OAI21_X1 U82120 ( .B1(n81315), .B2(n105495), .A(n95530), .ZN(
        \DLX_Datapath/RegisterFile/N25761 ) );
  AOI22_X1 U82121 ( .A1(n104845), .A2(n94686), .B1(n105494), .B2(n110232), 
        .ZN(n95530) );
  OAI21_X1 U82122 ( .B1(n106128), .B2(n105495), .A(n95531), .ZN(
        \DLX_Datapath/RegisterFile/N25760 ) );
  AOI22_X1 U82123 ( .A1(n104844), .A2(n94688), .B1(n105494), .B2(n110549), 
        .ZN(n95531) );
  OAI21_X1 U82124 ( .B1(n106188), .B2(n105495), .A(n95532), .ZN(
        \DLX_Datapath/RegisterFile/N25759 ) );
  AOI22_X1 U82125 ( .A1(n104846), .A2(n94690), .B1(n105494), .B2(n110340), 
        .ZN(n95532) );
  OAI21_X1 U82126 ( .B1(n106165), .B2(n105495), .A(n95533), .ZN(
        \DLX_Datapath/RegisterFile/N25758 ) );
  AOI22_X1 U82127 ( .A1(n104844), .A2(n94692), .B1(n105494), .B2(n110015), 
        .ZN(n95533) );
  OAI21_X1 U82128 ( .B1(n106105), .B2(n105495), .A(n95534), .ZN(
        \DLX_Datapath/RegisterFile/N25757 ) );
  AOI22_X1 U82129 ( .A1(n104845), .A2(n94694), .B1(n105494), .B2(n110122), 
        .ZN(n95534) );
  OAI21_X1 U82130 ( .B1(n81294), .B2(n105495), .A(n95535), .ZN(
        \DLX_Datapath/RegisterFile/N25756 ) );
  AOI22_X1 U82131 ( .A1(n104846), .A2(n94696), .B1(n105494), .B2(n109906), 
        .ZN(n95535) );
  OAI21_X1 U82132 ( .B1(n106109), .B2(n105495), .A(n95536), .ZN(
        \DLX_Datapath/RegisterFile/N25755 ) );
  AOI22_X1 U82133 ( .A1(n104845), .A2(n94698), .B1(n105494), .B2(n109788), 
        .ZN(n95536) );
  OAI21_X1 U82134 ( .B1(n106230), .B2(n105495), .A(n95537), .ZN(
        \DLX_Datapath/RegisterFile/N25754 ) );
  AOI22_X1 U82135 ( .A1(n104846), .A2(n94700), .B1(n105494), .B2(n108162), 
        .ZN(n95537) );
  OAI21_X1 U82136 ( .B1(n81340), .B2(n105495), .A(n95538), .ZN(
        \DLX_Datapath/RegisterFile/N25753 ) );
  AOI22_X1 U82137 ( .A1(n104846), .A2(n94702), .B1(n105494), .B2(n108285), 
        .ZN(n95538) );
  OAI21_X1 U82138 ( .B1(n106238), .B2(n105495), .A(n95539), .ZN(
        \DLX_Datapath/RegisterFile/N25752 ) );
  AOI22_X1 U82139 ( .A1(n104844), .A2(n94704), .B1(n105494), .B2(n108396), 
        .ZN(n95539) );
  OAI21_X1 U82140 ( .B1(n106069), .B2(n105495), .A(n95540), .ZN(
        \DLX_Datapath/RegisterFile/N25751 ) );
  AOI22_X1 U82141 ( .A1(n104846), .A2(n94706), .B1(n105494), .B2(n107634), 
        .ZN(n95540) );
  OAI21_X1 U82142 ( .B1(n81310), .B2(n105495), .A(n95541), .ZN(
        \DLX_Datapath/RegisterFile/N25750 ) );
  AOI22_X1 U82143 ( .A1(n104844), .A2(n94708), .B1(n105493), .B2(n109552), 
        .ZN(n95541) );
  OAI21_X1 U82144 ( .B1(n106244), .B2(n105495), .A(n95542), .ZN(
        \DLX_Datapath/RegisterFile/N25749 ) );
  AOI22_X1 U82145 ( .A1(n104845), .A2(n94710), .B1(n105493), .B2(n108513), 
        .ZN(n95542) );
  OAI21_X1 U82146 ( .B1(n106157), .B2(n105495), .A(n95543), .ZN(
        \DLX_Datapath/RegisterFile/N25748 ) );
  AOI22_X1 U82147 ( .A1(n104846), .A2(n94712), .B1(n105493), .B2(n109657), 
        .ZN(n95543) );
  OAI21_X1 U82148 ( .B1(n106113), .B2(n105495), .A(n95544), .ZN(
        \DLX_Datapath/RegisterFile/N25747 ) );
  AOI22_X1 U82149 ( .A1(n104844), .A2(n94714), .B1(n105493), .B2(n109441), 
        .ZN(n95544) );
  OAI21_X1 U82150 ( .B1(n106007), .B2(n105495), .A(n95545), .ZN(
        \DLX_Datapath/RegisterFile/N25746 ) );
  AOI22_X1 U82151 ( .A1(n104844), .A2(n81259), .B1(n105493), .B2(n108978), 
        .ZN(n95545) );
  OAI21_X1 U82152 ( .B1(n106259), .B2(n105495), .A(n95546), .ZN(
        \DLX_Datapath/RegisterFile/N25745 ) );
  AOI22_X1 U82153 ( .A1(n104844), .A2(n94717), .B1(n105493), .B2(n109326), 
        .ZN(n95546) );
  OAI21_X1 U82154 ( .B1(n81509), .B2(n105495), .A(n95547), .ZN(
        \DLX_Datapath/RegisterFile/N25744 ) );
  AOI22_X1 U82155 ( .A1(n104844), .A2(n94719), .B1(n105493), .B2(n109208), 
        .ZN(n95547) );
  OAI21_X1 U82156 ( .B1(n106048), .B2(n105495), .A(n95548), .ZN(
        \DLX_Datapath/RegisterFile/N25743 ) );
  AOI22_X1 U82157 ( .A1(n104845), .A2(n94721), .B1(n105493), .B2(n109100), 
        .ZN(n95548) );
  OAI21_X1 U82158 ( .B1(n106096), .B2(n105495), .A(n95549), .ZN(
        \DLX_Datapath/RegisterFile/N25742 ) );
  AOI22_X1 U82159 ( .A1(n104846), .A2(n94723), .B1(n105493), .B2(n108635), 
        .ZN(n95549) );
  OAI21_X1 U82160 ( .B1(n106053), .B2(n105495), .A(n95550), .ZN(
        \DLX_Datapath/RegisterFile/N25741 ) );
  AOI22_X1 U82161 ( .A1(n104845), .A2(n94725), .B1(n105493), .B2(n108862), 
        .ZN(n95550) );
  OAI21_X1 U82162 ( .B1(n105219), .B2(n105495), .A(n95551), .ZN(
        \DLX_Datapath/RegisterFile/N25740 ) );
  AOI22_X1 U82163 ( .A1(n104845), .A2(n94727), .B1(n105493), .B2(n108750), 
        .ZN(n95551) );
  OAI21_X1 U82164 ( .B1(n106266), .B2(n105495), .A(n95552), .ZN(
        \DLX_Datapath/RegisterFile/N25739 ) );
  AOI22_X1 U82165 ( .A1(n104846), .A2(n94729), .B1(n105493), .B2(n107290), 
        .ZN(n95552) );
  AOI21_X1 U82166 ( .B1(n95553), .B2(n105602), .A(n95554), .ZN(n95521) );
  OAI21_X1 U82167 ( .B1(n95555), .B2(n94999), .A(n105199), .ZN(n95553) );
  NOR2_X1 U82168 ( .A1(n95556), .A2(n95555), .ZN(n95520) );
  OR2_X1 U82169 ( .A1(n95554), .A2(n94999), .ZN(n95556) );
  NOR2_X1 U82170 ( .A1(n95518), .A2(n105089), .ZN(n95554) );
  NAND2_X1 U82171 ( .A1(n94367), .A2(n105133), .ZN(n95518) );
  OAI21_X1 U82172 ( .B1(n106146), .B2(n105918), .A(n95557), .ZN(
        \DLX_Datapath/RegisterFile/N25738 ) );
  AOI22_X1 U82173 ( .A1(n70295), .A2(n81776), .B1(n105916), .B2(n81360), .ZN(
        n95557) );
  OAI21_X1 U82174 ( .B1(n105968), .B2(n105918), .A(n95558), .ZN(
        \DLX_Datapath/RegisterFile/N25737 ) );
  AOI22_X1 U82175 ( .A1(n70437), .A2(n105001), .B1(n94511), .B2(n81777), .ZN(
        n95558) );
  OAI21_X1 U82176 ( .B1(n81299), .B2(n105917), .A(n95559), .ZN(
        \DLX_Datapath/RegisterFile/N25735 ) );
  AOI22_X1 U82177 ( .A1(n70151), .A2(n105000), .B1(n105916), .B2(n81301), .ZN(
        n95559) );
  OAI21_X1 U82178 ( .B1(n106203), .B2(n105918), .A(n95560), .ZN(
        \DLX_Datapath/RegisterFile/N25734 ) );
  AOI22_X1 U82179 ( .A1(n73997), .A2(n105000), .B1(n105915), .B2(n81308), .ZN(
        n95560) );
  OAI21_X1 U82180 ( .B1(n81408), .B2(n105917), .A(n95561), .ZN(
        \DLX_Datapath/RegisterFile/N25733 ) );
  AOI22_X1 U82181 ( .A1(n70584), .A2(n105001), .B1(n94516), .B2(n81777), .ZN(
        n95561) );
  OAI21_X1 U82182 ( .B1(n81629), .B2(n105918), .A(n95562), .ZN(
        \DLX_Datapath/RegisterFile/N25731 ) );
  AOI22_X1 U82183 ( .A1(n74278), .A2(n105000), .B1(n94519), .B2(n105916), .ZN(
        n95562) );
  OAI21_X1 U82184 ( .B1(n106332), .B2(n105918), .A(n95563), .ZN(
        \DLX_Datapath/RegisterFile/N25730 ) );
  AOI22_X1 U82185 ( .A1(n73714), .A2(n105001), .B1(n105915), .B2(n80192), .ZN(
        n95563) );
  OAI21_X1 U82186 ( .B1(n81315), .B2(n105918), .A(n95564), .ZN(
        \DLX_Datapath/RegisterFile/N25729 ) );
  AOI22_X1 U82187 ( .A1(n73418), .A2(n81776), .B1(n105916), .B2(n81474), .ZN(
        n95564) );
  OAI21_X1 U82188 ( .B1(n106129), .B2(n105918), .A(n95565), .ZN(
        \DLX_Datapath/RegisterFile/N25728 ) );
  AOI22_X1 U82189 ( .A1(n73855), .A2(n81776), .B1(n94523), .B2(n81777), .ZN(
        n95565) );
  OAI21_X1 U82190 ( .B1(n106186), .B2(n105918), .A(n95566), .ZN(
        \DLX_Datapath/RegisterFile/N25727 ) );
  AOI22_X1 U82191 ( .A1(n73567), .A2(n105000), .B1(n105915), .B2(n106061), 
        .ZN(n95566) );
  OAI21_X1 U82192 ( .B1(n106165), .B2(n105918), .A(n95567), .ZN(
        \DLX_Datapath/RegisterFile/N25726 ) );
  AOI22_X1 U82193 ( .A1(n73129), .A2(n105000), .B1(n105916), .B2(n81347), .ZN(
        n95567) );
  OAI21_X1 U82194 ( .B1(n106104), .B2(n105918), .A(n95568), .ZN(
        \DLX_Datapath/RegisterFile/N25725 ) );
  AOI22_X1 U82195 ( .A1(n73271), .A2(n105001), .B1(n94527), .B2(n81777), .ZN(
        n95568) );
  OAI21_X1 U82196 ( .B1(n81294), .B2(n105918), .A(n95569), .ZN(
        \DLX_Datapath/RegisterFile/N25724 ) );
  AOI22_X1 U82197 ( .A1(n72987), .A2(n105000), .B1(n105915), .B2(n81297), .ZN(
        n95569) );
  OAI21_X1 U82198 ( .B1(n106109), .B2(n105918), .A(n95570), .ZN(
        \DLX_Datapath/RegisterFile/N25723 ) );
  AOI22_X1 U82199 ( .A1(n72837), .A2(n105001), .B1(n94530), .B2(n105915), .ZN(
        n95570) );
  OAI21_X1 U82200 ( .B1(n106230), .B2(n105918), .A(n95571), .ZN(
        \DLX_Datapath/RegisterFile/N25722 ) );
  AOI22_X1 U82201 ( .A1(n70733), .A2(n105000), .B1(n105916), .B2(n81286), .ZN(
        n95571) );
  OAI21_X1 U82202 ( .B1(n106172), .B2(n105918), .A(n95572), .ZN(
        \DLX_Datapath/RegisterFile/N25721 ) );
  AOI22_X1 U82203 ( .A1(n70892), .A2(n105001), .B1(n105915), .B2(n106168), 
        .ZN(n95572) );
  OAI21_X1 U82204 ( .B1(n81281), .B2(n105918), .A(n95573), .ZN(
        \DLX_Datapath/RegisterFile/N25720 ) );
  AOI22_X1 U82205 ( .A1(n71037), .A2(n105001), .B1(n105916), .B2(n81283), .ZN(
        n95573) );
  OAI21_X1 U82206 ( .B1(n106069), .B2(n105917), .A(n95574), .ZN(
        \DLX_Datapath/RegisterFile/N25719 ) );
  AOI22_X1 U82207 ( .A1(n69998), .A2(n81776), .B1(n105915), .B2(n81453), .ZN(
        n95574) );
  OAI21_X1 U82208 ( .B1(n81310), .B2(n105917), .A(n95575), .ZN(
        \DLX_Datapath/RegisterFile/N25718 ) );
  AOI22_X1 U82209 ( .A1(n72527), .A2(n81776), .B1(n94536), .B2(n81777), .ZN(
        n95575) );
  OAI21_X1 U82210 ( .B1(n106158), .B2(n105917), .A(n95576), .ZN(
        \DLX_Datapath/RegisterFile/N25716 ) );
  AOI22_X1 U82211 ( .A1(n72669), .A2(n105000), .B1(n105916), .B2(n81351), .ZN(
        n95576) );
  OAI21_X1 U82212 ( .B1(n106116), .B2(n105917), .A(n95577), .ZN(
        \DLX_Datapath/RegisterFile/N25715 ) );
  AOI22_X1 U82213 ( .A1(n72379), .A2(n105000), .B1(n105915), .B2(n106020), 
        .ZN(n95577) );
  OAI21_X1 U82214 ( .B1(n81588), .B2(n105917), .A(n95578), .ZN(
        \DLX_Datapath/RegisterFile/N25714 ) );
  AOI22_X1 U82215 ( .A1(n71779), .A2(n105001), .B1(n94541), .B2(n81777), .ZN(
        n95578) );
  OAI21_X1 U82216 ( .B1(n81509), .B2(n105917), .A(n95579), .ZN(
        \DLX_Datapath/RegisterFile/N25712 ) );
  AOI22_X1 U82217 ( .A1(n72077), .A2(n81776), .B1(n105625), .B2(n81777), .ZN(
        n95579) );
  OAI21_X1 U82218 ( .B1(n106048), .B2(n105917), .A(n95580), .ZN(
        \DLX_Datapath/RegisterFile/N25711 ) );
  AOI22_X1 U82219 ( .A1(n71933), .A2(n105001), .B1(n94546), .B2(n105915), .ZN(
        n95580) );
  OAI21_X1 U82220 ( .B1(n106093), .B2(n105917), .A(n95581), .ZN(
        \DLX_Datapath/RegisterFile/N25710 ) );
  AOI22_X1 U82221 ( .A1(n71335), .A2(n105000), .B1(n94548), .B2(n81777), .ZN(
        n95581) );
  OAI21_X1 U82222 ( .B1(n106056), .B2(n105917), .A(n95582), .ZN(
        \DLX_Datapath/RegisterFile/N25709 ) );
  AOI22_X1 U82223 ( .A1(n71630), .A2(n105001), .B1(n81783), .B2(n105916), .ZN(
        n95582) );
  OAI21_X1 U82224 ( .B1(n105220), .B2(n105917), .A(n95583), .ZN(
        \DLX_Datapath/RegisterFile/N25708 ) );
  AOI22_X1 U82225 ( .A1(n71486), .A2(n105000), .B1(n105916), .B2(n80188), .ZN(
        n95583) );
  OAI21_X1 U82226 ( .B1(n106266), .B2(n105917), .A(n95584), .ZN(
        \DLX_Datapath/RegisterFile/N25707 ) );
  AOI22_X1 U82227 ( .A1(n69595), .A2(n81776), .B1(n105915), .B2(n81265), .ZN(
        n95584) );
  NOR2_X1 U82228 ( .A1(n95585), .A2(n95586), .ZN(n81777) );
  AOI21_X1 U82229 ( .B1(n95450), .B2(n94398), .A(n95586), .ZN(n81776) );
  NOR2_X1 U82230 ( .A1(n81774), .A2(n105089), .ZN(n95586) );
  NAND2_X1 U82231 ( .A1(n105134), .A2(n94399), .ZN(n81774) );
  OAI21_X1 U82232 ( .B1(n106146), .B2(n105492), .A(n95588), .ZN(
        \DLX_Datapath/RegisterFile/N25706 ) );
  AOI22_X1 U82233 ( .A1(n105490), .A2(n107858), .B1(n95590), .B2(n94559), .ZN(
        n95588) );
  OAI21_X1 U82234 ( .B1(n105968), .B2(n105492), .A(n95591), .ZN(
        \DLX_Datapath/RegisterFile/N25705 ) );
  AOI22_X1 U82235 ( .A1(n105489), .A2(n107955), .B1(n104972), .B2(n94562), 
        .ZN(n95591) );
  OAI21_X1 U82236 ( .B1(n106136), .B2(n105492), .A(n95592), .ZN(
        \DLX_Datapath/RegisterFile/N25704 ) );
  AOI22_X1 U82237 ( .A1(n105490), .A2(n107217), .B1(n95590), .B2(n94564), .ZN(
        n95592) );
  OAI21_X1 U82238 ( .B1(n81299), .B2(n105492), .A(n95593), .ZN(
        \DLX_Datapath/RegisterFile/N25703 ) );
  AOI22_X1 U82239 ( .A1(n105489), .A2(n107755), .B1(n104973), .B2(n94566), 
        .ZN(n95593) );
  OAI21_X1 U82240 ( .B1(n106203), .B2(n105492), .A(n95594), .ZN(
        \DLX_Datapath/RegisterFile/N25702 ) );
  AOI22_X1 U82241 ( .A1(n105490), .A2(n110658), .B1(n104972), .B2(n94568), 
        .ZN(n95594) );
  OAI21_X1 U82242 ( .B1(n81408), .B2(n105492), .A(n95595), .ZN(
        \DLX_Datapath/RegisterFile/N25701 ) );
  AOI22_X1 U82243 ( .A1(n105489), .A2(n108057), .B1(n104972), .B2(n94570), 
        .ZN(n95595) );
  OAI21_X1 U82244 ( .B1(n106256), .B2(n105492), .A(n95596), .ZN(
        \DLX_Datapath/RegisterFile/N25700 ) );
  AOI22_X1 U82245 ( .A1(n105490), .A2(n110755), .B1(n104972), .B2(n94572), 
        .ZN(n95596) );
  OAI21_X1 U82246 ( .B1(n105990), .B2(n105492), .A(n95597), .ZN(
        \DLX_Datapath/RegisterFile/N25699 ) );
  AOI22_X1 U82247 ( .A1(n105489), .A2(n110856), .B1(n104973), .B2(n94574), 
        .ZN(n95597) );
  OAI21_X1 U82248 ( .B1(n106331), .B2(n105492), .A(n95598), .ZN(
        \DLX_Datapath/RegisterFile/N25698 ) );
  AOI22_X1 U82249 ( .A1(n105489), .A2(n110451), .B1(n104972), .B2(n94576), 
        .ZN(n95598) );
  OAI21_X1 U82250 ( .B1(n81315), .B2(n105491), .A(n95599), .ZN(
        \DLX_Datapath/RegisterFile/N25697 ) );
  AOI22_X1 U82251 ( .A1(n105490), .A2(n110233), .B1(n104973), .B2(n94578), 
        .ZN(n95599) );
  OAI21_X1 U82252 ( .B1(n81383), .B2(n105491), .A(n95600), .ZN(
        \DLX_Datapath/RegisterFile/N25696 ) );
  AOI22_X1 U82253 ( .A1(n95589), .A2(n110550), .B1(n104972), .B2(n94580), .ZN(
        n95600) );
  OAI21_X1 U82254 ( .B1(n81318), .B2(n105491), .A(n95601), .ZN(
        \DLX_Datapath/RegisterFile/N25695 ) );
  AOI22_X1 U82255 ( .A1(n105489), .A2(n110341), .B1(n104973), .B2(n94582), 
        .ZN(n95601) );
  OAI21_X1 U82256 ( .B1(n106163), .B2(n105491), .A(n95602), .ZN(
        \DLX_Datapath/RegisterFile/N25694 ) );
  AOI22_X1 U82257 ( .A1(n95589), .A2(n110016), .B1(n104973), .B2(n94584), .ZN(
        n95602) );
  OAI21_X1 U82258 ( .B1(n106104), .B2(n105491), .A(n95603), .ZN(
        \DLX_Datapath/RegisterFile/N25693 ) );
  AOI22_X1 U82259 ( .A1(n95589), .A2(n110123), .B1(n95590), .B2(n94586), .ZN(
        n95603) );
  OAI21_X1 U82260 ( .B1(n81294), .B2(n105491), .A(n95604), .ZN(
        \DLX_Datapath/RegisterFile/N25692 ) );
  AOI22_X1 U82261 ( .A1(n105489), .A2(n109907), .B1(n104972), .B2(n94588), 
        .ZN(n95604) );
  OAI21_X1 U82262 ( .B1(n106110), .B2(n105491), .A(n95605), .ZN(
        \DLX_Datapath/RegisterFile/N25691 ) );
  AOI22_X1 U82263 ( .A1(n95589), .A2(n109789), .B1(n104972), .B2(n94590), .ZN(
        n95605) );
  OAI21_X1 U82264 ( .B1(n106230), .B2(n105491), .A(n95606), .ZN(
        \DLX_Datapath/RegisterFile/N25690 ) );
  AOI22_X1 U82265 ( .A1(n95589), .A2(n108163), .B1(n104973), .B2(n94592), .ZN(
        n95606) );
  OAI21_X1 U82266 ( .B1(n81340), .B2(n105491), .A(n95607), .ZN(
        \DLX_Datapath/RegisterFile/N25689 ) );
  AOI22_X1 U82267 ( .A1(n95589), .A2(n108286), .B1(n104972), .B2(n94594), .ZN(
        n95607) );
  OAI21_X1 U82268 ( .B1(n106235), .B2(n105491), .A(n95608), .ZN(
        \DLX_Datapath/RegisterFile/N25688 ) );
  AOI22_X1 U82269 ( .A1(n95589), .A2(n108397), .B1(n104972), .B2(n94596), .ZN(
        n95608) );
  OAI21_X1 U82270 ( .B1(n106069), .B2(n105491), .A(n95609), .ZN(
        \DLX_Datapath/RegisterFile/N25687 ) );
  AOI22_X1 U82271 ( .A1(n95589), .A2(n107635), .B1(n104972), .B2(n94598), .ZN(
        n95609) );
  OAI21_X1 U82272 ( .B1(n81310), .B2(n105491), .A(n95610), .ZN(
        \DLX_Datapath/RegisterFile/N25686 ) );
  AOI22_X1 U82273 ( .A1(n105489), .A2(n109553), .B1(n104973), .B2(n94600), 
        .ZN(n95610) );
  OAI21_X1 U82274 ( .B1(n106244), .B2(n105492), .A(n95611), .ZN(
        \DLX_Datapath/RegisterFile/N25685 ) );
  AOI22_X1 U82275 ( .A1(n105490), .A2(n108514), .B1(n104973), .B2(n94602), 
        .ZN(n95611) );
  OAI21_X1 U82276 ( .B1(n81349), .B2(n105492), .A(n95612), .ZN(
        \DLX_Datapath/RegisterFile/N25684 ) );
  AOI22_X1 U82277 ( .A1(n105489), .A2(n109658), .B1(n104973), .B2(n94604), 
        .ZN(n95612) );
  OAI21_X1 U82278 ( .B1(n106113), .B2(n105491), .A(n95613), .ZN(
        \DLX_Datapath/RegisterFile/N25683 ) );
  AOI22_X1 U82279 ( .A1(n105490), .A2(n109442), .B1(n95590), .B2(n94606), .ZN(
        n95613) );
  OAI21_X1 U82280 ( .B1(n106009), .B2(n105492), .A(n95614), .ZN(
        \DLX_Datapath/RegisterFile/N25682 ) );
  AOI22_X1 U82281 ( .A1(n105489), .A2(n108979), .B1(n95590), .B2(n94608), .ZN(
        n95614) );
  OAI21_X1 U82282 ( .B1(n106259), .B2(n105492), .A(n95615), .ZN(
        \DLX_Datapath/RegisterFile/N25681 ) );
  AOI22_X1 U82283 ( .A1(n105490), .A2(n109327), .B1(n104972), .B2(n94610), 
        .ZN(n95615) );
  OAI21_X1 U82284 ( .B1(n81509), .B2(n105491), .A(n95616), .ZN(
        \DLX_Datapath/RegisterFile/N25680 ) );
  AOI22_X1 U82285 ( .A1(n105489), .A2(n109209), .B1(n104973), .B2(n94612), 
        .ZN(n95616) );
  OAI21_X1 U82286 ( .B1(n106050), .B2(n105492), .A(n95617), .ZN(
        \DLX_Datapath/RegisterFile/N25679 ) );
  AOI22_X1 U82287 ( .A1(n105490), .A2(n109101), .B1(n104972), .B2(n94614), 
        .ZN(n95617) );
  OAI21_X1 U82288 ( .B1(n106094), .B2(n105491), .A(n95618), .ZN(
        \DLX_Datapath/RegisterFile/N25678 ) );
  AOI22_X1 U82289 ( .A1(n105489), .A2(n108636), .B1(n95590), .B2(n94616), .ZN(
        n95618) );
  OAI21_X1 U82290 ( .B1(n106054), .B2(n105492), .A(n95619), .ZN(
        \DLX_Datapath/RegisterFile/N25677 ) );
  AOI22_X1 U82291 ( .A1(n105490), .A2(n108863), .B1(n104972), .B2(n94618), 
        .ZN(n95619) );
  OAI21_X1 U82292 ( .B1(n105217), .B2(n105492), .A(n95620), .ZN(
        \DLX_Datapath/RegisterFile/N25676 ) );
  AOI22_X1 U82293 ( .A1(n105490), .A2(n108751), .B1(n95590), .B2(n94620), .ZN(
        n95620) );
  OAI21_X1 U82294 ( .B1(n106266), .B2(n105491), .A(n95621), .ZN(
        \DLX_Datapath/RegisterFile/N25675 ) );
  AOI22_X1 U82295 ( .A1(n105489), .A2(n107291), .B1(n104973), .B2(n94622), 
        .ZN(n95621) );
  NOR2_X1 U82296 ( .A1(n95585), .A2(n95622), .ZN(n95590) );
  NOR2_X1 U82297 ( .A1(n95623), .A2(n95622), .ZN(n95589) );
  NOR2_X1 U82298 ( .A1(n95587), .A2(n105089), .ZN(n95622) );
  NAND2_X1 U82299 ( .A1(n94434), .A2(n105134), .ZN(n95587) );
  OAI21_X1 U82300 ( .B1(n81299), .B2(n105966), .A(n95624), .ZN(
        \DLX_Datapath/RegisterFile/N25671 ) );
  AOI22_X1 U82301 ( .A1(n105964), .A2(n81377), .B1(n70153), .B2(n104990), .ZN(
        n95624) );
  OAI21_X1 U82302 ( .B1(n106203), .B2(n105966), .A(n95625), .ZN(
        \DLX_Datapath/RegisterFile/N25670 ) );
  AOI22_X1 U82303 ( .A1(n81660), .A2(n81428), .B1(n73999), .B2(n104991), .ZN(
        n95625) );
  OAI21_X1 U82304 ( .B1(n81408), .B2(n105966), .A(n95626), .ZN(
        \DLX_Datapath/RegisterFile/N25669 ) );
  AOI22_X1 U82305 ( .A1(n105964), .A2(n81410), .B1(n70586), .B2(n104991), .ZN(
        n95626) );
  OAI21_X1 U82306 ( .B1(n106256), .B2(n105967), .A(n95627), .ZN(
        \DLX_Datapath/RegisterFile/N25668 ) );
  AOI22_X1 U82307 ( .A1(n81700), .A2(n105965), .B1(n74140), .B2(n104991), .ZN(
        n95627) );
  OAI21_X1 U82308 ( .B1(n81629), .B2(n105967), .A(n95628), .ZN(
        \DLX_Datapath/RegisterFile/N25667 ) );
  AOI22_X1 U82309 ( .A1(n105965), .A2(n81632), .B1(n74280), .B2(n104990), .ZN(
        n95628) );
  OAI21_X1 U82310 ( .B1(n106331), .B2(n105967), .A(n95629), .ZN(
        \DLX_Datapath/RegisterFile/N25666 ) );
  AOI22_X1 U82311 ( .A1(n105965), .A2(n81414), .B1(n73716), .B2(n104991), .ZN(
        n95629) );
  OAI21_X1 U82312 ( .B1(n106192), .B2(n105967), .A(n95630), .ZN(
        \DLX_Datapath/RegisterFile/N25665 ) );
  AOI22_X1 U82313 ( .A1(n105965), .A2(n81317), .B1(n73420), .B2(n81661), .ZN(
        n95630) );
  OAI21_X1 U82314 ( .B1(n106129), .B2(n105967), .A(n95631), .ZN(
        \DLX_Datapath/RegisterFile/N25664 ) );
  AOI22_X1 U82315 ( .A1(n105964), .A2(n81386), .B1(n73857), .B2(n81661), .ZN(
        n95631) );
  OAI21_X1 U82316 ( .B1(n106186), .B2(n105967), .A(n95632), .ZN(
        \DLX_Datapath/RegisterFile/N25663 ) );
  AOI22_X1 U82317 ( .A1(n105965), .A2(n81320), .B1(n73569), .B2(n104990), .ZN(
        n95632) );
  OAI21_X1 U82318 ( .B1(n106164), .B2(n105967), .A(n95633), .ZN(
        \DLX_Datapath/RegisterFile/N25662 ) );
  AOI22_X1 U82319 ( .A1(n105964), .A2(n81604), .B1(n73131), .B2(n104990), .ZN(
        n95633) );
  OAI21_X1 U82320 ( .B1(n106106), .B2(n105967), .A(n95634), .ZN(
        \DLX_Datapath/RegisterFile/N25661 ) );
  AOI22_X1 U82321 ( .A1(n105965), .A2(n81405), .B1(n73273), .B2(n104991), .ZN(
        n95634) );
  OAI21_X1 U82322 ( .B1(n81294), .B2(n105967), .A(n95635), .ZN(
        \DLX_Datapath/RegisterFile/N25660 ) );
  AOI22_X1 U82323 ( .A1(n105965), .A2(n81402), .B1(n72989), .B2(n104990), .ZN(
        n95635) );
  OAI21_X1 U82324 ( .B1(n106110), .B2(n105967), .A(n95636), .ZN(
        \DLX_Datapath/RegisterFile/N25659 ) );
  AOI22_X1 U82325 ( .A1(n105965), .A2(n81400), .B1(n72839), .B2(n104991), .ZN(
        n95636) );
  OAI21_X1 U82326 ( .B1(n106171), .B2(n105967), .A(n95637), .ZN(
        \DLX_Datapath/RegisterFile/N25657 ) );
  AOI22_X1 U82327 ( .A1(n105965), .A2(n81373), .B1(n70894), .B2(n104990), .ZN(
        n95637) );
  OAI21_X1 U82328 ( .B1(n81281), .B2(n105967), .A(n95638), .ZN(
        \DLX_Datapath/RegisterFile/N25656 ) );
  AOI22_X1 U82329 ( .A1(n105965), .A2(n81322), .B1(n71039), .B2(n104991), .ZN(
        n95638) );
  OAI21_X1 U82330 ( .B1(n106069), .B2(n105967), .A(n95639), .ZN(
        \DLX_Datapath/RegisterFile/N25655 ) );
  AOI22_X1 U82331 ( .A1(n105965), .A2(n81506), .B1(n70000), .B2(n104991), .ZN(
        n95639) );
  OAI21_X1 U82332 ( .B1(n81310), .B2(n105966), .A(n95640), .ZN(
        \DLX_Datapath/RegisterFile/N25654 ) );
  AOI22_X1 U82333 ( .A1(n105964), .A2(n81313), .B1(n72529), .B2(n104990), .ZN(
        n95640) );
  OAI21_X1 U82334 ( .B1(n106244), .B2(n105966), .A(n95641), .ZN(
        \DLX_Datapath/RegisterFile/N25653 ) );
  AOI22_X1 U82335 ( .A1(n81660), .A2(n81330), .B1(n71188), .B2(n81661), .ZN(
        n95641) );
  OAI21_X1 U82336 ( .B1(n81349), .B2(n105966), .A(n95642), .ZN(
        \DLX_Datapath/RegisterFile/N25652 ) );
  AOI22_X1 U82337 ( .A1(n105964), .A2(n81425), .B1(n72671), .B2(n104991), .ZN(
        n95642) );
  OAI21_X1 U82338 ( .B1(n106113), .B2(n105966), .A(n95643), .ZN(
        \DLX_Datapath/RegisterFile/N25651 ) );
  AOI22_X1 U82339 ( .A1(n81660), .A2(n81396), .B1(n72381), .B2(n81661), .ZN(
        n95643) );
  OAI21_X1 U82340 ( .B1(n81588), .B2(n105966), .A(n95644), .ZN(
        \DLX_Datapath/RegisterFile/N25650 ) );
  AOI22_X1 U82341 ( .A1(n81660), .A2(n81590), .B1(n71781), .B2(n104990), .ZN(
        n95644) );
  OAI21_X1 U82342 ( .B1(n81267), .B2(n105966), .A(n95645), .ZN(
        \DLX_Datapath/RegisterFile/N25649 ) );
  AOI22_X1 U82343 ( .A1(n105964), .A2(n81423), .B1(n72230), .B2(n104990), .ZN(
        n95645) );
  OAI21_X1 U82344 ( .B1(n81509), .B2(n105966), .A(n95646), .ZN(
        \DLX_Datapath/RegisterFile/N25648 ) );
  AOI22_X1 U82345 ( .A1(n81660), .A2(n81511), .B1(n72079), .B2(n104991), .ZN(
        n95646) );
  OAI21_X1 U82346 ( .B1(n106049), .B2(n105966), .A(n95647), .ZN(
        \DLX_Datapath/RegisterFile/N25647 ) );
  AOI22_X1 U82347 ( .A1(n105964), .A2(n81503), .B1(n71935), .B2(n104991), .ZN(
        n95647) );
  OAI21_X1 U82348 ( .B1(n81415), .B2(n105966), .A(n95648), .ZN(
        \DLX_Datapath/RegisterFile/N25646 ) );
  AOI22_X1 U82349 ( .A1(n105965), .A2(n81417), .B1(n71337), .B2(n81661), .ZN(
        n95648) );
  OAI21_X1 U82350 ( .B1(n105216), .B2(n105966), .A(n95649), .ZN(
        \DLX_Datapath/RegisterFile/N25644 ) );
  AOI22_X1 U82351 ( .A1(n105964), .A2(n81335), .B1(n71488), .B2(n81661), .ZN(
        n95649) );
  OAI21_X1 U82352 ( .B1(n106266), .B2(n105966), .A(n95650), .ZN(
        \DLX_Datapath/RegisterFile/N25643 ) );
  AOI22_X1 U82353 ( .A1(n105964), .A2(n81327), .B1(n69597), .B2(n104990), .ZN(
        n95650) );
  NOR2_X1 U82354 ( .A1(n95651), .A2(n95623), .ZN(n81661) );
  AOI21_X1 U82355 ( .B1(n105205), .B2(n95585), .A(n105601), .ZN(n95623) );
  NOR2_X1 U82356 ( .A1(n95585), .A2(n95651), .ZN(n81660) );
  NOR2_X1 U82357 ( .A1(n81658), .A2(n105091), .ZN(n95651) );
  OR2_X1 U82358 ( .A1(n95517), .A2(n95131), .ZN(n95585) );
  NAND2_X1 U82359 ( .A1(n105133), .A2(n95132), .ZN(n81658) );
  OAI21_X1 U82360 ( .B1(n106146), .B2(n95652), .A(n95653), .ZN(
        \DLX_Datapath/RegisterFile/N25642 ) );
  AOI22_X1 U82361 ( .A1(n105487), .A2(n94667), .B1(n104938), .B2(n107859), 
        .ZN(n95653) );
  OAI21_X1 U82362 ( .B1(n105969), .B2(n95652), .A(n95656), .ZN(
        \DLX_Datapath/RegisterFile/N25641 ) );
  AOI22_X1 U82363 ( .A1(n105486), .A2(n94670), .B1(n104939), .B2(n107956), 
        .ZN(n95656) );
  OAI21_X1 U82364 ( .B1(n106135), .B2(n95652), .A(n95657), .ZN(
        \DLX_Datapath/RegisterFile/N25640 ) );
  AOI22_X1 U82365 ( .A1(n105487), .A2(n94672), .B1(n104938), .B2(n107218), 
        .ZN(n95657) );
  OAI21_X1 U82366 ( .B1(n106210), .B2(n95652), .A(n95658), .ZN(
        \DLX_Datapath/RegisterFile/N25639 ) );
  AOI22_X1 U82367 ( .A1(n105486), .A2(n94674), .B1(n104940), .B2(n107756), 
        .ZN(n95658) );
  OAI21_X1 U82368 ( .B1(n106203), .B2(n95652), .A(n95659), .ZN(
        \DLX_Datapath/RegisterFile/N25638 ) );
  AOI22_X1 U82369 ( .A1(n105487), .A2(n94676), .B1(n104938), .B2(n110659), 
        .ZN(n95659) );
  OAI21_X1 U82370 ( .B1(n81408), .B2(n105488), .A(n95660), .ZN(
        \DLX_Datapath/RegisterFile/N25637 ) );
  AOI22_X1 U82371 ( .A1(n105486), .A2(n94678), .B1(n104939), .B2(n108058), 
        .ZN(n95660) );
  OAI21_X1 U82372 ( .B1(n106254), .B2(n95652), .A(n95661), .ZN(
        \DLX_Datapath/RegisterFile/N25636 ) );
  AOI22_X1 U82373 ( .A1(n105487), .A2(n94680), .B1(n104939), .B2(n110756), 
        .ZN(n95661) );
  OAI21_X1 U82374 ( .B1(n81629), .B2(n105488), .A(n95662), .ZN(
        \DLX_Datapath/RegisterFile/N25635 ) );
  AOI22_X1 U82375 ( .A1(n105486), .A2(n94682), .B1(n104940), .B2(n110857), 
        .ZN(n95662) );
  OAI21_X1 U82376 ( .B1(n80190), .B2(n105488), .A(n95663), .ZN(
        \DLX_Datapath/RegisterFile/N25634 ) );
  AOI22_X1 U82377 ( .A1(n105486), .A2(n94684), .B1(n104939), .B2(n110452), 
        .ZN(n95663) );
  OAI21_X1 U82378 ( .B1(n81315), .B2(n105488), .A(n95664), .ZN(
        \DLX_Datapath/RegisterFile/N25633 ) );
  AOI22_X1 U82379 ( .A1(n105485), .A2(n94686), .B1(n104938), .B2(n110234), 
        .ZN(n95664) );
  OAI21_X1 U82380 ( .B1(n81383), .B2(n105488), .A(n95665), .ZN(
        \DLX_Datapath/RegisterFile/N25632 ) );
  AOI22_X1 U82381 ( .A1(n105485), .A2(n94688), .B1(n104939), .B2(n110551), 
        .ZN(n95665) );
  OAI21_X1 U82382 ( .B1(n81318), .B2(n105488), .A(n95666), .ZN(
        \DLX_Datapath/RegisterFile/N25631 ) );
  AOI22_X1 U82383 ( .A1(n105485), .A2(n94690), .B1(n104940), .B2(n110342), 
        .ZN(n95666) );
  OAI21_X1 U82384 ( .B1(n106162), .B2(n105488), .A(n95667), .ZN(
        \DLX_Datapath/RegisterFile/N25630 ) );
  AOI22_X1 U82385 ( .A1(n105485), .A2(n94692), .B1(n104940), .B2(n110017), 
        .ZN(n95667) );
  OAI21_X1 U82386 ( .B1(n106106), .B2(n105488), .A(n95668), .ZN(
        \DLX_Datapath/RegisterFile/N25629 ) );
  AOI22_X1 U82387 ( .A1(n105485), .A2(n94694), .B1(n104938), .B2(n110124), 
        .ZN(n95668) );
  OAI21_X1 U82388 ( .B1(n81294), .B2(n105488), .A(n95669), .ZN(
        \DLX_Datapath/RegisterFile/N25628 ) );
  AOI22_X1 U82389 ( .A1(n105485), .A2(n94696), .B1(n104938), .B2(n109908), 
        .ZN(n95669) );
  OAI21_X1 U82390 ( .B1(n106111), .B2(n105488), .A(n95670), .ZN(
        \DLX_Datapath/RegisterFile/N25627 ) );
  AOI22_X1 U82391 ( .A1(n105485), .A2(n94698), .B1(n104939), .B2(n109790), 
        .ZN(n95670) );
  OAI21_X1 U82392 ( .B1(n106230), .B2(n105488), .A(n95671), .ZN(
        \DLX_Datapath/RegisterFile/N25626 ) );
  AOI22_X1 U82393 ( .A1(n105485), .A2(n94700), .B1(n104940), .B2(n108164), 
        .ZN(n95671) );
  OAI21_X1 U82394 ( .B1(n81340), .B2(n105488), .A(n95672), .ZN(
        \DLX_Datapath/RegisterFile/N25625 ) );
  AOI22_X1 U82395 ( .A1(n105485), .A2(n94702), .B1(n104939), .B2(n108287), 
        .ZN(n95672) );
  OAI21_X1 U82396 ( .B1(n106237), .B2(n105488), .A(n95673), .ZN(
        \DLX_Datapath/RegisterFile/N25624 ) );
  AOI22_X1 U82397 ( .A1(n105485), .A2(n94704), .B1(n104938), .B2(n108398), 
        .ZN(n95673) );
  OAI21_X1 U82398 ( .B1(n106069), .B2(n105488), .A(n95674), .ZN(
        \DLX_Datapath/RegisterFile/N25623 ) );
  AOI22_X1 U82399 ( .A1(n105485), .A2(n94706), .B1(n104939), .B2(n107636), 
        .ZN(n95674) );
  OAI21_X1 U82400 ( .B1(n81310), .B2(n105488), .A(n95675), .ZN(
        \DLX_Datapath/RegisterFile/N25622 ) );
  AOI22_X1 U82401 ( .A1(n105486), .A2(n94708), .B1(n104940), .B2(n109554), 
        .ZN(n95675) );
  OAI21_X1 U82402 ( .B1(n106244), .B2(n105488), .A(n95676), .ZN(
        \DLX_Datapath/RegisterFile/N25621 ) );
  AOI22_X1 U82403 ( .A1(n105487), .A2(n94710), .B1(n104940), .B2(n108515), 
        .ZN(n95676) );
  OAI21_X1 U82404 ( .B1(n81349), .B2(n105488), .A(n95677), .ZN(
        \DLX_Datapath/RegisterFile/N25620 ) );
  AOI22_X1 U82405 ( .A1(n105486), .A2(n94712), .B1(n104940), .B2(n109659), 
        .ZN(n95677) );
  OAI21_X1 U82406 ( .B1(n106113), .B2(n105488), .A(n95678), .ZN(
        \DLX_Datapath/RegisterFile/N25619 ) );
  AOI22_X1 U82407 ( .A1(n105487), .A2(n94714), .B1(n104938), .B2(n109443), 
        .ZN(n95678) );
  OAI21_X1 U82408 ( .B1(n106011), .B2(n105488), .A(n95679), .ZN(
        \DLX_Datapath/RegisterFile/N25618 ) );
  AOI22_X1 U82409 ( .A1(n105486), .A2(n81259), .B1(n104938), .B2(n108980), 
        .ZN(n95679) );
  OAI21_X1 U82410 ( .B1(n106260), .B2(n95652), .A(n95680), .ZN(
        \DLX_Datapath/RegisterFile/N25617 ) );
  AOI22_X1 U82411 ( .A1(n105487), .A2(n94717), .B1(n104939), .B2(n109328), 
        .ZN(n95680) );
  OAI21_X1 U82412 ( .B1(n81509), .B2(n105488), .A(n95681), .ZN(
        \DLX_Datapath/RegisterFile/N25616 ) );
  AOI22_X1 U82413 ( .A1(n105486), .A2(n94719), .B1(n104940), .B2(n109210), 
        .ZN(n95681) );
  OAI21_X1 U82414 ( .B1(n81501), .B2(n105488), .A(n95682), .ZN(
        \DLX_Datapath/RegisterFile/N25615 ) );
  AOI22_X1 U82415 ( .A1(n105487), .A2(n94721), .B1(n104939), .B2(n109102), 
        .ZN(n95682) );
  OAI21_X1 U82416 ( .B1(n81415), .B2(n105488), .A(n95683), .ZN(
        \DLX_Datapath/RegisterFile/N25614 ) );
  AOI22_X1 U82417 ( .A1(n105486), .A2(n94723), .B1(n104938), .B2(n108637), 
        .ZN(n95683) );
  OAI21_X1 U82418 ( .B1(n81498), .B2(n105488), .A(n95684), .ZN(
        \DLX_Datapath/RegisterFile/N25613 ) );
  AOI22_X1 U82419 ( .A1(n105487), .A2(n94725), .B1(n104939), .B2(n108864), 
        .ZN(n95684) );
  OAI21_X1 U82420 ( .B1(n105217), .B2(n105488), .A(n95685), .ZN(
        \DLX_Datapath/RegisterFile/N25612 ) );
  AOI22_X1 U82421 ( .A1(n105487), .A2(n94727), .B1(n104938), .B2(n108752), 
        .ZN(n95685) );
  OAI21_X1 U82422 ( .B1(n106266), .B2(n105488), .A(n95686), .ZN(
        \DLX_Datapath/RegisterFile/N25611 ) );
  AOI22_X1 U82423 ( .A1(n105486), .A2(n94729), .B1(n104940), .B2(n107292), 
        .ZN(n95686) );
  AOI21_X1 U82424 ( .B1(n95687), .B2(n105602), .A(n104703), .ZN(n95655) );
  OAI21_X1 U82425 ( .B1(n95555), .B2(n95131), .A(n107022), .ZN(n95687) );
  NOR2_X1 U82426 ( .A1(n95689), .A2(n95555), .ZN(n95654) );
  OR2_X1 U82427 ( .A1(n95688), .A2(n95131), .ZN(n95689) );
  NOR2_X1 U82428 ( .A1(n95652), .A2(n105089), .ZN(n95688) );
  NAND2_X1 U82429 ( .A1(n105134), .A2(n94505), .ZN(n95652) );
  OAI21_X1 U82430 ( .B1(n106146), .B2(n105484), .A(n95691), .ZN(
        \DLX_Datapath/RegisterFile/N25610 ) );
  AOI22_X1 U82431 ( .A1(n104969), .A2(n107860), .B1(n105483), .B2(n81360), 
        .ZN(n95691) );
  OAI21_X1 U82432 ( .B1(n105969), .B2(n105484), .A(n95694), .ZN(
        \DLX_Datapath/RegisterFile/N25609 ) );
  AOI22_X1 U82433 ( .A1(n104970), .A2(n107957), .B1(n105482), .B2(n94511), 
        .ZN(n95694) );
  OAI21_X1 U82434 ( .B1(n106135), .B2(n105484), .A(n95695), .ZN(
        \DLX_Datapath/RegisterFile/N25608 ) );
  AOI22_X1 U82435 ( .A1(n104969), .A2(n107219), .B1(n105482), .B2(n81539), 
        .ZN(n95695) );
  OAI21_X1 U82436 ( .B1(n81299), .B2(n105484), .A(n95696), .ZN(
        \DLX_Datapath/RegisterFile/N25607 ) );
  AOI22_X1 U82437 ( .A1(n104970), .A2(n107757), .B1(n105483), .B2(n81301), 
        .ZN(n95696) );
  OAI21_X1 U82438 ( .B1(n106203), .B2(n105484), .A(n95697), .ZN(
        \DLX_Datapath/RegisterFile/N25606 ) );
  AOI22_X1 U82439 ( .A1(n104971), .A2(n110660), .B1(n105482), .B2(n81308), 
        .ZN(n95697) );
  OAI21_X1 U82440 ( .B1(n81408), .B2(n105484), .A(n95698), .ZN(
        \DLX_Datapath/RegisterFile/N25605 ) );
  AOI22_X1 U82441 ( .A1(n104970), .A2(n108059), .B1(n105483), .B2(n94516), 
        .ZN(n95698) );
  OAI21_X1 U82442 ( .B1(n106254), .B2(n105484), .A(n95699), .ZN(
        \DLX_Datapath/RegisterFile/N25604 ) );
  AOI22_X1 U82443 ( .A1(n104969), .A2(n110757), .B1(n105483), .B2(n81272), 
        .ZN(n95699) );
  OAI21_X1 U82444 ( .B1(n81629), .B2(n105484), .A(n95700), .ZN(
        \DLX_Datapath/RegisterFile/N25603 ) );
  AOI22_X1 U82445 ( .A1(n104971), .A2(n110858), .B1(n105482), .B2(n94519), 
        .ZN(n95700) );
  OAI21_X1 U82446 ( .B1(n106331), .B2(n105484), .A(n95701), .ZN(
        \DLX_Datapath/RegisterFile/N25602 ) );
  AOI22_X1 U82447 ( .A1(n104970), .A2(n110453), .B1(n105482), .B2(n80192), 
        .ZN(n95701) );
  OAI21_X1 U82448 ( .B1(n106190), .B2(n105484), .A(n95702), .ZN(
        \DLX_Datapath/RegisterFile/N25601 ) );
  AOI22_X1 U82449 ( .A1(n104969), .A2(n110235), .B1(n105481), .B2(n81474), 
        .ZN(n95702) );
  OAI21_X1 U82450 ( .B1(n106130), .B2(n105484), .A(n95703), .ZN(
        \DLX_Datapath/RegisterFile/N25600 ) );
  AOI22_X1 U82451 ( .A1(n104970), .A2(n110552), .B1(n105481), .B2(n94523), 
        .ZN(n95703) );
  OAI21_X1 U82452 ( .B1(n106187), .B2(n105484), .A(n95704), .ZN(
        \DLX_Datapath/RegisterFile/N25599 ) );
  AOI22_X1 U82453 ( .A1(n104971), .A2(n110343), .B1(n105481), .B2(n106061), 
        .ZN(n95704) );
  OAI21_X1 U82454 ( .B1(n106163), .B2(n105484), .A(n95705), .ZN(
        \DLX_Datapath/RegisterFile/N25598 ) );
  AOI22_X1 U82455 ( .A1(n104971), .A2(n110018), .B1(n105481), .B2(n81347), 
        .ZN(n95705) );
  OAI21_X1 U82456 ( .B1(n106103), .B2(n105484), .A(n95706), .ZN(
        \DLX_Datapath/RegisterFile/N25597 ) );
  AOI22_X1 U82457 ( .A1(n104969), .A2(n110125), .B1(n105481), .B2(n94527), 
        .ZN(n95706) );
  OAI21_X1 U82458 ( .B1(n81294), .B2(n105484), .A(n95707), .ZN(
        \DLX_Datapath/RegisterFile/N25596 ) );
  AOI22_X1 U82459 ( .A1(n104969), .A2(n109909), .B1(n105481), .B2(n81297), 
        .ZN(n95707) );
  OAI21_X1 U82460 ( .B1(n106110), .B2(n105484), .A(n95708), .ZN(
        \DLX_Datapath/RegisterFile/N25595 ) );
  AOI22_X1 U82461 ( .A1(n104970), .A2(n109791), .B1(n105483), .B2(n94530), 
        .ZN(n95708) );
  OAI21_X1 U82462 ( .B1(n106230), .B2(n105484), .A(n95709), .ZN(
        \DLX_Datapath/RegisterFile/N25594 ) );
  AOI22_X1 U82463 ( .A1(n104971), .A2(n108165), .B1(n105481), .B2(n81286), 
        .ZN(n95709) );
  OAI21_X1 U82464 ( .B1(n106170), .B2(n105484), .A(n95710), .ZN(
        \DLX_Datapath/RegisterFile/N25593 ) );
  AOI22_X1 U82465 ( .A1(n104970), .A2(n108288), .B1(n105481), .B2(n106168), 
        .ZN(n95710) );
  OAI21_X1 U82466 ( .B1(n81281), .B2(n105484), .A(n95711), .ZN(
        \DLX_Datapath/RegisterFile/N25592 ) );
  AOI22_X1 U82467 ( .A1(n104969), .A2(n108399), .B1(n105481), .B2(n81283), 
        .ZN(n95711) );
  OAI21_X1 U82468 ( .B1(n106069), .B2(n105484), .A(n95712), .ZN(
        \DLX_Datapath/RegisterFile/N25591 ) );
  AOI22_X1 U82469 ( .A1(n104970), .A2(n107637), .B1(n105481), .B2(n81453), 
        .ZN(n95712) );
  OAI21_X1 U82470 ( .B1(n106197), .B2(n105484), .A(n95713), .ZN(
        \DLX_Datapath/RegisterFile/N25590 ) );
  AOI22_X1 U82471 ( .A1(n104971), .A2(n109555), .B1(n105482), .B2(n94536), 
        .ZN(n95713) );
  OAI21_X1 U82472 ( .B1(n106244), .B2(n95690), .A(n95714), .ZN(
        \DLX_Datapath/RegisterFile/N25589 ) );
  AOI22_X1 U82473 ( .A1(n104971), .A2(n108516), .B1(n105483), .B2(n106241), 
        .ZN(n95714) );
  OAI21_X1 U82474 ( .B1(n81349), .B2(n105484), .A(n95715), .ZN(
        \DLX_Datapath/RegisterFile/N25588 ) );
  AOI22_X1 U82475 ( .A1(n104971), .A2(n109660), .B1(n105482), .B2(n81351), 
        .ZN(n95715) );
  OAI21_X1 U82476 ( .B1(n106113), .B2(n95690), .A(n95716), .ZN(
        \DLX_Datapath/RegisterFile/N25587 ) );
  AOI22_X1 U82477 ( .A1(n104969), .A2(n109444), .B1(n105483), .B2(n106020), 
        .ZN(n95716) );
  OAI21_X1 U82478 ( .B1(n81588), .B2(n95690), .A(n95717), .ZN(
        \DLX_Datapath/RegisterFile/N25586 ) );
  AOI22_X1 U82479 ( .A1(n104969), .A2(n108981), .B1(n105482), .B2(n94541), 
        .ZN(n95717) );
  OAI21_X1 U82480 ( .B1(n81267), .B2(n105484), .A(n95718), .ZN(
        \DLX_Datapath/RegisterFile/N25585 ) );
  AOI22_X1 U82481 ( .A1(n104970), .A2(n109329), .B1(n105482), .B2(n81269), 
        .ZN(n95718) );
  OAI21_X1 U82482 ( .B1(n106044), .B2(n95690), .A(n95719), .ZN(
        \DLX_Datapath/RegisterFile/N25584 ) );
  AOI22_X1 U82483 ( .A1(n104971), .A2(n109211), .B1(n105483), .B2(n105624), 
        .ZN(n95719) );
  OAI21_X1 U82484 ( .B1(n106048), .B2(n95690), .A(n95720), .ZN(
        \DLX_Datapath/RegisterFile/N25583 ) );
  AOI22_X1 U82485 ( .A1(n104970), .A2(n109103), .B1(n105482), .B2(n94546), 
        .ZN(n95720) );
  OAI21_X1 U82486 ( .B1(n81415), .B2(n95690), .A(n95721), .ZN(
        \DLX_Datapath/RegisterFile/N25582 ) );
  AOI22_X1 U82487 ( .A1(n104969), .A2(n108638), .B1(n105483), .B2(n94548), 
        .ZN(n95721) );
  OAI21_X1 U82488 ( .B1(n106053), .B2(n95690), .A(n95722), .ZN(
        \DLX_Datapath/RegisterFile/N25581 ) );
  AOI22_X1 U82489 ( .A1(n104970), .A2(n108865), .B1(n105483), .B2(n81783), 
        .ZN(n95722) );
  OAI21_X1 U82490 ( .B1(n105216), .B2(n95690), .A(n95723), .ZN(
        \DLX_Datapath/RegisterFile/N25580 ) );
  AOI22_X1 U82491 ( .A1(n104969), .A2(n108753), .B1(n105483), .B2(n80188), 
        .ZN(n95723) );
  OAI21_X1 U82492 ( .B1(n106266), .B2(n95690), .A(n95724), .ZN(
        \DLX_Datapath/RegisterFile/N25579 ) );
  AOI22_X1 U82493 ( .A1(n104971), .A2(n107293), .B1(n105482), .B2(n81265), 
        .ZN(n95724) );
  NOR2_X1 U82496 ( .A1(n95690), .A2(n105094), .ZN(n95726) );
  NAND2_X1 U82497 ( .A1(n105133), .A2(n94555), .ZN(n95690) );
  OAI21_X1 U82498 ( .B1(n106146), .B2(n105480), .A(n95728), .ZN(
        \DLX_Datapath/RegisterFile/N25578 ) );
  AOI22_X1 U82499 ( .A1(n104947), .A2(n94559), .B1(n104956), .B2(n107861), 
        .ZN(n95728) );
  OAI21_X1 U82500 ( .B1(n105969), .B2(n105480), .A(n95731), .ZN(
        \DLX_Datapath/RegisterFile/N25577 ) );
  AOI22_X1 U82501 ( .A1(n104948), .A2(n94562), .B1(n104957), .B2(n107958), 
        .ZN(n95731) );
  OAI21_X1 U82502 ( .B1(n106135), .B2(n105480), .A(n95732), .ZN(
        \DLX_Datapath/RegisterFile/N25576 ) );
  AOI22_X1 U82503 ( .A1(n104947), .A2(n94564), .B1(n104956), .B2(n107220), 
        .ZN(n95732) );
  OAI21_X1 U82504 ( .B1(n81299), .B2(n105480), .A(n95733), .ZN(
        \DLX_Datapath/RegisterFile/N25575 ) );
  AOI22_X1 U82505 ( .A1(n104949), .A2(n94566), .B1(n104958), .B2(n107758), 
        .ZN(n95733) );
  OAI21_X1 U82506 ( .B1(n106203), .B2(n105480), .A(n95734), .ZN(
        \DLX_Datapath/RegisterFile/N25574 ) );
  AOI22_X1 U82507 ( .A1(n104947), .A2(n94568), .B1(n104956), .B2(n110661), 
        .ZN(n95734) );
  OAI21_X1 U82508 ( .B1(n81408), .B2(n105480), .A(n95735), .ZN(
        \DLX_Datapath/RegisterFile/N25573 ) );
  AOI22_X1 U82509 ( .A1(n104948), .A2(n94570), .B1(n104957), .B2(n108060), 
        .ZN(n95735) );
  OAI21_X1 U82510 ( .B1(n106255), .B2(n105480), .A(n95736), .ZN(
        \DLX_Datapath/RegisterFile/N25572 ) );
  AOI22_X1 U82511 ( .A1(n104948), .A2(n94572), .B1(n104957), .B2(n110758), 
        .ZN(n95736) );
  OAI21_X1 U82512 ( .B1(n81629), .B2(n105480), .A(n95737), .ZN(
        \DLX_Datapath/RegisterFile/N25571 ) );
  AOI22_X1 U82513 ( .A1(n104949), .A2(n94574), .B1(n104958), .B2(n110859), 
        .ZN(n95737) );
  OAI21_X1 U82514 ( .B1(n106330), .B2(n105480), .A(n95738), .ZN(
        \DLX_Datapath/RegisterFile/N25570 ) );
  AOI22_X1 U82515 ( .A1(n104948), .A2(n94576), .B1(n104957), .B2(n110454), 
        .ZN(n95738) );
  OAI21_X1 U82516 ( .B1(n106191), .B2(n105480), .A(n95739), .ZN(
        \DLX_Datapath/RegisterFile/N25569 ) );
  AOI22_X1 U82517 ( .A1(n104947), .A2(n94578), .B1(n104956), .B2(n110236), 
        .ZN(n95739) );
  OAI21_X1 U82518 ( .B1(n106128), .B2(n105480), .A(n95740), .ZN(
        \DLX_Datapath/RegisterFile/N25568 ) );
  AOI22_X1 U82519 ( .A1(n104948), .A2(n94580), .B1(n104957), .B2(n110553), 
        .ZN(n95740) );
  OAI21_X1 U82520 ( .B1(n106187), .B2(n105480), .A(n95741), .ZN(
        \DLX_Datapath/RegisterFile/N25567 ) );
  AOI22_X1 U82521 ( .A1(n104949), .A2(n94582), .B1(n104958), .B2(n110344), 
        .ZN(n95741) );
  OAI21_X1 U82522 ( .B1(n106163), .B2(n105480), .A(n95742), .ZN(
        \DLX_Datapath/RegisterFile/N25566 ) );
  AOI22_X1 U82523 ( .A1(n104949), .A2(n94584), .B1(n104958), .B2(n110019), 
        .ZN(n95742) );
  OAI21_X1 U82524 ( .B1(n81403), .B2(n105480), .A(n95743), .ZN(
        \DLX_Datapath/RegisterFile/N25565 ) );
  AOI22_X1 U82525 ( .A1(n104947), .A2(n94586), .B1(n104956), .B2(n110126), 
        .ZN(n95743) );
  OAI21_X1 U82526 ( .B1(n81294), .B2(n105480), .A(n95744), .ZN(
        \DLX_Datapath/RegisterFile/N25564 ) );
  AOI22_X1 U82527 ( .A1(n104947), .A2(n94588), .B1(n104956), .B2(n109910), 
        .ZN(n95744) );
  OAI21_X1 U82528 ( .B1(n106108), .B2(n105480), .A(n95745), .ZN(
        \DLX_Datapath/RegisterFile/N25563 ) );
  AOI22_X1 U82529 ( .A1(n104948), .A2(n94590), .B1(n104957), .B2(n109792), 
        .ZN(n95745) );
  OAI21_X1 U82530 ( .B1(n106230), .B2(n105480), .A(n95746), .ZN(
        \DLX_Datapath/RegisterFile/N25562 ) );
  AOI22_X1 U82531 ( .A1(n104949), .A2(n94592), .B1(n104958), .B2(n108166), 
        .ZN(n95746) );
  OAI21_X1 U82532 ( .B1(n81340), .B2(n105480), .A(n95747), .ZN(
        \DLX_Datapath/RegisterFile/N25561 ) );
  AOI22_X1 U82533 ( .A1(n104948), .A2(n94594), .B1(n104957), .B2(n108289), 
        .ZN(n95747) );
  OAI21_X1 U82534 ( .B1(n106237), .B2(n105480), .A(n95748), .ZN(
        \DLX_Datapath/RegisterFile/N25560 ) );
  AOI22_X1 U82535 ( .A1(n104947), .A2(n94596), .B1(n104956), .B2(n108400), 
        .ZN(n95748) );
  OAI21_X1 U82536 ( .B1(n106070), .B2(n105480), .A(n95749), .ZN(
        \DLX_Datapath/RegisterFile/N25559 ) );
  AOI22_X1 U82537 ( .A1(n104948), .A2(n94598), .B1(n104957), .B2(n107638), 
        .ZN(n95749) );
  OAI21_X1 U82538 ( .B1(n106200), .B2(n105480), .A(n95750), .ZN(
        \DLX_Datapath/RegisterFile/N25558 ) );
  AOI22_X1 U82539 ( .A1(n104949), .A2(n94600), .B1(n104958), .B2(n109556), 
        .ZN(n95750) );
  OAI21_X1 U82540 ( .B1(n106244), .B2(n95727), .A(n95751), .ZN(
        \DLX_Datapath/RegisterFile/N25557 ) );
  AOI22_X1 U82541 ( .A1(n104949), .A2(n94602), .B1(n104958), .B2(n108517), 
        .ZN(n95751) );
  OAI21_X1 U82542 ( .B1(n81349), .B2(n95727), .A(n95752), .ZN(
        \DLX_Datapath/RegisterFile/N25556 ) );
  AOI22_X1 U82543 ( .A1(n104949), .A2(n94604), .B1(n104958), .B2(n109661), 
        .ZN(n95752) );
  OAI21_X1 U82544 ( .B1(n106113), .B2(n95727), .A(n95753), .ZN(
        \DLX_Datapath/RegisterFile/N25555 ) );
  AOI22_X1 U82545 ( .A1(n104947), .A2(n94606), .B1(n104956), .B2(n109445), 
        .ZN(n95753) );
  OAI21_X1 U82546 ( .B1(n81588), .B2(n95727), .A(n95754), .ZN(
        \DLX_Datapath/RegisterFile/N25554 ) );
  AOI22_X1 U82547 ( .A1(n104949), .A2(n94608), .B1(n104958), .B2(n108982), 
        .ZN(n95754) );
  OAI21_X1 U82548 ( .B1(n81267), .B2(n105480), .A(n95755), .ZN(
        \DLX_Datapath/RegisterFile/N25553 ) );
  AOI22_X1 U82549 ( .A1(n104948), .A2(n94610), .B1(n104957), .B2(n109330), 
        .ZN(n95755) );
  OAI21_X1 U82550 ( .B1(n106043), .B2(n95727), .A(n95756), .ZN(
        \DLX_Datapath/RegisterFile/N25552 ) );
  AOI22_X1 U82551 ( .A1(n104949), .A2(n94612), .B1(n104958), .B2(n109212), 
        .ZN(n95756) );
  OAI21_X1 U82552 ( .B1(n106048), .B2(n95727), .A(n95757), .ZN(
        \DLX_Datapath/RegisterFile/N25551 ) );
  AOI22_X1 U82553 ( .A1(n104947), .A2(n94614), .B1(n104956), .B2(n109104), 
        .ZN(n95757) );
  OAI21_X1 U82554 ( .B1(n81415), .B2(n95727), .A(n95758), .ZN(
        \DLX_Datapath/RegisterFile/N25550 ) );
  AOI22_X1 U82555 ( .A1(n104947), .A2(n94616), .B1(n104956), .B2(n108639), 
        .ZN(n95758) );
  OAI21_X1 U82556 ( .B1(n106056), .B2(n95727), .A(n95759), .ZN(
        \DLX_Datapath/RegisterFile/N25549 ) );
  AOI22_X1 U82557 ( .A1(n104948), .A2(n94618), .B1(n104957), .B2(n108866), 
        .ZN(n95759) );
  OAI21_X1 U82558 ( .B1(n105215), .B2(n95727), .A(n95760), .ZN(
        \DLX_Datapath/RegisterFile/N25548 ) );
  AOI22_X1 U82559 ( .A1(n104947), .A2(n94620), .B1(n104956), .B2(n108754), 
        .ZN(n95760) );
  OAI21_X1 U82560 ( .B1(n81262), .B2(n105480), .A(n95761), .ZN(
        \DLX_Datapath/RegisterFile/N25547 ) );
  AOI22_X1 U82561 ( .A1(n104948), .A2(n94622), .B1(n104957), .B2(n107294), 
        .ZN(n95761) );
  NOR2_X1 U82563 ( .A1(n95725), .A2(n95762), .ZN(n95729) );
  NOR2_X1 U82564 ( .A1(n95727), .A2(n105089), .ZN(n95762) );
  NAND2_X1 U82565 ( .A1(n94625), .A2(n105133), .ZN(n95727) );
  OAI21_X1 U82566 ( .B1(n106146), .B2(n105479), .A(n95765), .ZN(
        \DLX_Datapath/RegisterFile/N25546 ) );
  AOI22_X1 U82567 ( .A1(n105478), .A2(n107862), .B1(n104935), .B2(n81521), 
        .ZN(n95765) );
  OAI21_X1 U82568 ( .B1(n105969), .B2(n105479), .A(n95768), .ZN(
        \DLX_Datapath/RegisterFile/N25545 ) );
  AOI22_X1 U82569 ( .A1(n105477), .A2(n107959), .B1(n104936), .B2(n81653), 
        .ZN(n95768) );
  OAI21_X1 U82570 ( .B1(n106135), .B2(n105479), .A(n95769), .ZN(
        \DLX_Datapath/RegisterFile/N25544 ) );
  AOI22_X1 U82571 ( .A1(n105478), .A2(n107221), .B1(n104935), .B2(n81380), 
        .ZN(n95769) );
  OAI21_X1 U82572 ( .B1(n81299), .B2(n105479), .A(n95770), .ZN(
        \DLX_Datapath/RegisterFile/N25543 ) );
  AOI22_X1 U82573 ( .A1(n105477), .A2(n107759), .B1(n104937), .B2(n81377), 
        .ZN(n95770) );
  OAI21_X1 U82574 ( .B1(n106203), .B2(n105479), .A(n95771), .ZN(
        \DLX_Datapath/RegisterFile/N25542 ) );
  AOI22_X1 U82575 ( .A1(n105478), .A2(n110662), .B1(n104935), .B2(n81428), 
        .ZN(n95771) );
  OAI21_X1 U82576 ( .B1(n81408), .B2(n105479), .A(n95772), .ZN(
        \DLX_Datapath/RegisterFile/N25541 ) );
  AOI22_X1 U82577 ( .A1(n105477), .A2(n108061), .B1(n104936), .B2(n81410), 
        .ZN(n95772) );
  OAI21_X1 U82578 ( .B1(n106257), .B2(n105479), .A(n95773), .ZN(
        \DLX_Datapath/RegisterFile/N25540 ) );
  AOI22_X1 U82579 ( .A1(n105477), .A2(n110759), .B1(n104937), .B2(n81700), 
        .ZN(n95773) );
  OAI21_X1 U82580 ( .B1(n81629), .B2(n105479), .A(n95774), .ZN(
        \DLX_Datapath/RegisterFile/N25539 ) );
  AOI22_X1 U82581 ( .A1(n105478), .A2(n110860), .B1(n104936), .B2(n81632), 
        .ZN(n95774) );
  OAI21_X1 U82582 ( .B1(n106333), .B2(n105479), .A(n95775), .ZN(
        \DLX_Datapath/RegisterFile/N25538 ) );
  AOI22_X1 U82583 ( .A1(n105477), .A2(n110455), .B1(n104936), .B2(n81414), 
        .ZN(n95775) );
  OAI21_X1 U82584 ( .B1(n106192), .B2(n105479), .A(n95776), .ZN(
        \DLX_Datapath/RegisterFile/N25537 ) );
  AOI22_X1 U82585 ( .A1(n105476), .A2(n110237), .B1(n104935), .B2(n81317), 
        .ZN(n95776) );
  OAI21_X1 U82586 ( .B1(n106128), .B2(n105479), .A(n95777), .ZN(
        \DLX_Datapath/RegisterFile/N25536 ) );
  AOI22_X1 U82587 ( .A1(n105476), .A2(n110554), .B1(n104936), .B2(n81386), 
        .ZN(n95777) );
  OAI21_X1 U82588 ( .B1(n106188), .B2(n105479), .A(n95778), .ZN(
        \DLX_Datapath/RegisterFile/N25535 ) );
  AOI22_X1 U82589 ( .A1(n105476), .A2(n110345), .B1(n104937), .B2(n81320), 
        .ZN(n95778) );
  OAI21_X1 U82590 ( .B1(n106162), .B2(n105479), .A(n95779), .ZN(
        \DLX_Datapath/RegisterFile/N25534 ) );
  AOI22_X1 U82591 ( .A1(n105476), .A2(n110020), .B1(n104937), .B2(n81604), 
        .ZN(n95779) );
  OAI21_X1 U82592 ( .B1(n81403), .B2(n105479), .A(n95780), .ZN(
        \DLX_Datapath/RegisterFile/N25533 ) );
  AOI22_X1 U82593 ( .A1(n105476), .A2(n110127), .B1(n104935), .B2(n81405), 
        .ZN(n95780) );
  OAI21_X1 U82594 ( .B1(n106219), .B2(n105479), .A(n95781), .ZN(
        \DLX_Datapath/RegisterFile/N25532 ) );
  AOI22_X1 U82595 ( .A1(n105476), .A2(n109911), .B1(n104935), .B2(n81402), 
        .ZN(n95781) );
  OAI21_X1 U82596 ( .B1(n106111), .B2(n105479), .A(n95782), .ZN(
        \DLX_Datapath/RegisterFile/N25531 ) );
  AOI22_X1 U82597 ( .A1(n105476), .A2(n109793), .B1(n104936), .B2(n81400), 
        .ZN(n95782) );
  OAI21_X1 U82598 ( .B1(n106230), .B2(n105479), .A(n95783), .ZN(
        \DLX_Datapath/RegisterFile/N25530 ) );
  AOI22_X1 U82599 ( .A1(n105476), .A2(n108167), .B1(n104937), .B2(n81332), 
        .ZN(n95783) );
  OAI21_X1 U82600 ( .B1(n106173), .B2(n105479), .A(n95784), .ZN(
        \DLX_Datapath/RegisterFile/N25529 ) );
  AOI22_X1 U82601 ( .A1(n105476), .A2(n108290), .B1(n104936), .B2(n81373), 
        .ZN(n95784) );
  OAI21_X1 U82602 ( .B1(n81281), .B2(n105479), .A(n95785), .ZN(
        \DLX_Datapath/RegisterFile/N25528 ) );
  AOI22_X1 U82603 ( .A1(n105476), .A2(n108401), .B1(n104935), .B2(n81322), 
        .ZN(n95785) );
  OAI21_X1 U82604 ( .B1(n106071), .B2(n105479), .A(n95786), .ZN(
        \DLX_Datapath/RegisterFile/N25527 ) );
  AOI22_X1 U82605 ( .A1(n105476), .A2(n107639), .B1(n104936), .B2(n81506), 
        .ZN(n95786) );
  OAI21_X1 U82606 ( .B1(n106199), .B2(n105479), .A(n95787), .ZN(
        \DLX_Datapath/RegisterFile/N25526 ) );
  AOI22_X1 U82607 ( .A1(n105477), .A2(n109557), .B1(n104937), .B2(n81313), 
        .ZN(n95787) );
  OAI21_X1 U82608 ( .B1(n106244), .B2(n95764), .A(n95788), .ZN(
        \DLX_Datapath/RegisterFile/N25525 ) );
  AOI22_X1 U82609 ( .A1(n105478), .A2(n108518), .B1(n104937), .B2(n81330), 
        .ZN(n95788) );
  OAI21_X1 U82610 ( .B1(n81349), .B2(n95764), .A(n95789), .ZN(
        \DLX_Datapath/RegisterFile/N25524 ) );
  AOI22_X1 U82611 ( .A1(n105477), .A2(n109662), .B1(n104937), .B2(n81425), 
        .ZN(n95789) );
  OAI21_X1 U82612 ( .B1(n106113), .B2(n95764), .A(n95790), .ZN(
        \DLX_Datapath/RegisterFile/N25523 ) );
  AOI22_X1 U82613 ( .A1(n105478), .A2(n109446), .B1(n104935), .B2(n81396), 
        .ZN(n95790) );
  OAI21_X1 U82614 ( .B1(n81588), .B2(n95764), .A(n95791), .ZN(
        \DLX_Datapath/RegisterFile/N25522 ) );
  AOI22_X1 U82615 ( .A1(n105477), .A2(n108983), .B1(n104935), .B2(n81590), 
        .ZN(n95791) );
  OAI21_X1 U82616 ( .B1(n81267), .B2(n105479), .A(n95792), .ZN(
        \DLX_Datapath/RegisterFile/N25521 ) );
  AOI22_X1 U82617 ( .A1(n105478), .A2(n109331), .B1(n104936), .B2(n81423), 
        .ZN(n95792) );
  OAI21_X1 U82618 ( .B1(n106046), .B2(n95764), .A(n95793), .ZN(
        \DLX_Datapath/RegisterFile/N25520 ) );
  AOI22_X1 U82619 ( .A1(n105477), .A2(n109213), .B1(n104937), .B2(n81511), 
        .ZN(n95793) );
  OAI21_X1 U82620 ( .B1(n106048), .B2(n95764), .A(n95794), .ZN(
        \DLX_Datapath/RegisterFile/N25519 ) );
  AOI22_X1 U82621 ( .A1(n105478), .A2(n109105), .B1(n104936), .B2(n81503), 
        .ZN(n95794) );
  OAI21_X1 U82622 ( .B1(n81415), .B2(n95764), .A(n95795), .ZN(
        \DLX_Datapath/RegisterFile/N25518 ) );
  AOI22_X1 U82623 ( .A1(n105477), .A2(n108640), .B1(n104935), .B2(n81417), 
        .ZN(n95795) );
  OAI21_X1 U82624 ( .B1(n106054), .B2(n95764), .A(n95796), .ZN(
        \DLX_Datapath/RegisterFile/N25517 ) );
  AOI22_X1 U82625 ( .A1(n105478), .A2(n108867), .B1(n104936), .B2(n81500), 
        .ZN(n95796) );
  OAI21_X1 U82626 ( .B1(n105217), .B2(n95764), .A(n95797), .ZN(
        \DLX_Datapath/RegisterFile/N25516 ) );
  AOI22_X1 U82627 ( .A1(n105478), .A2(n108755), .B1(n104935), .B2(n81335), 
        .ZN(n95797) );
  OAI21_X1 U82628 ( .B1(n81262), .B2(n105479), .A(n95798), .ZN(
        \DLX_Datapath/RegisterFile/N25515 ) );
  AOI22_X1 U82629 ( .A1(n105477), .A2(n107295), .B1(n104937), .B2(n81327), 
        .ZN(n95798) );
  AOI21_X1 U82632 ( .B1(n105199), .B2(n95725), .A(n94663), .ZN(n95763) );
  OR2_X1 U82633 ( .A1(n95517), .A2(n86230), .ZN(n95725) );
  NOR2_X1 U82634 ( .A1(n95764), .A2(n105090), .ZN(n95799) );
  NAND2_X1 U82635 ( .A1(n105134), .A2(n94664), .ZN(n95764) );
  OAI21_X1 U82636 ( .B1(n106146), .B2(n105475), .A(n95801), .ZN(
        \DLX_Datapath/RegisterFile/N25514 ) );
  AOI22_X1 U82637 ( .A1(n104840), .A2(n94667), .B1(n105473), .B2(n107863), 
        .ZN(n95801) );
  OAI21_X1 U82638 ( .B1(n105968), .B2(n105474), .A(n95804), .ZN(
        \DLX_Datapath/RegisterFile/N25513 ) );
  AOI22_X1 U82639 ( .A1(n104840), .A2(n94670), .B1(n95803), .B2(n107960), .ZN(
        n95804) );
  OAI21_X1 U82640 ( .B1(n106135), .B2(n105475), .A(n95805), .ZN(
        \DLX_Datapath/RegisterFile/N25512 ) );
  AOI22_X1 U82641 ( .A1(n104840), .A2(n94672), .B1(n105473), .B2(n107222), 
        .ZN(n95805) );
  OAI21_X1 U82642 ( .B1(n106208), .B2(n105475), .A(n95806), .ZN(
        \DLX_Datapath/RegisterFile/N25511 ) );
  AOI22_X1 U82643 ( .A1(n104840), .A2(n94674), .B1(n95803), .B2(n107760), .ZN(
        n95806) );
  OAI21_X1 U82644 ( .B1(n106203), .B2(n105474), .A(n95807), .ZN(
        \DLX_Datapath/RegisterFile/N25510 ) );
  AOI22_X1 U82645 ( .A1(n104841), .A2(n94676), .B1(n105473), .B2(n110663), 
        .ZN(n95807) );
  OAI21_X1 U82646 ( .B1(n81408), .B2(n105474), .A(n95808), .ZN(
        \DLX_Datapath/RegisterFile/N25509 ) );
  AOI22_X1 U82647 ( .A1(n104842), .A2(n94678), .B1(n105472), .B2(n108062), 
        .ZN(n95808) );
  OAI21_X1 U82648 ( .B1(n106255), .B2(n105475), .A(n95809), .ZN(
        \DLX_Datapath/RegisterFile/N25508 ) );
  AOI22_X1 U82649 ( .A1(n104841), .A2(n94680), .B1(n105473), .B2(n110760), 
        .ZN(n95809) );
  OAI21_X1 U82650 ( .B1(n105990), .B2(n105474), .A(n95810), .ZN(
        \DLX_Datapath/RegisterFile/N25507 ) );
  AOI22_X1 U82651 ( .A1(n104842), .A2(n94682), .B1(n95803), .B2(n110861), .ZN(
        n95810) );
  OAI21_X1 U82652 ( .B1(n80190), .B2(n105474), .A(n95811), .ZN(
        \DLX_Datapath/RegisterFile/N25506 ) );
  AOI22_X1 U82653 ( .A1(n104842), .A2(n94684), .B1(n95803), .B2(n110456), .ZN(
        n95811) );
  OAI21_X1 U82654 ( .B1(n81315), .B2(n105474), .A(n95812), .ZN(
        \DLX_Datapath/RegisterFile/N25505 ) );
  AOI22_X1 U82655 ( .A1(n104842), .A2(n94686), .B1(n105472), .B2(n110238), 
        .ZN(n95812) );
  OAI21_X1 U82656 ( .B1(n106128), .B2(n105475), .A(n95813), .ZN(
        \DLX_Datapath/RegisterFile/N25504 ) );
  AOI22_X1 U82657 ( .A1(n104840), .A2(n94688), .B1(n105472), .B2(n110555), 
        .ZN(n95813) );
  OAI21_X1 U82658 ( .B1(n81318), .B2(n105475), .A(n95814), .ZN(
        \DLX_Datapath/RegisterFile/N25503 ) );
  AOI22_X1 U82659 ( .A1(n104842), .A2(n94690), .B1(n105472), .B2(n110346), 
        .ZN(n95814) );
  OAI21_X1 U82660 ( .B1(n106165), .B2(n105475), .A(n95815), .ZN(
        \DLX_Datapath/RegisterFile/N25502 ) );
  AOI22_X1 U82661 ( .A1(n104840), .A2(n94692), .B1(n105472), .B2(n110021), 
        .ZN(n95815) );
  OAI21_X1 U82662 ( .B1(n81403), .B2(n105474), .A(n95816), .ZN(
        \DLX_Datapath/RegisterFile/N25501 ) );
  AOI22_X1 U82663 ( .A1(n104841), .A2(n94694), .B1(n105472), .B2(n110128), 
        .ZN(n95816) );
  OAI21_X1 U82664 ( .B1(n106218), .B2(n105474), .A(n95817), .ZN(
        \DLX_Datapath/RegisterFile/N25500 ) );
  AOI22_X1 U82665 ( .A1(n104842), .A2(n94696), .B1(n105472), .B2(n109912), 
        .ZN(n95817) );
  OAI21_X1 U82666 ( .B1(n106108), .B2(n105475), .A(n95818), .ZN(
        \DLX_Datapath/RegisterFile/N25499 ) );
  AOI22_X1 U82667 ( .A1(n104841), .A2(n94698), .B1(n105472), .B2(n109794), 
        .ZN(n95818) );
  OAI21_X1 U82668 ( .B1(n106231), .B2(n105475), .A(n95819), .ZN(
        \DLX_Datapath/RegisterFile/N25498 ) );
  AOI22_X1 U82669 ( .A1(n104842), .A2(n94700), .B1(n105472), .B2(n108168), 
        .ZN(n95819) );
  OAI21_X1 U82670 ( .B1(n106171), .B2(n105474), .A(n95820), .ZN(
        \DLX_Datapath/RegisterFile/N25497 ) );
  AOI22_X1 U82671 ( .A1(n104842), .A2(n94702), .B1(n105472), .B2(n108291), 
        .ZN(n95820) );
  OAI21_X1 U82672 ( .B1(n106238), .B2(n105474), .A(n95821), .ZN(
        \DLX_Datapath/RegisterFile/N25496 ) );
  AOI22_X1 U82673 ( .A1(n104840), .A2(n94704), .B1(n105472), .B2(n108402), 
        .ZN(n95821) );
  OAI21_X1 U82674 ( .B1(n81451), .B2(n105475), .A(n95822), .ZN(
        \DLX_Datapath/RegisterFile/N25495 ) );
  AOI22_X1 U82675 ( .A1(n104841), .A2(n94706), .B1(n105472), .B2(n107640), 
        .ZN(n95822) );
  OAI21_X1 U82676 ( .B1(n81310), .B2(n105474), .A(n95823), .ZN(
        \DLX_Datapath/RegisterFile/N25494 ) );
  AOI22_X1 U82677 ( .A1(n104840), .A2(n94708), .B1(n95803), .B2(n109558), .ZN(
        n95823) );
  OAI21_X1 U82678 ( .B1(n106244), .B2(n105475), .A(n95824), .ZN(
        \DLX_Datapath/RegisterFile/N25493 ) );
  AOI22_X1 U82679 ( .A1(n104841), .A2(n94710), .B1(n105473), .B2(n108519), 
        .ZN(n95824) );
  OAI21_X1 U82680 ( .B1(n81349), .B2(n105474), .A(n95825), .ZN(
        \DLX_Datapath/RegisterFile/N25492 ) );
  AOI22_X1 U82681 ( .A1(n104842), .A2(n94712), .B1(n105472), .B2(n109663), 
        .ZN(n95825) );
  OAI21_X1 U82682 ( .B1(n106113), .B2(n105475), .A(n95826), .ZN(
        \DLX_Datapath/RegisterFile/N25491 ) );
  AOI22_X1 U82683 ( .A1(n104840), .A2(n94714), .B1(n105473), .B2(n109447), 
        .ZN(n95826) );
  OAI21_X1 U82684 ( .B1(n106008), .B2(n105474), .A(n95827), .ZN(
        \DLX_Datapath/RegisterFile/N25490 ) );
  AOI22_X1 U82685 ( .A1(n104840), .A2(n81259), .B1(n105472), .B2(n108984), 
        .ZN(n95827) );
  OAI21_X1 U82686 ( .B1(n106259), .B2(n105474), .A(n95828), .ZN(
        \DLX_Datapath/RegisterFile/N25489 ) );
  AOI22_X1 U82687 ( .A1(n104840), .A2(n94717), .B1(n105473), .B2(n109332), 
        .ZN(n95828) );
  OAI21_X1 U82688 ( .B1(n106043), .B2(n105475), .A(n95829), .ZN(
        \DLX_Datapath/RegisterFile/N25488 ) );
  AOI22_X1 U82689 ( .A1(n104840), .A2(n94719), .B1(n95803), .B2(n109214), .ZN(
        n95829) );
  OAI21_X1 U82690 ( .B1(n106048), .B2(n105474), .A(n95830), .ZN(
        \DLX_Datapath/RegisterFile/N25487 ) );
  AOI22_X1 U82691 ( .A1(n104841), .A2(n94721), .B1(n105473), .B2(n109106), 
        .ZN(n95830) );
  OAI21_X1 U82692 ( .B1(n81415), .B2(n105475), .A(n95831), .ZN(
        \DLX_Datapath/RegisterFile/N25486 ) );
  AOI22_X1 U82693 ( .A1(n104842), .A2(n94723), .B1(n105473), .B2(n108641), 
        .ZN(n95831) );
  OAI21_X1 U82694 ( .B1(n81498), .B2(n105475), .A(n95832), .ZN(
        \DLX_Datapath/RegisterFile/N25485 ) );
  AOI22_X1 U82695 ( .A1(n104841), .A2(n94725), .B1(n105473), .B2(n108868), 
        .ZN(n95832) );
  OAI21_X1 U82696 ( .B1(n105216), .B2(n105475), .A(n95833), .ZN(
        \DLX_Datapath/RegisterFile/N25484 ) );
  AOI22_X1 U82697 ( .A1(n104841), .A2(n94727), .B1(n105473), .B2(n108756), 
        .ZN(n95833) );
  OAI21_X1 U82698 ( .B1(n106268), .B2(n105474), .A(n95834), .ZN(
        \DLX_Datapath/RegisterFile/N25483 ) );
  AOI22_X1 U82699 ( .A1(n104842), .A2(n94729), .B1(n95803), .B2(n107296), .ZN(
        n95834) );
  AOI21_X1 U82700 ( .B1(n95835), .B2(n105602), .A(n95836), .ZN(n95803) );
  OAI21_X1 U82701 ( .B1(n95555), .B2(n86230), .A(n105199), .ZN(n95835) );
  NOR2_X1 U82702 ( .A1(n95837), .A2(n95555), .ZN(n95802) );
  OR2_X1 U82703 ( .A1(n95836), .A2(n86230), .ZN(n95837) );
  NOR2_X1 U82704 ( .A1(n95800), .A2(n105091), .ZN(n95836) );
  NAND2_X1 U82705 ( .A1(n94734), .A2(n105134), .ZN(n95800) );
  OAI21_X1 U82706 ( .B1(n81358), .B2(n105471), .A(n95839), .ZN(
        \DLX_Datapath/RegisterFile/N25482 ) );
  AOI22_X1 U82707 ( .A1(n104816), .A2(n81360), .B1(n105469), .B2(n70303), .ZN(
        n95839) );
  OAI21_X1 U82708 ( .B1(n105969), .B2(n105471), .A(n95842), .ZN(
        \DLX_Datapath/RegisterFile/N25481 ) );
  AOI22_X1 U82709 ( .A1(n104817), .A2(n94511), .B1(n105469), .B2(n70445), .ZN(
        n95842) );
  OAI21_X1 U82710 ( .B1(n106135), .B2(n105471), .A(n95843), .ZN(
        \DLX_Datapath/RegisterFile/N25480 ) );
  AOI22_X1 U82711 ( .A1(n104816), .A2(n81539), .B1(n105469), .B2(n69498), .ZN(
        n95843) );
  OAI21_X1 U82712 ( .B1(n106208), .B2(n105471), .A(n95844), .ZN(
        \DLX_Datapath/RegisterFile/N25479 ) );
  AOI22_X1 U82713 ( .A1(n104817), .A2(n81301), .B1(n105469), .B2(n70159), .ZN(
        n95844) );
  OAI21_X1 U82714 ( .B1(n106203), .B2(n105471), .A(n95845), .ZN(
        \DLX_Datapath/RegisterFile/N25478 ) );
  AOI22_X1 U82715 ( .A1(n104816), .A2(n81308), .B1(n105469), .B2(n74005), .ZN(
        n95845) );
  OAI21_X1 U82716 ( .B1(n81408), .B2(n105471), .A(n95846), .ZN(
        \DLX_Datapath/RegisterFile/N25477 ) );
  AOI22_X1 U82717 ( .A1(n104818), .A2(n94516), .B1(n105469), .B2(n70592), .ZN(
        n95846) );
  OAI21_X1 U82718 ( .B1(n106256), .B2(n105471), .A(n95847), .ZN(
        \DLX_Datapath/RegisterFile/N25476 ) );
  AOI22_X1 U82719 ( .A1(n104816), .A2(n81272), .B1(n105469), .B2(n74146), .ZN(
        n95847) );
  OAI21_X1 U82720 ( .B1(n105992), .B2(n105471), .A(n95848), .ZN(
        \DLX_Datapath/RegisterFile/N25475 ) );
  AOI22_X1 U82721 ( .A1(n104818), .A2(n94519), .B1(n105469), .B2(n74286), .ZN(
        n95848) );
  OAI21_X1 U82722 ( .B1(n106330), .B2(n105471), .A(n95849), .ZN(
        \DLX_Datapath/RegisterFile/N25474 ) );
  AOI22_X1 U82723 ( .A1(n104818), .A2(n80192), .B1(n105468), .B2(n73722), .ZN(
        n95849) );
  OAI21_X1 U82724 ( .B1(n81315), .B2(n105470), .A(n95850), .ZN(
        \DLX_Datapath/RegisterFile/N25473 ) );
  AOI22_X1 U82725 ( .A1(n104816), .A2(n81474), .B1(n105468), .B2(n73426), .ZN(
        n95850) );
  OAI21_X1 U82726 ( .B1(n106128), .B2(n105470), .A(n95851), .ZN(
        \DLX_Datapath/RegisterFile/N25472 ) );
  AOI22_X1 U82727 ( .A1(n104818), .A2(n94523), .B1(n105468), .B2(n73863), .ZN(
        n95851) );
  OAI21_X1 U82728 ( .B1(n81318), .B2(n105470), .A(n95852), .ZN(
        \DLX_Datapath/RegisterFile/N25471 ) );
  AOI22_X1 U82729 ( .A1(n104816), .A2(n106060), .B1(n105468), .B2(n73575), 
        .ZN(n95852) );
  OAI21_X1 U82730 ( .B1(n106164), .B2(n105470), .A(n95853), .ZN(
        \DLX_Datapath/RegisterFile/N25470 ) );
  AOI22_X1 U82731 ( .A1(n104816), .A2(n81347), .B1(n105468), .B2(n73137), .ZN(
        n95853) );
  OAI21_X1 U82732 ( .B1(n81403), .B2(n105470), .A(n95854), .ZN(
        \DLX_Datapath/RegisterFile/N25469 ) );
  AOI22_X1 U82733 ( .A1(n104816), .A2(n94527), .B1(n105468), .B2(n73279), .ZN(
        n95854) );
  OAI21_X1 U82734 ( .B1(n106220), .B2(n105470), .A(n95855), .ZN(
        \DLX_Datapath/RegisterFile/N25468 ) );
  AOI22_X1 U82735 ( .A1(n104816), .A2(n81297), .B1(n105468), .B2(n72995), .ZN(
        n95855) );
  OAI21_X1 U82736 ( .B1(n106108), .B2(n105470), .A(n95856), .ZN(
        \DLX_Datapath/RegisterFile/N25467 ) );
  AOI22_X1 U82737 ( .A1(n104817), .A2(n94530), .B1(n105468), .B2(n72845), .ZN(
        n95856) );
  OAI21_X1 U82738 ( .B1(n106230), .B2(n105470), .A(n95857), .ZN(
        \DLX_Datapath/RegisterFile/N25466 ) );
  AOI22_X1 U82739 ( .A1(n104817), .A2(n81286), .B1(n105468), .B2(n70741), .ZN(
        n95857) );
  OAI21_X1 U82740 ( .B1(n106170), .B2(n105470), .A(n95858), .ZN(
        \DLX_Datapath/RegisterFile/N25465 ) );
  AOI22_X1 U82741 ( .A1(n104817), .A2(n106167), .B1(n105468), .B2(n70900), 
        .ZN(n95858) );
  AOI22_X1 U82743 ( .A1(n104818), .A2(n81283), .B1(n105468), .B2(n71045), .ZN(
        n95859) );
  OAI21_X1 U82744 ( .B1(n81451), .B2(n105470), .A(n95860), .ZN(
        \DLX_Datapath/RegisterFile/N25463 ) );
  AOI22_X1 U82745 ( .A1(n104818), .A2(n81453), .B1(n105468), .B2(n70006), .ZN(
        n95860) );
  OAI21_X1 U82746 ( .B1(n81310), .B2(n105470), .A(n95861), .ZN(
        \DLX_Datapath/RegisterFile/N25462 ) );
  AOI22_X1 U82747 ( .A1(n104816), .A2(n105626), .B1(n105469), .B2(n72535), 
        .ZN(n95861) );
  OAI21_X1 U82748 ( .B1(n106245), .B2(n105471), .A(n95862), .ZN(
        \DLX_Datapath/RegisterFile/N25461 ) );
  AOI22_X1 U82749 ( .A1(n104817), .A2(n106240), .B1(n105469), .B2(n71194), 
        .ZN(n95862) );
  OAI21_X1 U82750 ( .B1(n81349), .B2(n105471), .A(n95863), .ZN(
        \DLX_Datapath/RegisterFile/N25460 ) );
  AOI22_X1 U82751 ( .A1(n104818), .A2(n81351), .B1(n105469), .B2(n72677), .ZN(
        n95863) );
  OAI21_X1 U82752 ( .B1(n106113), .B2(n105471), .A(n95864), .ZN(
        \DLX_Datapath/RegisterFile/N25459 ) );
  AOI22_X1 U82753 ( .A1(n104817), .A2(n106019), .B1(n105468), .B2(n72387), 
        .ZN(n95864) );
  OAI21_X1 U82754 ( .B1(n106008), .B2(n105471), .A(n95865), .ZN(
        \DLX_Datapath/RegisterFile/N25458 ) );
  AOI22_X1 U82755 ( .A1(n104816), .A2(n94541), .B1(n95841), .B2(n71787), .ZN(
        n95865) );
  OAI21_X1 U82756 ( .B1(n106261), .B2(n105471), .A(n95866), .ZN(
        \DLX_Datapath/RegisterFile/N25457 ) );
  AOI22_X1 U82757 ( .A1(n104817), .A2(n81269), .B1(n95841), .B2(n72236), .ZN(
        n95866) );
  OAI21_X1 U82758 ( .B1(n106043), .B2(n105471), .A(n95867), .ZN(
        \DLX_Datapath/RegisterFile/N25456 ) );
  AOI22_X1 U82759 ( .A1(n104817), .A2(n105623), .B1(n95841), .B2(n72085), .ZN(
        n95867) );
  OAI21_X1 U82760 ( .B1(n106048), .B2(n105471), .A(n95868), .ZN(
        \DLX_Datapath/RegisterFile/N25455 ) );
  AOI22_X1 U82761 ( .A1(n104817), .A2(n105622), .B1(n95841), .B2(n71941), .ZN(
        n95868) );
  OAI21_X1 U82762 ( .B1(n81415), .B2(n105471), .A(n95869), .ZN(
        \DLX_Datapath/RegisterFile/N25454 ) );
  AOI22_X1 U82763 ( .A1(n104818), .A2(n105621), .B1(n105469), .B2(n71343), 
        .ZN(n95869) );
  OAI21_X1 U82764 ( .B1(n81498), .B2(n105470), .A(n95870), .ZN(
        \DLX_Datapath/RegisterFile/N25453 ) );
  AOI22_X1 U82765 ( .A1(n104818), .A2(n105911), .B1(n105469), .B2(n71638), 
        .ZN(n95870) );
  OAI21_X1 U82766 ( .B1(n105215), .B2(n105471), .A(n95871), .ZN(
        \DLX_Datapath/RegisterFile/N25452 ) );
  AOI22_X1 U82767 ( .A1(n104817), .A2(n80188), .B1(n95841), .B2(n71494), .ZN(
        n95871) );
  OAI21_X1 U82768 ( .B1(n106267), .B2(n105471), .A(n95872), .ZN(
        \DLX_Datapath/RegisterFile/N25451 ) );
  AOI22_X1 U82769 ( .A1(n104816), .A2(n81265), .B1(n95841), .B2(n69603), .ZN(
        n95872) );
  AOI21_X1 U82770 ( .B1(n95450), .B2(n94771), .A(n104701), .ZN(n95841) );
  NAND2_X1 U82771 ( .A1(n95517), .A2(n105205), .ZN(n95450) );
  NOR2_X1 U82772 ( .A1(n95874), .A2(n95517), .ZN(n95840) );
  OR2_X1 U82773 ( .A1(n95873), .A2(n94848), .ZN(n95874) );
  NOR2_X1 U82774 ( .A1(n95838), .A2(n105091), .ZN(n95873) );
  NAND2_X1 U82775 ( .A1(n105133), .A2(n94772), .ZN(n95838) );
  OAI21_X1 U82776 ( .B1(n106147), .B2(n105467), .A(n95876), .ZN(
        \DLX_Datapath/RegisterFile/N25450 ) );
  AOI22_X1 U82777 ( .A1(n105466), .A2(n70304), .B1(n105463), .B2(n94559), .ZN(
        n95876) );
  OAI21_X1 U82778 ( .B1(n105970), .B2(n105467), .A(n95879), .ZN(
        \DLX_Datapath/RegisterFile/N25449 ) );
  AOI22_X1 U82779 ( .A1(n105465), .A2(n70446), .B1(n105462), .B2(n94562), .ZN(
        n95879) );
  OAI21_X1 U82780 ( .B1(n106135), .B2(n105467), .A(n95880), .ZN(
        \DLX_Datapath/RegisterFile/N25448 ) );
  AOI22_X1 U82781 ( .A1(n105466), .A2(n107223), .B1(n105463), .B2(n94564), 
        .ZN(n95880) );
  OAI21_X1 U82782 ( .B1(n106211), .B2(n105467), .A(n95881), .ZN(
        \DLX_Datapath/RegisterFile/N25447 ) );
  AOI22_X1 U82783 ( .A1(n105465), .A2(n107761), .B1(n105462), .B2(n94566), 
        .ZN(n95881) );
  OAI21_X1 U82784 ( .B1(n106203), .B2(n105467), .A(n95882), .ZN(
        \DLX_Datapath/RegisterFile/N25446 ) );
  AOI22_X1 U82785 ( .A1(n105466), .A2(n110664), .B1(n105463), .B2(n94568), 
        .ZN(n95882) );
  OAI21_X1 U82786 ( .B1(n106100), .B2(n105467), .A(n95883), .ZN(
        \DLX_Datapath/RegisterFile/N25445 ) );
  AOI22_X1 U82787 ( .A1(n105465), .A2(n108063), .B1(n105462), .B2(n94570), 
        .ZN(n95883) );
  OAI21_X1 U82788 ( .B1(n106256), .B2(n105467), .A(n95884), .ZN(
        \DLX_Datapath/RegisterFile/N25444 ) );
  AOI22_X1 U82789 ( .A1(n105466), .A2(n110761), .B1(n105463), .B2(n94572), 
        .ZN(n95884) );
  OAI21_X1 U82790 ( .B1(n105990), .B2(n105467), .A(n95885), .ZN(
        \DLX_Datapath/RegisterFile/N25443 ) );
  AOI22_X1 U82791 ( .A1(n105465), .A2(n110862), .B1(n105462), .B2(n94574), 
        .ZN(n95885) );
  OAI21_X1 U82792 ( .B1(n106332), .B2(n105467), .A(n95886), .ZN(
        \DLX_Datapath/RegisterFile/N25442 ) );
  AOI22_X1 U82793 ( .A1(n105465), .A2(n110457), .B1(n105462), .B2(n94576), 
        .ZN(n95886) );
  OAI21_X1 U82794 ( .B1(n106192), .B2(n105467), .A(n95887), .ZN(
        \DLX_Datapath/RegisterFile/N25441 ) );
  AOI22_X1 U82795 ( .A1(n105464), .A2(n110239), .B1(n105461), .B2(n94578), 
        .ZN(n95887) );
  OAI21_X1 U82796 ( .B1(n106128), .B2(n105467), .A(n95888), .ZN(
        \DLX_Datapath/RegisterFile/N25440 ) );
  AOI22_X1 U82797 ( .A1(n105464), .A2(n110556), .B1(n105461), .B2(n94580), 
        .ZN(n95888) );
  OAI21_X1 U82798 ( .B1(n106188), .B2(n105467), .A(n95889), .ZN(
        \DLX_Datapath/RegisterFile/N25439 ) );
  AOI22_X1 U82799 ( .A1(n105464), .A2(n110347), .B1(n105461), .B2(n94582), 
        .ZN(n95889) );
  OAI21_X1 U82800 ( .B1(n106162), .B2(n105467), .A(n95890), .ZN(
        \DLX_Datapath/RegisterFile/N25438 ) );
  AOI22_X1 U82801 ( .A1(n105464), .A2(n110022), .B1(n105461), .B2(n94584), 
        .ZN(n95890) );
  OAI21_X1 U82802 ( .B1(n81403), .B2(n105467), .A(n95891), .ZN(
        \DLX_Datapath/RegisterFile/N25437 ) );
  AOI22_X1 U82803 ( .A1(n105464), .A2(n110129), .B1(n105461), .B2(n94586), 
        .ZN(n95891) );
  OAI21_X1 U82804 ( .B1(n81294), .B2(n105467), .A(n95892), .ZN(
        \DLX_Datapath/RegisterFile/N25436 ) );
  AOI22_X1 U82805 ( .A1(n105464), .A2(n109913), .B1(n105461), .B2(n94588), 
        .ZN(n95892) );
  OAI21_X1 U82806 ( .B1(n106108), .B2(n105467), .A(n95893), .ZN(
        \DLX_Datapath/RegisterFile/N25435 ) );
  AOI22_X1 U82807 ( .A1(n105464), .A2(n109795), .B1(n105461), .B2(n94590), 
        .ZN(n95893) );
  OAI21_X1 U82808 ( .B1(n81284), .B2(n105467), .A(n95894), .ZN(
        \DLX_Datapath/RegisterFile/N25434 ) );
  AOI22_X1 U82809 ( .A1(n105464), .A2(n108169), .B1(n105461), .B2(n94592), 
        .ZN(n95894) );
  OAI21_X1 U82810 ( .B1(n106172), .B2(n105467), .A(n95895), .ZN(
        \DLX_Datapath/RegisterFile/N25433 ) );
  AOI22_X1 U82811 ( .A1(n105464), .A2(n108292), .B1(n105461), .B2(n94594), 
        .ZN(n95895) );
  OAI21_X1 U82812 ( .B1(n106236), .B2(n105467), .A(n95896), .ZN(
        \DLX_Datapath/RegisterFile/N25432 ) );
  AOI22_X1 U82813 ( .A1(n105464), .A2(n108403), .B1(n105461), .B2(n94596), 
        .ZN(n95896) );
  OAI21_X1 U82814 ( .B1(n81451), .B2(n105467), .A(n95897), .ZN(
        \DLX_Datapath/RegisterFile/N25431 ) );
  AOI22_X1 U82815 ( .A1(n105464), .A2(n107641), .B1(n105461), .B2(n94598), 
        .ZN(n95897) );
  OAI21_X1 U82816 ( .B1(n106199), .B2(n105467), .A(n95898), .ZN(
        \DLX_Datapath/RegisterFile/N25430 ) );
  AOI22_X1 U82817 ( .A1(n105465), .A2(n109559), .B1(n105462), .B2(n94600), 
        .ZN(n95898) );
  OAI21_X1 U82818 ( .B1(n106245), .B2(n95875), .A(n95899), .ZN(
        \DLX_Datapath/RegisterFile/N25429 ) );
  AOI22_X1 U82819 ( .A1(n105466), .A2(n108520), .B1(n105463), .B2(n94602), 
        .ZN(n95899) );
  OAI21_X1 U82820 ( .B1(n81349), .B2(n95875), .A(n95900), .ZN(
        \DLX_Datapath/RegisterFile/N25428 ) );
  AOI22_X1 U82821 ( .A1(n105465), .A2(n109664), .B1(n105462), .B2(n94604), 
        .ZN(n95900) );
  OAI21_X1 U82822 ( .B1(n106113), .B2(n95875), .A(n95901), .ZN(
        \DLX_Datapath/RegisterFile/N25427 ) );
  AOI22_X1 U82823 ( .A1(n105466), .A2(n109448), .B1(n105463), .B2(n94606), 
        .ZN(n95901) );
  OAI21_X1 U82824 ( .B1(n106011), .B2(n95875), .A(n95902), .ZN(
        \DLX_Datapath/RegisterFile/N25426 ) );
  AOI22_X1 U82825 ( .A1(n105465), .A2(n108985), .B1(n105462), .B2(n94608), 
        .ZN(n95902) );
  OAI21_X1 U82826 ( .B1(n106262), .B2(n95875), .A(n95903), .ZN(
        \DLX_Datapath/RegisterFile/N25425 ) );
  AOI22_X1 U82827 ( .A1(n105466), .A2(n109333), .B1(n105463), .B2(n94610), 
        .ZN(n95903) );
  OAI21_X1 U82828 ( .B1(n106043), .B2(n95875), .A(n95904), .ZN(
        \DLX_Datapath/RegisterFile/N25424 ) );
  AOI22_X1 U82829 ( .A1(n105465), .A2(n109215), .B1(n105462), .B2(n94612), 
        .ZN(n95904) );
  OAI21_X1 U82830 ( .B1(n106048), .B2(n95875), .A(n95905), .ZN(
        \DLX_Datapath/RegisterFile/N25423 ) );
  AOI22_X1 U82831 ( .A1(n105466), .A2(n109107), .B1(n105463), .B2(n94614), 
        .ZN(n95905) );
  OAI21_X1 U82832 ( .B1(n81415), .B2(n95875), .A(n95906), .ZN(
        \DLX_Datapath/RegisterFile/N25422 ) );
  AOI22_X1 U82833 ( .A1(n105465), .A2(n108642), .B1(n105462), .B2(n94616), 
        .ZN(n95906) );
  OAI21_X1 U82834 ( .B1(n106053), .B2(n95875), .A(n95907), .ZN(
        \DLX_Datapath/RegisterFile/N25421 ) );
  AOI22_X1 U82835 ( .A1(n105466), .A2(n108869), .B1(n105463), .B2(n94618), 
        .ZN(n95907) );
  OAI21_X1 U82836 ( .B1(n105215), .B2(n95875), .A(n95908), .ZN(
        \DLX_Datapath/RegisterFile/N25420 ) );
  AOI22_X1 U82837 ( .A1(n105466), .A2(n108757), .B1(n105463), .B2(n94620), 
        .ZN(n95908) );
  OAI21_X1 U82838 ( .B1(n106267), .B2(n105467), .A(n95909), .ZN(
        \DLX_Datapath/RegisterFile/N25419 ) );
  AOI22_X1 U82839 ( .A1(n105465), .A2(n107297), .B1(n105462), .B2(n94622), 
        .ZN(n95909) );
  NOR2_X1 U82843 ( .A1(n95875), .A2(n105091), .ZN(n95911) );
  NAND2_X1 U82844 ( .A1(n105134), .A2(n94810), .ZN(n95875) );
  OAI21_X1 U82845 ( .B1(n106148), .B2(n105460), .A(n95914), .ZN(
        \DLX_Datapath/RegisterFile/N25418 ) );
  AOI22_X1 U82846 ( .A1(n105459), .A2(n107864), .B1(n105457), .B2(n81521), 
        .ZN(n95914) );
  OAI21_X1 U82847 ( .B1(n105968), .B2(n105460), .A(n95917), .ZN(
        \DLX_Datapath/RegisterFile/N25417 ) );
  AOI22_X1 U82848 ( .A1(n95915), .A2(n107961), .B1(n105456), .B2(n81653), .ZN(
        n95917) );
  OAI21_X1 U82849 ( .B1(n106135), .B2(n105460), .A(n95918), .ZN(
        \DLX_Datapath/RegisterFile/N25416 ) );
  AOI22_X1 U82850 ( .A1(n105459), .A2(n107224), .B1(n105457), .B2(n81380), 
        .ZN(n95918) );
  OAI21_X1 U82851 ( .B1(n106208), .B2(n105460), .A(n95919), .ZN(
        \DLX_Datapath/RegisterFile/N25415 ) );
  AOI22_X1 U82852 ( .A1(n105459), .A2(n107762), .B1(n105456), .B2(n81377), 
        .ZN(n95919) );
  OAI21_X1 U82853 ( .B1(n106203), .B2(n105460), .A(n95920), .ZN(
        \DLX_Datapath/RegisterFile/N25414 ) );
  AOI22_X1 U82854 ( .A1(n105459), .A2(n110665), .B1(n105457), .B2(n81428), 
        .ZN(n95920) );
  OAI21_X1 U82855 ( .B1(n106099), .B2(n105460), .A(n95921), .ZN(
        \DLX_Datapath/RegisterFile/N25413 ) );
  AOI22_X1 U82856 ( .A1(n105458), .A2(n108064), .B1(n105456), .B2(n81410), 
        .ZN(n95921) );
  OAI21_X1 U82857 ( .B1(n106254), .B2(n105460), .A(n95922), .ZN(
        \DLX_Datapath/RegisterFile/N25412 ) );
  AOI22_X1 U82858 ( .A1(n95915), .A2(n110762), .B1(n105456), .B2(n81700), .ZN(
        n95922) );
  OAI21_X1 U82859 ( .B1(n105991), .B2(n105460), .A(n95923), .ZN(
        \DLX_Datapath/RegisterFile/N25411 ) );
  AOI22_X1 U82860 ( .A1(n105459), .A2(n110863), .B1(n105457), .B2(n81632), 
        .ZN(n95923) );
  OAI21_X1 U82861 ( .B1(n106331), .B2(n105460), .A(n95924), .ZN(
        \DLX_Datapath/RegisterFile/N25410 ) );
  AOI22_X1 U82862 ( .A1(n95915), .A2(n110458), .B1(n105456), .B2(n81414), .ZN(
        n95924) );
  OAI21_X1 U82863 ( .B1(n106193), .B2(n105460), .A(n95925), .ZN(
        \DLX_Datapath/RegisterFile/N25409 ) );
  AOI22_X1 U82864 ( .A1(n105458), .A2(n110240), .B1(n105455), .B2(n81317), 
        .ZN(n95925) );
  OAI21_X1 U82865 ( .B1(n106128), .B2(n105460), .A(n95926), .ZN(
        \DLX_Datapath/RegisterFile/N25408 ) );
  AOI22_X1 U82866 ( .A1(n105458), .A2(n110557), .B1(n105455), .B2(n81386), 
        .ZN(n95926) );
  OAI21_X1 U82867 ( .B1(n106185), .B2(n105460), .A(n95927), .ZN(
        \DLX_Datapath/RegisterFile/N25407 ) );
  AOI22_X1 U82868 ( .A1(n105458), .A2(n110348), .B1(n105455), .B2(n81320), 
        .ZN(n95927) );
  OAI21_X1 U82869 ( .B1(n106163), .B2(n105460), .A(n95928), .ZN(
        \DLX_Datapath/RegisterFile/N25406 ) );
  AOI22_X1 U82870 ( .A1(n105458), .A2(n110023), .B1(n105455), .B2(n81604), 
        .ZN(n95928) );
  OAI21_X1 U82871 ( .B1(n81403), .B2(n105460), .A(n95929), .ZN(
        \DLX_Datapath/RegisterFile/N25405 ) );
  AOI22_X1 U82872 ( .A1(n105458), .A2(n110130), .B1(n105455), .B2(n81405), 
        .ZN(n95929) );
  OAI21_X1 U82873 ( .B1(n106221), .B2(n105460), .A(n95930), .ZN(
        \DLX_Datapath/RegisterFile/N25404 ) );
  AOI22_X1 U82874 ( .A1(n105458), .A2(n109914), .B1(n105455), .B2(n81402), 
        .ZN(n95930) );
  OAI21_X1 U82875 ( .B1(n106108), .B2(n105460), .A(n95931), .ZN(
        \DLX_Datapath/RegisterFile/N25403 ) );
  AOI22_X1 U82876 ( .A1(n105458), .A2(n109796), .B1(n105455), .B2(n81400), 
        .ZN(n95931) );
  OAI21_X1 U82877 ( .B1(n106232), .B2(n105460), .A(n95932), .ZN(
        \DLX_Datapath/RegisterFile/N25402 ) );
  AOI22_X1 U82878 ( .A1(n105458), .A2(n108170), .B1(n105455), .B2(n81332), 
        .ZN(n95932) );
  OAI21_X1 U82879 ( .B1(n106173), .B2(n105460), .A(n95933), .ZN(
        \DLX_Datapath/RegisterFile/N25401 ) );
  AOI22_X1 U82880 ( .A1(n105458), .A2(n108293), .B1(n105455), .B2(n81373), 
        .ZN(n95933) );
  OAI21_X1 U82881 ( .B1(n106236), .B2(n105460), .A(n95934), .ZN(
        \DLX_Datapath/RegisterFile/N25400 ) );
  AOI22_X1 U82882 ( .A1(n105458), .A2(n108404), .B1(n105455), .B2(n81322), 
        .ZN(n95934) );
  OAI21_X1 U82883 ( .B1(n106072), .B2(n105460), .A(n95935), .ZN(
        \DLX_Datapath/RegisterFile/N25399 ) );
  AOI22_X1 U82884 ( .A1(n105458), .A2(n107642), .B1(n105455), .B2(n81506), 
        .ZN(n95935) );
  OAI21_X1 U82885 ( .B1(n106200), .B2(n105460), .A(n95936), .ZN(
        \DLX_Datapath/RegisterFile/N25398 ) );
  AOI22_X1 U82886 ( .A1(n105458), .A2(n109560), .B1(n105456), .B2(n81313), 
        .ZN(n95936) );
  OAI21_X1 U82887 ( .B1(n81278), .B2(n105460), .A(n95937), .ZN(
        \DLX_Datapath/RegisterFile/N25397 ) );
  AOI22_X1 U82888 ( .A1(n105459), .A2(n108521), .B1(n105457), .B2(n81330), 
        .ZN(n95937) );
  OAI21_X1 U82889 ( .B1(n81349), .B2(n105460), .A(n95938), .ZN(
        \DLX_Datapath/RegisterFile/N25396 ) );
  AOI22_X1 U82890 ( .A1(n95915), .A2(n109665), .B1(n105456), .B2(n81425), .ZN(
        n95938) );
  OAI21_X1 U82891 ( .B1(n106113), .B2(n105460), .A(n95939), .ZN(
        \DLX_Datapath/RegisterFile/N25395 ) );
  AOI22_X1 U82892 ( .A1(n105459), .A2(n109449), .B1(n105457), .B2(n81396), 
        .ZN(n95939) );
  OAI21_X1 U82893 ( .B1(n81588), .B2(n105460), .A(n95940), .ZN(
        \DLX_Datapath/RegisterFile/N25394 ) );
  AOI22_X1 U82894 ( .A1(n105458), .A2(n108986), .B1(n105456), .B2(n81590), 
        .ZN(n95940) );
  OAI21_X1 U82895 ( .B1(n81267), .B2(n105460), .A(n95941), .ZN(
        \DLX_Datapath/RegisterFile/N25393 ) );
  AOI22_X1 U82896 ( .A1(n105459), .A2(n109334), .B1(n105457), .B2(n81423), 
        .ZN(n95941) );
  OAI21_X1 U82897 ( .B1(n106043), .B2(n105460), .A(n95942), .ZN(
        \DLX_Datapath/RegisterFile/N25392 ) );
  AOI22_X1 U82898 ( .A1(n95915), .A2(n109216), .B1(n105456), .B2(n81511), .ZN(
        n95942) );
  OAI21_X1 U82899 ( .B1(n106048), .B2(n105460), .A(n95943), .ZN(
        \DLX_Datapath/RegisterFile/N25391 ) );
  AOI22_X1 U82900 ( .A1(n105459), .A2(n109108), .B1(n105457), .B2(n81503), 
        .ZN(n95943) );
  OAI21_X1 U82901 ( .B1(n81415), .B2(n105460), .A(n95944), .ZN(
        \DLX_Datapath/RegisterFile/N25390 ) );
  AOI22_X1 U82902 ( .A1(n95915), .A2(n108643), .B1(n105456), .B2(n81417), .ZN(
        n95944) );
  OAI21_X1 U82903 ( .B1(n106055), .B2(n105460), .A(n95945), .ZN(
        \DLX_Datapath/RegisterFile/N25389 ) );
  AOI22_X1 U82904 ( .A1(n105459), .A2(n108870), .B1(n105457), .B2(n81500), 
        .ZN(n95945) );
  OAI21_X1 U82905 ( .B1(n105217), .B2(n105460), .A(n95946), .ZN(
        \DLX_Datapath/RegisterFile/N25388 ) );
  AOI22_X1 U82906 ( .A1(n105459), .A2(n108758), .B1(n105457), .B2(n81335), 
        .ZN(n95946) );
  OAI21_X1 U82907 ( .B1(n81262), .B2(n105460), .A(n95947), .ZN(
        \DLX_Datapath/RegisterFile/N25387 ) );
  AOI22_X1 U82908 ( .A1(n95915), .A2(n107298), .B1(n105456), .B2(n81327), .ZN(
        n95947) );
  OR2_X1 U82910 ( .A1(n95949), .A2(n94848), .ZN(n95948) );
  NOR2_X1 U82911 ( .A1(n95949), .A2(n95912), .ZN(n95915) );
  AOI21_X1 U82912 ( .B1(n105204), .B2(n95950), .A(n94663), .ZN(n95912) );
  OR2_X1 U82913 ( .A1(n94848), .A2(n95517), .ZN(n95950) );
  NAND2_X1 U82914 ( .A1(n95951), .A2(n94850), .ZN(n95517) );
  NOR2_X1 U82915 ( .A1(n94852), .A2(n106763), .ZN(n95951) );
  NOR2_X1 U82916 ( .A1(n95913), .A2(n105089), .ZN(n95949) );
  NAND2_X1 U82917 ( .A1(n105133), .A2(n94853), .ZN(n95913) );
  OAI21_X1 U82918 ( .B1(n106146), .B2(n105454), .A(n95953), .ZN(
        \DLX_Datapath/RegisterFile/N25386 ) );
  AOI22_X1 U82919 ( .A1(n105453), .A2(n94667), .B1(n95955), .B2(n107865), .ZN(
        n95953) );
  OAI21_X1 U82920 ( .B1(n105969), .B2(n105454), .A(n95956), .ZN(
        \DLX_Datapath/RegisterFile/N25385 ) );
  AOI22_X1 U82921 ( .A1(n105452), .A2(n94670), .B1(n104965), .B2(n107962), 
        .ZN(n95956) );
  OAI21_X1 U82922 ( .B1(n106135), .B2(n105454), .A(n95957), .ZN(
        \DLX_Datapath/RegisterFile/N25384 ) );
  AOI22_X1 U82923 ( .A1(n105453), .A2(n94672), .B1(n95955), .B2(n107225), .ZN(
        n95957) );
  OAI21_X1 U82924 ( .B1(n106209), .B2(n105454), .A(n95958), .ZN(
        \DLX_Datapath/RegisterFile/N25383 ) );
  AOI22_X1 U82925 ( .A1(n105452), .A2(n94674), .B1(n104966), .B2(n107763), 
        .ZN(n95958) );
  OAI21_X1 U82926 ( .B1(n106203), .B2(n105454), .A(n95959), .ZN(
        \DLX_Datapath/RegisterFile/N25382 ) );
  AOI22_X1 U82927 ( .A1(n105453), .A2(n94676), .B1(n95955), .B2(n110666), .ZN(
        n95959) );
  OAI21_X1 U82928 ( .B1(n106098), .B2(n105454), .A(n95960), .ZN(
        \DLX_Datapath/RegisterFile/N25381 ) );
  AOI22_X1 U82929 ( .A1(n105452), .A2(n94678), .B1(n104965), .B2(n108065), 
        .ZN(n95960) );
  OAI21_X1 U82930 ( .B1(n106255), .B2(n105454), .A(n95961), .ZN(
        \DLX_Datapath/RegisterFile/N25380 ) );
  AOI22_X1 U82931 ( .A1(n105453), .A2(n94680), .B1(n104965), .B2(n110763), 
        .ZN(n95961) );
  OAI21_X1 U82932 ( .B1(n105992), .B2(n105454), .A(n95962), .ZN(
        \DLX_Datapath/RegisterFile/N25379 ) );
  AOI22_X1 U82933 ( .A1(n105452), .A2(n94682), .B1(n104966), .B2(n110864), 
        .ZN(n95962) );
  OAI21_X1 U82934 ( .B1(n80190), .B2(n105454), .A(n95963), .ZN(
        \DLX_Datapath/RegisterFile/N25378 ) );
  AOI22_X1 U82935 ( .A1(n105452), .A2(n94684), .B1(n104965), .B2(n110459), 
        .ZN(n95963) );
  OAI21_X1 U82936 ( .B1(n106190), .B2(n105454), .A(n95964), .ZN(
        \DLX_Datapath/RegisterFile/N25377 ) );
  AOI22_X1 U82937 ( .A1(n105451), .A2(n94686), .B1(n95955), .B2(n110241), .ZN(
        n95964) );
  OAI21_X1 U82938 ( .B1(n106128), .B2(n105454), .A(n95965), .ZN(
        \DLX_Datapath/RegisterFile/N25376 ) );
  AOI22_X1 U82939 ( .A1(n105451), .A2(n94688), .B1(n104965), .B2(n110558), 
        .ZN(n95965) );
  OAI21_X1 U82940 ( .B1(n106185), .B2(n105454), .A(n95966), .ZN(
        \DLX_Datapath/RegisterFile/N25375 ) );
  AOI22_X1 U82941 ( .A1(n105451), .A2(n94690), .B1(n104966), .B2(n110349), 
        .ZN(n95966) );
  OAI21_X1 U82942 ( .B1(n81345), .B2(n105454), .A(n95967), .ZN(
        \DLX_Datapath/RegisterFile/N25374 ) );
  AOI22_X1 U82943 ( .A1(n105451), .A2(n94692), .B1(n104966), .B2(n110024), 
        .ZN(n95967) );
  OAI21_X1 U82944 ( .B1(n81403), .B2(n105454), .A(n95968), .ZN(
        \DLX_Datapath/RegisterFile/N25373 ) );
  AOI22_X1 U82945 ( .A1(n105451), .A2(n94694), .B1(n104965), .B2(n110131), 
        .ZN(n95968) );
  OAI21_X1 U82946 ( .B1(n81294), .B2(n105454), .A(n95969), .ZN(
        \DLX_Datapath/RegisterFile/N25372 ) );
  AOI22_X1 U82947 ( .A1(n105451), .A2(n94696), .B1(n104966), .B2(n109915), 
        .ZN(n95969) );
  OAI21_X1 U82948 ( .B1(n106108), .B2(n105454), .A(n95970), .ZN(
        \DLX_Datapath/RegisterFile/N25371 ) );
  AOI22_X1 U82949 ( .A1(n105451), .A2(n94698), .B1(n104965), .B2(n109797), 
        .ZN(n95970) );
  OAI21_X1 U82950 ( .B1(n81284), .B2(n105454), .A(n95971), .ZN(
        \DLX_Datapath/RegisterFile/N25370 ) );
  AOI22_X1 U82951 ( .A1(n105451), .A2(n94700), .B1(n104966), .B2(n108171), 
        .ZN(n95971) );
  OAI21_X1 U82952 ( .B1(n106173), .B2(n105454), .A(n95972), .ZN(
        \DLX_Datapath/RegisterFile/N25369 ) );
  AOI22_X1 U82953 ( .A1(n105451), .A2(n94702), .B1(n104965), .B2(n108294), 
        .ZN(n95972) );
  OAI21_X1 U82954 ( .B1(n106236), .B2(n105454), .A(n95973), .ZN(
        \DLX_Datapath/RegisterFile/N25368 ) );
  AOI22_X1 U82955 ( .A1(n105451), .A2(n94704), .B1(n104965), .B2(n108405), 
        .ZN(n95973) );
  OAI21_X1 U82956 ( .B1(n106072), .B2(n105454), .A(n95974), .ZN(
        \DLX_Datapath/RegisterFile/N25367 ) );
  AOI22_X1 U82957 ( .A1(n105451), .A2(n94706), .B1(n104965), .B2(n107643), 
        .ZN(n95974) );
  OAI21_X1 U82958 ( .B1(n106197), .B2(n105454), .A(n95975), .ZN(
        \DLX_Datapath/RegisterFile/N25366 ) );
  AOI22_X1 U82959 ( .A1(n105452), .A2(n94708), .B1(n104966), .B2(n109561), 
        .ZN(n95975) );
  OAI21_X1 U82960 ( .B1(n81278), .B2(n105454), .A(n95976), .ZN(
        \DLX_Datapath/RegisterFile/N25365 ) );
  AOI22_X1 U82961 ( .A1(n105453), .A2(n94710), .B1(n104966), .B2(n108522), 
        .ZN(n95976) );
  OAI21_X1 U82962 ( .B1(n81349), .B2(n105454), .A(n95977), .ZN(
        \DLX_Datapath/RegisterFile/N25364 ) );
  AOI22_X1 U82963 ( .A1(n105452), .A2(n94712), .B1(n104966), .B2(n109666), 
        .ZN(n95977) );
  OAI21_X1 U82964 ( .B1(n106113), .B2(n105454), .A(n95978), .ZN(
        \DLX_Datapath/RegisterFile/N25363 ) );
  AOI22_X1 U82965 ( .A1(n105453), .A2(n94714), .B1(n95955), .B2(n109450), .ZN(
        n95978) );
  OAI21_X1 U82966 ( .B1(n106007), .B2(n105454), .A(n95979), .ZN(
        \DLX_Datapath/RegisterFile/N25362 ) );
  AOI22_X1 U82967 ( .A1(n105452), .A2(n81259), .B1(n95955), .B2(n108987), .ZN(
        n95979) );
  OAI21_X1 U82968 ( .B1(n81267), .B2(n105454), .A(n95980), .ZN(
        \DLX_Datapath/RegisterFile/N25361 ) );
  AOI22_X1 U82969 ( .A1(n105453), .A2(n94717), .B1(n104965), .B2(n109335), 
        .ZN(n95980) );
  OAI21_X1 U82970 ( .B1(n106043), .B2(n105454), .A(n95981), .ZN(
        \DLX_Datapath/RegisterFile/N25360 ) );
  AOI22_X1 U82971 ( .A1(n105452), .A2(n94719), .B1(n104966), .B2(n109217), 
        .ZN(n95981) );
  OAI21_X1 U82972 ( .B1(n106048), .B2(n105454), .A(n95982), .ZN(
        \DLX_Datapath/RegisterFile/N25359 ) );
  AOI22_X1 U82973 ( .A1(n105453), .A2(n94721), .B1(n104965), .B2(n109109), 
        .ZN(n95982) );
  OAI21_X1 U82974 ( .B1(n81415), .B2(n105454), .A(n95983), .ZN(
        \DLX_Datapath/RegisterFile/N25358 ) );
  AOI22_X1 U82975 ( .A1(n105452), .A2(n94723), .B1(n95955), .B2(n108644), .ZN(
        n95983) );
  OAI21_X1 U82976 ( .B1(n106055), .B2(n105454), .A(n95984), .ZN(
        \DLX_Datapath/RegisterFile/N25357 ) );
  AOI22_X1 U82977 ( .A1(n105453), .A2(n94725), .B1(n104965), .B2(n108871), 
        .ZN(n95984) );
  OAI21_X1 U82978 ( .B1(n105216), .B2(n105454), .A(n95985), .ZN(
        \DLX_Datapath/RegisterFile/N25356 ) );
  AOI22_X1 U82979 ( .A1(n105453), .A2(n94727), .B1(n95955), .B2(n108759), .ZN(
        n95985) );
  OAI21_X1 U82980 ( .B1(n81262), .B2(n105454), .A(n95986), .ZN(
        \DLX_Datapath/RegisterFile/N25355 ) );
  AOI22_X1 U82981 ( .A1(n105452), .A2(n94729), .B1(n104966), .B2(n107299), 
        .ZN(n95986) );
  AOI21_X1 U82982 ( .B1(n95987), .B2(n105602), .A(n95988), .ZN(n95955) );
  OAI21_X1 U82983 ( .B1(n95555), .B2(n94848), .A(n105199), .ZN(n95987) );
  OR2_X1 U82985 ( .A1(n95990), .A2(n94852), .ZN(n95555) );
  NAND2_X1 U82986 ( .A1(n59515), .A2(n94851), .ZN(n95990) );
  OR2_X1 U82987 ( .A1(n95988), .A2(n94848), .ZN(n95989) );
  NOR2_X1 U82988 ( .A1(n95952), .A2(n105089), .ZN(n95988) );
  NAND2_X1 U82989 ( .A1(n94892), .A2(n105133), .ZN(n95952) );
  NOR2_X1 U82990 ( .A1(n95991), .A2(n94894), .ZN(n95452) );
  OAI21_X1 U82991 ( .B1(n105970), .B2(n105921), .A(n95992), .ZN(
        \DLX_Datapath/RegisterFile/N25353 ) );
  AOI22_X1 U82992 ( .A1(n94511), .A2(n104843), .B1(n105920), .B2(n107963), 
        .ZN(n95992) );
  OAI21_X1 U82993 ( .B1(n81408), .B2(n105921), .A(n95993), .ZN(
        \DLX_Datapath/RegisterFile/N25349 ) );
  AOI22_X1 U82994 ( .A1(n94516), .A2(n104843), .B1(n105920), .B2(n108066), 
        .ZN(n95993) );
  OAI21_X1 U82995 ( .B1(n106257), .B2(n105921), .A(n95994), .ZN(
        \DLX_Datapath/RegisterFile/N25348 ) );
  AOI22_X1 U82996 ( .A1(n81759), .A2(n81272), .B1(n105919), .B2(n110764), .ZN(
        n95994) );
  OAI21_X1 U82997 ( .B1(n105991), .B2(n105921), .A(n95995), .ZN(
        \DLX_Datapath/RegisterFile/N25347 ) );
  AOI22_X1 U82998 ( .A1(n94519), .A2(n104843), .B1(n105920), .B2(n110865), 
        .ZN(n95995) );
  OAI21_X1 U82999 ( .B1(n106332), .B2(n105921), .A(n95996), .ZN(
        \DLX_Datapath/RegisterFile/N25346 ) );
  AOI22_X1 U83000 ( .A1(n104719), .A2(n80192), .B1(n105919), .B2(n110460), 
        .ZN(n95996) );
  OAI21_X1 U83001 ( .B1(n106128), .B2(n105921), .A(n95997), .ZN(
        \DLX_Datapath/RegisterFile/N25344 ) );
  AOI22_X1 U83002 ( .A1(n94523), .A2(n104843), .B1(n81760), .B2(n110559), .ZN(
        n95997) );
  OAI21_X1 U83003 ( .B1(n81403), .B2(n105921), .A(n95998), .ZN(
        \DLX_Datapath/RegisterFile/N25341 ) );
  AOI22_X1 U83004 ( .A1(n94527), .A2(n104843), .B1(n105920), .B2(n110132), 
        .ZN(n95998) );
  OAI21_X1 U83005 ( .B1(n106221), .B2(n105922), .A(n95999), .ZN(
        \DLX_Datapath/RegisterFile/N25340 ) );
  AOI22_X1 U83006 ( .A1(n104820), .A2(n81297), .B1(n105919), .B2(n109916), 
        .ZN(n95999) );
  OAI21_X1 U83007 ( .B1(n106108), .B2(n105922), .A(n96000), .ZN(
        \DLX_Datapath/RegisterFile/N25339 ) );
  AOI22_X1 U83008 ( .A1(n94530), .A2(n81759), .B1(n81760), .B2(n109798), .ZN(
        n96000) );
  OAI21_X1 U83009 ( .B1(n106172), .B2(n105922), .A(n96001), .ZN(
        \DLX_Datapath/RegisterFile/N25337 ) );
  AOI22_X1 U83010 ( .A1(n104719), .A2(n106167), .B1(n105920), .B2(n108295), 
        .ZN(n96001) );
  OAI21_X1 U83011 ( .B1(n106072), .B2(n105921), .A(n96002), .ZN(
        \DLX_Datapath/RegisterFile/N25335 ) );
  AOI22_X1 U83012 ( .A1(n81759), .A2(n81453), .B1(n81760), .B2(n107644), .ZN(
        n96002) );
  OAI21_X1 U83013 ( .B1(n81310), .B2(n105922), .A(n96003), .ZN(
        \DLX_Datapath/RegisterFile/N25334 ) );
  AOI22_X1 U83014 ( .A1(n105626), .A2(n104820), .B1(n105920), .B2(n109562), 
        .ZN(n96003) );
  OAI21_X1 U83015 ( .B1(n106009), .B2(n105922), .A(n96004), .ZN(
        \DLX_Datapath/RegisterFile/N25330 ) );
  AOI22_X1 U83016 ( .A1(n94541), .A2(n104718), .B1(n81760), .B2(n108988), .ZN(
        n96004) );
  OAI21_X1 U83017 ( .B1(n106043), .B2(n105921), .A(n96005), .ZN(
        \DLX_Datapath/RegisterFile/N25328 ) );
  AOI22_X1 U83018 ( .A1(n105623), .A2(n104820), .B1(n105920), .B2(n109218), 
        .ZN(n96005) );
  OAI21_X1 U83019 ( .B1(n106048), .B2(n105922), .A(n96006), .ZN(
        \DLX_Datapath/RegisterFile/N25327 ) );
  AOI22_X1 U83020 ( .A1(n105622), .A2(n104819), .B1(n81760), .B2(n109110), 
        .ZN(n96006) );
  OAI21_X1 U83021 ( .B1(n81415), .B2(n105921), .A(n96007), .ZN(
        \DLX_Datapath/RegisterFile/N25326 ) );
  AOI22_X1 U83022 ( .A1(n105621), .A2(n81759), .B1(n105920), .B2(n108645), 
        .ZN(n96007) );
  OAI21_X1 U83023 ( .B1(n106054), .B2(n105922), .A(n96008), .ZN(
        \DLX_Datapath/RegisterFile/N25325 ) );
  AOI22_X1 U83024 ( .A1(n105911), .A2(n104719), .B1(n81760), .B2(n108872), 
        .ZN(n96008) );
  OAI21_X1 U83025 ( .B1(n106269), .B2(n105921), .A(n96009), .ZN(
        \DLX_Datapath/RegisterFile/N25323 ) );
  AOI22_X1 U83026 ( .A1(n81759), .A2(n81265), .B1(n105919), .B2(n107300), .ZN(
        n96009) );
  AOI21_X1 U83027 ( .B1(n96010), .B2(n94258), .A(n96011), .ZN(n81760) );
  NOR2_X1 U83028 ( .A1(n96012), .A2(n96013), .ZN(n81759) );
  OR2_X1 U83029 ( .A1(n96011), .A2(n94999), .ZN(n96012) );
  NOR2_X1 U83030 ( .A1(n81757), .A2(n105089), .ZN(n96011) );
  NAND2_X1 U83031 ( .A1(n105132), .A2(n94934), .ZN(n81757) );
  OAI21_X1 U83032 ( .B1(n81358), .B2(n105450), .A(n96016), .ZN(
        \DLX_Datapath/RegisterFile/N25322 ) );
  AOI22_X1 U83033 ( .A1(n105449), .A2(n70308), .B1(n105447), .B2(n94559), .ZN(
        n96016) );
  OAI21_X1 U83034 ( .B1(n105970), .B2(n105450), .A(n96019), .ZN(
        \DLX_Datapath/RegisterFile/N25321 ) );
  AOI22_X1 U83035 ( .A1(n105449), .A2(n70450), .B1(n105447), .B2(n94562), .ZN(
        n96019) );
  OAI21_X1 U83036 ( .B1(n106135), .B2(n105450), .A(n96020), .ZN(
        \DLX_Datapath/RegisterFile/N25320 ) );
  AOI22_X1 U83037 ( .A1(n105449), .A2(n69503), .B1(n105447), .B2(n94564), .ZN(
        n96020) );
  OAI21_X1 U83038 ( .B1(n106209), .B2(n105450), .A(n96021), .ZN(
        \DLX_Datapath/RegisterFile/N25319 ) );
  AOI22_X1 U83039 ( .A1(n105449), .A2(n107765), .B1(n105447), .B2(n94566), 
        .ZN(n96021) );
  OAI21_X1 U83040 ( .B1(n81306), .B2(n105450), .A(n96022), .ZN(
        \DLX_Datapath/RegisterFile/N25318 ) );
  AOI22_X1 U83041 ( .A1(n105449), .A2(n110668), .B1(n105447), .B2(n94568), 
        .ZN(n96022) );
  OAI21_X1 U83042 ( .B1(n81408), .B2(n105450), .A(n96023), .ZN(
        \DLX_Datapath/RegisterFile/N25317 ) );
  AOI22_X1 U83043 ( .A1(n105449), .A2(n108067), .B1(n105447), .B2(n94570), 
        .ZN(n96023) );
  OAI21_X1 U83044 ( .B1(n81270), .B2(n105450), .A(n96024), .ZN(
        \DLX_Datapath/RegisterFile/N25316 ) );
  AOI22_X1 U83045 ( .A1(n105449), .A2(n110765), .B1(n105447), .B2(n94572), 
        .ZN(n96024) );
  OAI21_X1 U83046 ( .B1(n105991), .B2(n105450), .A(n96025), .ZN(
        \DLX_Datapath/RegisterFile/N25315 ) );
  AOI22_X1 U83047 ( .A1(n105449), .A2(n110866), .B1(n105447), .B2(n94574), 
        .ZN(n96025) );
  OAI21_X1 U83048 ( .B1(n106331), .B2(n105450), .A(n96026), .ZN(
        \DLX_Datapath/RegisterFile/N25314 ) );
  AOI22_X1 U83049 ( .A1(n105448), .A2(n110461), .B1(n105446), .B2(n94576), 
        .ZN(n96026) );
  OAI21_X1 U83050 ( .B1(n106193), .B2(n105450), .A(n96027), .ZN(
        \DLX_Datapath/RegisterFile/N25313 ) );
  AOI22_X1 U83051 ( .A1(n105448), .A2(n110243), .B1(n105446), .B2(n94578), 
        .ZN(n96027) );
  OAI21_X1 U83052 ( .B1(n106128), .B2(n105450), .A(n96028), .ZN(
        \DLX_Datapath/RegisterFile/N25312 ) );
  AOI22_X1 U83053 ( .A1(n105448), .A2(n110560), .B1(n105446), .B2(n94580), 
        .ZN(n96028) );
  OAI21_X1 U83054 ( .B1(n106185), .B2(n105450), .A(n96029), .ZN(
        \DLX_Datapath/RegisterFile/N25311 ) );
  AOI22_X1 U83055 ( .A1(n105448), .A2(n110351), .B1(n105446), .B2(n94582), 
        .ZN(n96029) );
  OAI21_X1 U83056 ( .B1(n81345), .B2(n105450), .A(n96030), .ZN(
        \DLX_Datapath/RegisterFile/N25310 ) );
  AOI22_X1 U83057 ( .A1(n105448), .A2(n110026), .B1(n105446), .B2(n94584), 
        .ZN(n96030) );
  OAI21_X1 U83058 ( .B1(n81403), .B2(n105450), .A(n96031), .ZN(
        \DLX_Datapath/RegisterFile/N25309 ) );
  AOI22_X1 U83059 ( .A1(n105448), .A2(n110133), .B1(n105446), .B2(n94586), 
        .ZN(n96031) );
  OAI21_X1 U83060 ( .B1(n81294), .B2(n105450), .A(n96032), .ZN(
        \DLX_Datapath/RegisterFile/N25308 ) );
  AOI22_X1 U83061 ( .A1(n105448), .A2(n109917), .B1(n105446), .B2(n94588), 
        .ZN(n96032) );
  OAI21_X1 U83062 ( .B1(n106108), .B2(n105450), .A(n96033), .ZN(
        \DLX_Datapath/RegisterFile/N25307 ) );
  AOI22_X1 U83063 ( .A1(n105448), .A2(n109799), .B1(n105446), .B2(n94590), 
        .ZN(n96033) );
  OAI21_X1 U83064 ( .B1(n81284), .B2(n105450), .A(n96034), .ZN(
        \DLX_Datapath/RegisterFile/N25306 ) );
  AOI22_X1 U83065 ( .A1(n105448), .A2(n108173), .B1(n105446), .B2(n94592), 
        .ZN(n96034) );
  OAI21_X1 U83066 ( .B1(n106171), .B2(n105450), .A(n96035), .ZN(
        \DLX_Datapath/RegisterFile/N25305 ) );
  AOI22_X1 U83067 ( .A1(n96017), .A2(n108296), .B1(n105446), .B2(n94594), .ZN(
        n96035) );
  OAI21_X1 U83068 ( .B1(n106236), .B2(n105450), .A(n96036), .ZN(
        \DLX_Datapath/RegisterFile/N25304 ) );
  AOI22_X1 U83069 ( .A1(n96017), .A2(n108407), .B1(n105446), .B2(n94596), .ZN(
        n96036) );
  OAI21_X1 U83070 ( .B1(n106072), .B2(n105450), .A(n96037), .ZN(
        \DLX_Datapath/RegisterFile/N25303 ) );
  AOI22_X1 U83071 ( .A1(n96017), .A2(n107645), .B1(n105446), .B2(n94598), .ZN(
        n96037) );
  OAI21_X1 U83072 ( .B1(n81310), .B2(n105450), .A(n96038), .ZN(
        \DLX_Datapath/RegisterFile/N25302 ) );
  AOI22_X1 U83073 ( .A1(n105448), .A2(n109563), .B1(n105445), .B2(n94600), 
        .ZN(n96038) );
  OAI21_X1 U83074 ( .B1(n106243), .B2(n105450), .A(n96039), .ZN(
        \DLX_Datapath/RegisterFile/N25301 ) );
  AOI22_X1 U83075 ( .A1(n105448), .A2(n108524), .B1(n105445), .B2(n94602), 
        .ZN(n96039) );
  OAI21_X1 U83076 ( .B1(n81349), .B2(n105450), .A(n96040), .ZN(
        \DLX_Datapath/RegisterFile/N25300 ) );
  AOI22_X1 U83077 ( .A1(n105448), .A2(n109668), .B1(n105445), .B2(n94604), 
        .ZN(n96040) );
  OAI21_X1 U83078 ( .B1(n106113), .B2(n105450), .A(n96041), .ZN(
        \DLX_Datapath/RegisterFile/N25299 ) );
  AOI22_X1 U83079 ( .A1(n105448), .A2(n109452), .B1(n105445), .B2(n94606), 
        .ZN(n96041) );
  OAI21_X1 U83080 ( .B1(n81588), .B2(n105450), .A(n96042), .ZN(
        \DLX_Datapath/RegisterFile/N25298 ) );
  AOI22_X1 U83081 ( .A1(n105448), .A2(n108989), .B1(n105445), .B2(n94608), 
        .ZN(n96042) );
  OAI21_X1 U83082 ( .B1(n106261), .B2(n105450), .A(n96043), .ZN(
        \DLX_Datapath/RegisterFile/N25297 ) );
  AOI22_X1 U83083 ( .A1(n105448), .A2(n109337), .B1(n105445), .B2(n94610), 
        .ZN(n96043) );
  OAI21_X1 U83084 ( .B1(n106043), .B2(n105450), .A(n96044), .ZN(
        \DLX_Datapath/RegisterFile/N25296 ) );
  AOI22_X1 U83085 ( .A1(n105448), .A2(n109219), .B1(n105445), .B2(n94612), 
        .ZN(n96044) );
  OAI21_X1 U83086 ( .B1(n106048), .B2(n105450), .A(n96045), .ZN(
        \DLX_Datapath/RegisterFile/N25295 ) );
  AOI22_X1 U83087 ( .A1(n105448), .A2(n109111), .B1(n105445), .B2(n94614), 
        .ZN(n96045) );
  OAI21_X1 U83088 ( .B1(n81415), .B2(n105450), .A(n96046), .ZN(
        \DLX_Datapath/RegisterFile/N25294 ) );
  AOI22_X1 U83089 ( .A1(n105448), .A2(n108646), .B1(n105445), .B2(n94616), 
        .ZN(n96046) );
  OAI21_X1 U83090 ( .B1(n81498), .B2(n105450), .A(n96047), .ZN(
        \DLX_Datapath/RegisterFile/N25293 ) );
  AOI22_X1 U83091 ( .A1(n105448), .A2(n108873), .B1(n105445), .B2(n94618), 
        .ZN(n96047) );
  OAI21_X1 U83092 ( .B1(n105215), .B2(n105450), .A(n96048), .ZN(
        \DLX_Datapath/RegisterFile/N25292 ) );
  AOI22_X1 U83093 ( .A1(n105448), .A2(n108761), .B1(n105445), .B2(n94620), 
        .ZN(n96048) );
  OAI21_X1 U83094 ( .B1(n106266), .B2(n105450), .A(n96049), .ZN(
        \DLX_Datapath/RegisterFile/N25291 ) );
  AOI22_X1 U83095 ( .A1(n105448), .A2(n107301), .B1(n105445), .B2(n94622), 
        .ZN(n96049) );
  OR2_X1 U83097 ( .A1(n96051), .A2(n94999), .ZN(n96050) );
  NOR2_X1 U83098 ( .A1(n96052), .A2(n96051), .ZN(n96017) );
  NOR2_X1 U83099 ( .A1(n96015), .A2(n105091), .ZN(n96051) );
  NAND2_X1 U83100 ( .A1(n94296), .A2(n105132), .ZN(n96015) );
  OAI21_X1 U83101 ( .B1(n106149), .B2(n105444), .A(n96054), .ZN(
        \DLX_Datapath/RegisterFile/N25290 ) );
  AOI22_X1 U83102 ( .A1(n104888), .A2(n107868), .B1(n104770), .B2(n81521), 
        .ZN(n96054) );
  OAI21_X1 U83103 ( .B1(n105970), .B2(n105444), .A(n96057), .ZN(
        \DLX_Datapath/RegisterFile/N25289 ) );
  AOI22_X1 U83104 ( .A1(n104889), .A2(n107965), .B1(n104767), .B2(n81653), 
        .ZN(n96057) );
  OAI21_X1 U83105 ( .B1(n106135), .B2(n105444), .A(n96058), .ZN(
        \DLX_Datapath/RegisterFile/N25288 ) );
  AOI22_X1 U83106 ( .A1(n104888), .A2(n107228), .B1(n104768), .B2(n81380), 
        .ZN(n96058) );
  OAI21_X1 U83107 ( .B1(n106210), .B2(n105444), .A(n96059), .ZN(
        \DLX_Datapath/RegisterFile/N25287 ) );
  AOI22_X1 U83108 ( .A1(n104890), .A2(n107766), .B1(n104767), .B2(n81377), 
        .ZN(n96059) );
  OAI21_X1 U83109 ( .B1(n106204), .B2(n105444), .A(n96060), .ZN(
        \DLX_Datapath/RegisterFile/N25286 ) );
  AOI22_X1 U83110 ( .A1(n104888), .A2(n110669), .B1(n104768), .B2(n81428), 
        .ZN(n96060) );
  OAI21_X1 U83111 ( .B1(n106099), .B2(n105444), .A(n96061), .ZN(
        \DLX_Datapath/RegisterFile/N25285 ) );
  AOI22_X1 U83112 ( .A1(n104889), .A2(n108068), .B1(n104769), .B2(n81410), 
        .ZN(n96061) );
  OAI21_X1 U83113 ( .B1(n106257), .B2(n105444), .A(n96062), .ZN(
        \DLX_Datapath/RegisterFile/N25284 ) );
  AOI22_X1 U83114 ( .A1(n104890), .A2(n110766), .B1(n104770), .B2(n81700), 
        .ZN(n96062) );
  OAI21_X1 U83115 ( .B1(n105991), .B2(n105444), .A(n96063), .ZN(
        \DLX_Datapath/RegisterFile/N25283 ) );
  AOI22_X1 U83116 ( .A1(n104889), .A2(n110867), .B1(n104769), .B2(n81632), 
        .ZN(n96063) );
  OAI21_X1 U83117 ( .B1(n80190), .B2(n105444), .A(n96064), .ZN(
        \DLX_Datapath/RegisterFile/N25282 ) );
  AOI22_X1 U83118 ( .A1(n104890), .A2(n110462), .B1(n104767), .B2(n81414), 
        .ZN(n96064) );
  OAI21_X1 U83119 ( .B1(n106191), .B2(n105444), .A(n96065), .ZN(
        \DLX_Datapath/RegisterFile/N25281 ) );
  AOI22_X1 U83120 ( .A1(n104888), .A2(n110244), .B1(n104768), .B2(n81317), 
        .ZN(n96065) );
  OAI21_X1 U83121 ( .B1(n106128), .B2(n105444), .A(n96066), .ZN(
        \DLX_Datapath/RegisterFile/N25280 ) );
  AOI22_X1 U83122 ( .A1(n104889), .A2(n110561), .B1(n104767), .B2(n81386), 
        .ZN(n96066) );
  OAI21_X1 U83123 ( .B1(n106185), .B2(n105444), .A(n96067), .ZN(
        \DLX_Datapath/RegisterFile/N25279 ) );
  AOI22_X1 U83124 ( .A1(n104890), .A2(n110352), .B1(n104768), .B2(n81320), 
        .ZN(n96067) );
  OAI21_X1 U83125 ( .B1(n81345), .B2(n105444), .A(n96068), .ZN(
        \DLX_Datapath/RegisterFile/N25278 ) );
  AOI22_X1 U83126 ( .A1(n104890), .A2(n110027), .B1(n104769), .B2(n81604), 
        .ZN(n96068) );
  OAI21_X1 U83127 ( .B1(n81403), .B2(n105444), .A(n96069), .ZN(
        \DLX_Datapath/RegisterFile/N25277 ) );
  AOI22_X1 U83128 ( .A1(n104888), .A2(n110134), .B1(n104770), .B2(n81405), 
        .ZN(n96069) );
  OAI21_X1 U83129 ( .B1(n81294), .B2(n105444), .A(n96070), .ZN(
        \DLX_Datapath/RegisterFile/N25276 ) );
  AOI22_X1 U83130 ( .A1(n104888), .A2(n109918), .B1(n104769), .B2(n81402), 
        .ZN(n96070) );
  OAI21_X1 U83131 ( .B1(n106108), .B2(n105444), .A(n96071), .ZN(
        \DLX_Datapath/RegisterFile/N25275 ) );
  AOI22_X1 U83132 ( .A1(n104889), .A2(n109800), .B1(n104770), .B2(n81400), 
        .ZN(n96071) );
  OAI21_X1 U83133 ( .B1(n81284), .B2(n105444), .A(n96072), .ZN(
        \DLX_Datapath/RegisterFile/N25274 ) );
  AOI22_X1 U83134 ( .A1(n104890), .A2(n108174), .B1(n104767), .B2(n81332), 
        .ZN(n96072) );
  OAI21_X1 U83135 ( .B1(n106173), .B2(n105444), .A(n96073), .ZN(
        \DLX_Datapath/RegisterFile/N25273 ) );
  AOI22_X1 U83136 ( .A1(n104889), .A2(n108297), .B1(n104768), .B2(n81373), 
        .ZN(n96073) );
  OAI21_X1 U83137 ( .B1(n106236), .B2(n105444), .A(n96074), .ZN(
        \DLX_Datapath/RegisterFile/N25272 ) );
  AOI22_X1 U83138 ( .A1(n104888), .A2(n108408), .B1(n104767), .B2(n81322), 
        .ZN(n96074) );
  OAI21_X1 U83139 ( .B1(n106072), .B2(n105444), .A(n96075), .ZN(
        \DLX_Datapath/RegisterFile/N25271 ) );
  AOI22_X1 U83140 ( .A1(n104889), .A2(n107646), .B1(n104768), .B2(n81506), 
        .ZN(n96075) );
  OAI21_X1 U83141 ( .B1(n106200), .B2(n105444), .A(n96076), .ZN(
        \DLX_Datapath/RegisterFile/N25270 ) );
  AOI22_X1 U83142 ( .A1(n104890), .A2(n109564), .B1(n104767), .B2(n81313), 
        .ZN(n96076) );
  OAI21_X1 U83143 ( .B1(n106246), .B2(n96053), .A(n96077), .ZN(
        \DLX_Datapath/RegisterFile/N25269 ) );
  AOI22_X1 U83144 ( .A1(n104888), .A2(n108525), .B1(n104770), .B2(n81330), 
        .ZN(n96077) );
  OAI21_X1 U83145 ( .B1(n106159), .B2(n96053), .A(n96078), .ZN(
        \DLX_Datapath/RegisterFile/N25268 ) );
  AOI22_X1 U83146 ( .A1(n104889), .A2(n109669), .B1(n104767), .B2(n81425), 
        .ZN(n96078) );
  OAI21_X1 U83147 ( .B1(n81394), .B2(n96053), .A(n96079), .ZN(
        \DLX_Datapath/RegisterFile/N25267 ) );
  AOI22_X1 U83148 ( .A1(n104889), .A2(n109453), .B1(n104768), .B2(n81396), 
        .ZN(n96079) );
  OAI21_X1 U83149 ( .B1(n106010), .B2(n96053), .A(n96080), .ZN(
        \DLX_Datapath/RegisterFile/N25266 ) );
  AOI22_X1 U83150 ( .A1(n104889), .A2(n108990), .B1(n104770), .B2(n81590), 
        .ZN(n96080) );
  OAI21_X1 U83151 ( .B1(n106262), .B2(n96053), .A(n96081), .ZN(
        \DLX_Datapath/RegisterFile/N25265 ) );
  AOI22_X1 U83152 ( .A1(n104890), .A2(n109338), .B1(n104768), .B2(n81423), 
        .ZN(n96081) );
  OAI21_X1 U83153 ( .B1(n106043), .B2(n96053), .A(n96082), .ZN(
        \DLX_Datapath/RegisterFile/N25264 ) );
  AOI22_X1 U83154 ( .A1(n104890), .A2(n109220), .B1(n104769), .B2(n81511), 
        .ZN(n96082) );
  OAI21_X1 U83155 ( .B1(n106048), .B2(n96053), .A(n96083), .ZN(
        \DLX_Datapath/RegisterFile/N25263 ) );
  AOI22_X1 U83156 ( .A1(n104888), .A2(n109112), .B1(n104769), .B2(n81503), 
        .ZN(n96083) );
  OAI21_X1 U83157 ( .B1(n106094), .B2(n96053), .A(n96084), .ZN(
        \DLX_Datapath/RegisterFile/N25262 ) );
  AOI22_X1 U83158 ( .A1(n104888), .A2(n108647), .B1(n104770), .B2(n81417), 
        .ZN(n96084) );
  OAI21_X1 U83159 ( .B1(n106056), .B2(n96053), .A(n96085), .ZN(
        \DLX_Datapath/RegisterFile/N25261 ) );
  AOI22_X1 U83160 ( .A1(n104890), .A2(n108874), .B1(n104769), .B2(n81500), 
        .ZN(n96085) );
  OAI21_X1 U83161 ( .B1(n105219), .B2(n96053), .A(n96086), .ZN(
        \DLX_Datapath/RegisterFile/N25260 ) );
  AOI22_X1 U83162 ( .A1(n104888), .A2(n108762), .B1(n104769), .B2(n81335), 
        .ZN(n96086) );
  OAI21_X1 U83163 ( .B1(n106268), .B2(n105444), .A(n96087), .ZN(
        \DLX_Datapath/RegisterFile/N25259 ) );
  AOI22_X1 U83164 ( .A1(n104889), .A2(n107302), .B1(n104770), .B2(n81327), 
        .ZN(n96087) );
  NOR2_X1 U83165 ( .A1(n96088), .A2(n96013), .ZN(n96056) );
  OR2_X1 U83166 ( .A1(n96089), .A2(n94999), .ZN(n96088) );
  AOI21_X1 U83168 ( .B1(n105199), .B2(n96090), .A(n94663), .ZN(n96052) );
  OR2_X1 U83169 ( .A1(n94999), .A2(n96013), .ZN(n96090) );
  NOR2_X1 U83170 ( .A1(n96053), .A2(n105089), .ZN(n96089) );
  NAND2_X1 U83171 ( .A1(n105131), .A2(n94331), .ZN(n96053) );
  OAI21_X1 U83172 ( .B1(n102174), .B2(n96091), .A(n96092), .ZN(
        \DLX_Datapath/RegisterFile/N25258 ) );
  AOI22_X1 U83173 ( .A1(n96093), .A2(n106150), .B1(n105440), .B2(n94667), .ZN(
        n96092) );
  OAI21_X1 U83174 ( .B1(n102160), .B2(n96091), .A(n96095), .ZN(
        \DLX_Datapath/RegisterFile/N25257 ) );
  AOI22_X1 U83175 ( .A1(n96093), .A2(n105972), .B1(n105438), .B2(n94670), .ZN(
        n96095) );
  OAI21_X1 U83176 ( .B1(n102145), .B2(n96091), .A(n96096), .ZN(
        \DLX_Datapath/RegisterFile/N25256 ) );
  AOI22_X1 U83177 ( .A1(n105441), .A2(n106139), .B1(n105440), .B2(n94672), 
        .ZN(n96096) );
  OAI21_X1 U83178 ( .B1(n102131), .B2(n96091), .A(n96097), .ZN(
        \DLX_Datapath/RegisterFile/N25255 ) );
  AOI22_X1 U83179 ( .A1(n96093), .A2(n106212), .B1(n105438), .B2(n94674), .ZN(
        n96097) );
  OAI21_X1 U83180 ( .B1(n102115), .B2(n96091), .A(n96098), .ZN(
        \DLX_Datapath/RegisterFile/N25254 ) );
  AOI22_X1 U83181 ( .A1(n96093), .A2(n106207), .B1(n105440), .B2(n94676), .ZN(
        n96098) );
  OAI21_X1 U83182 ( .B1(n102101), .B2(n96091), .A(n96099), .ZN(
        \DLX_Datapath/RegisterFile/N25253 ) );
  AOI22_X1 U83183 ( .A1(n96093), .A2(n106102), .B1(n105438), .B2(n94678), .ZN(
        n96099) );
  OAI21_X1 U83184 ( .B1(n102087), .B2(n96091), .A(n96100), .ZN(
        \DLX_Datapath/RegisterFile/N25252 ) );
  AOI22_X1 U83185 ( .A1(n96093), .A2(n106258), .B1(n105440), .B2(n94680), .ZN(
        n96100) );
  OAI21_X1 U83186 ( .B1(n102070), .B2(n96091), .A(n96101), .ZN(
        \DLX_Datapath/RegisterFile/N25251 ) );
  AOI22_X1 U83187 ( .A1(n96093), .A2(n105993), .B1(n105438), .B2(n94682), .ZN(
        n96101) );
  OAI21_X1 U83188 ( .B1(n102052), .B2(n105443), .A(n96102), .ZN(
        \DLX_Datapath/RegisterFile/N25250 ) );
  AOI22_X1 U83189 ( .A1(n105441), .A2(n106334), .B1(n105439), .B2(n94684), 
        .ZN(n96102) );
  OAI21_X1 U83190 ( .B1(n102036), .B2(n105443), .A(n96103), .ZN(
        \DLX_Datapath/RegisterFile/N25249 ) );
  AOI22_X1 U83191 ( .A1(n105441), .A2(n106194), .B1(n105439), .B2(n94686), 
        .ZN(n96103) );
  OAI21_X1 U83192 ( .B1(n102019), .B2(n105443), .A(n96104), .ZN(
        \DLX_Datapath/RegisterFile/N25248 ) );
  AOI22_X1 U83193 ( .A1(n105441), .A2(n106132), .B1(n105439), .B2(n94688), 
        .ZN(n96104) );
  OAI21_X1 U83194 ( .B1(n102001), .B2(n105443), .A(n96105), .ZN(
        \DLX_Datapath/RegisterFile/N25247 ) );
  AOI22_X1 U83195 ( .A1(n105441), .A2(n106189), .B1(n105439), .B2(n94690), 
        .ZN(n96105) );
  OAI21_X1 U83196 ( .B1(n101985), .B2(n105443), .A(n96106), .ZN(
        \DLX_Datapath/RegisterFile/N25246 ) );
  AOI22_X1 U83197 ( .A1(n105441), .A2(n106166), .B1(n105439), .B2(n94692), 
        .ZN(n96106) );
  OAI21_X1 U83198 ( .B1(n101969), .B2(n105443), .A(n96107), .ZN(
        \DLX_Datapath/RegisterFile/N25245 ) );
  AOI22_X1 U83199 ( .A1(n105441), .A2(n106107), .B1(n105439), .B2(n94694), 
        .ZN(n96107) );
  OAI21_X1 U83200 ( .B1(n101953), .B2(n105443), .A(n96108), .ZN(
        \DLX_Datapath/RegisterFile/N25244 ) );
  AOI22_X1 U83201 ( .A1(n105441), .A2(n106222), .B1(n105439), .B2(n94696), 
        .ZN(n96108) );
  OAI21_X1 U83202 ( .B1(n101937), .B2(n105443), .A(n96109), .ZN(
        \DLX_Datapath/RegisterFile/N25243 ) );
  AOI22_X1 U83203 ( .A1(n105441), .A2(n106112), .B1(n105439), .B2(n94698), 
        .ZN(n96109) );
  OAI21_X1 U83204 ( .B1(n101921), .B2(n105443), .A(n96110), .ZN(
        \DLX_Datapath/RegisterFile/N25242 ) );
  AOI22_X1 U83205 ( .A1(n105441), .A2(n106234), .B1(n105439), .B2(n94700), 
        .ZN(n96110) );
  OAI21_X1 U83206 ( .B1(n101905), .B2(n105443), .A(n96111), .ZN(
        \DLX_Datapath/RegisterFile/N25241 ) );
  AOI22_X1 U83207 ( .A1(n105441), .A2(n106174), .B1(n105439), .B2(n94702), 
        .ZN(n96111) );
  OAI21_X1 U83208 ( .B1(n101889), .B2(n105443), .A(n96112), .ZN(
        \DLX_Datapath/RegisterFile/N25240 ) );
  AOI22_X1 U83209 ( .A1(n105441), .A2(n106239), .B1(n105439), .B2(n94704), 
        .ZN(n96112) );
  OAI21_X1 U83210 ( .B1(n101871), .B2(n105443), .A(n96113), .ZN(
        \DLX_Datapath/RegisterFile/N25239 ) );
  AOI22_X1 U83211 ( .A1(n105441), .A2(n106073), .B1(n105438), .B2(n94706), 
        .ZN(n96113) );
  OAI21_X1 U83212 ( .B1(n101855), .B2(n105442), .A(n96114), .ZN(
        \DLX_Datapath/RegisterFile/N25238 ) );
  AOI22_X1 U83213 ( .A1(n105441), .A2(n106201), .B1(n105440), .B2(n94708), 
        .ZN(n96114) );
  OAI21_X1 U83214 ( .B1(n101837), .B2(n105442), .A(n96115), .ZN(
        \DLX_Datapath/RegisterFile/N25237 ) );
  AOI22_X1 U83215 ( .A1(n105441), .A2(n106247), .B1(n105438), .B2(n94710), 
        .ZN(n96115) );
  OAI21_X1 U83216 ( .B1(n101819), .B2(n105442), .A(n96116), .ZN(
        \DLX_Datapath/RegisterFile/N25236 ) );
  AOI22_X1 U83217 ( .A1(n105441), .A2(n106161), .B1(n105440), .B2(n94712), 
        .ZN(n96116) );
  OAI21_X1 U83218 ( .B1(n101803), .B2(n105442), .A(n96117), .ZN(
        \DLX_Datapath/RegisterFile/N25235 ) );
  AOI22_X1 U83219 ( .A1(n105441), .A2(n106117), .B1(n105438), .B2(n94714), 
        .ZN(n96117) );
  OAI21_X1 U83220 ( .B1(n101785), .B2(n105442), .A(n96118), .ZN(
        \DLX_Datapath/RegisterFile/N25234 ) );
  AOI22_X1 U83221 ( .A1(n96093), .A2(n106012), .B1(n105440), .B2(n81259), .ZN(
        n96118) );
  OAI21_X1 U83222 ( .B1(n101769), .B2(n105442), .A(n96119), .ZN(
        \DLX_Datapath/RegisterFile/N25233 ) );
  AOI22_X1 U83223 ( .A1(n96093), .A2(n106263), .B1(n105438), .B2(n94717), .ZN(
        n96119) );
  OAI21_X1 U83224 ( .B1(n101751), .B2(n105442), .A(n96120), .ZN(
        \DLX_Datapath/RegisterFile/N25232 ) );
  AOI22_X1 U83225 ( .A1(n96093), .A2(n106047), .B1(n105440), .B2(n94719), .ZN(
        n96120) );
  OAI21_X1 U83226 ( .B1(n101733), .B2(n105442), .A(n96121), .ZN(
        \DLX_Datapath/RegisterFile/N25231 ) );
  AOI22_X1 U83227 ( .A1(n105441), .A2(n106052), .B1(n105438), .B2(n94721), 
        .ZN(n96121) );
  OAI21_X1 U83228 ( .B1(n101715), .B2(n105442), .A(n96122), .ZN(
        \DLX_Datapath/RegisterFile/N25230 ) );
  AOI22_X1 U83229 ( .A1(n105441), .A2(n106097), .B1(n105440), .B2(n94723), 
        .ZN(n96122) );
  OAI21_X1 U83230 ( .B1(n101697), .B2(n105442), .A(n96123), .ZN(
        \DLX_Datapath/RegisterFile/N25229 ) );
  AOI22_X1 U83231 ( .A1(n96093), .A2(n106057), .B1(n105438), .B2(n94725), .ZN(
        n96123) );
  OAI21_X1 U83232 ( .B1(n101679), .B2(n105442), .A(n96124), .ZN(
        \DLX_Datapath/RegisterFile/N25228 ) );
  AOI22_X1 U83233 ( .A1(n105441), .A2(n96125), .B1(n105440), .B2(n94727), .ZN(
        n96124) );
  OAI21_X1 U83234 ( .B1(n101661), .B2(n105442), .A(n96126), .ZN(
        \DLX_Datapath/RegisterFile/N25227 ) );
  AOI22_X1 U83235 ( .A1(n105441), .A2(n106270), .B1(n105438), .B2(n94729), 
        .ZN(n96126) );
  NAND2_X1 U83237 ( .A1(n96128), .A2(n111025), .ZN(n96127) );
  OAI21_X1 U83238 ( .B1(n96129), .B2(n94663), .A(n96128), .ZN(n96091) );
  NAND2_X1 U83239 ( .A1(n96093), .A2(n105502), .ZN(n96128) );
  AND2_X2 U83240 ( .A1(n94367), .A2(n105131), .ZN(n96093) );
  AOI21_X1 U83241 ( .B1(n96130), .B2(n111025), .A(n94366), .ZN(n96129) );
  OAI21_X1 U83242 ( .B1(n106149), .B2(n105437), .A(n96132), .ZN(
        \DLX_Datapath/RegisterFile/N25226 ) );
  AOI22_X1 U83243 ( .A1(n104987), .A2(n107870), .B1(n105436), .B2(n81360), 
        .ZN(n96132) );
  OAI21_X1 U83244 ( .B1(n105970), .B2(n105437), .A(n96135), .ZN(
        \DLX_Datapath/RegisterFile/N25225 ) );
  AOI22_X1 U83245 ( .A1(n104988), .A2(n107967), .B1(n105435), .B2(n94511), 
        .ZN(n96135) );
  OAI21_X1 U83246 ( .B1(n106135), .B2(n105437), .A(n96136), .ZN(
        \DLX_Datapath/RegisterFile/N25224 ) );
  AOI22_X1 U83247 ( .A1(n104987), .A2(n107230), .B1(n105435), .B2(n81539), 
        .ZN(n96136) );
  OAI21_X1 U83248 ( .B1(n106211), .B2(n105437), .A(n96137), .ZN(
        \DLX_Datapath/RegisterFile/N25223 ) );
  AOI22_X1 U83249 ( .A1(n104988), .A2(n107768), .B1(n105436), .B2(n81301), 
        .ZN(n96137) );
  OAI21_X1 U83250 ( .B1(n106204), .B2(n105437), .A(n96138), .ZN(
        \DLX_Datapath/RegisterFile/N25222 ) );
  AOI22_X1 U83251 ( .A1(n104989), .A2(n110671), .B1(n105435), .B2(n81308), 
        .ZN(n96138) );
  OAI21_X1 U83252 ( .B1(n106101), .B2(n105437), .A(n96139), .ZN(
        \DLX_Datapath/RegisterFile/N25221 ) );
  AOI22_X1 U83253 ( .A1(n104988), .A2(n108070), .B1(n105436), .B2(n94516), 
        .ZN(n96139) );
  OAI21_X1 U83254 ( .B1(n81270), .B2(n105437), .A(n96140), .ZN(
        \DLX_Datapath/RegisterFile/N25220 ) );
  AOI22_X1 U83255 ( .A1(n104987), .A2(n110768), .B1(n105436), .B2(n81272), 
        .ZN(n96140) );
  OAI21_X1 U83256 ( .B1(n105991), .B2(n105437), .A(n96141), .ZN(
        \DLX_Datapath/RegisterFile/N25219 ) );
  AOI22_X1 U83257 ( .A1(n104989), .A2(n110869), .B1(n105435), .B2(n94519), 
        .ZN(n96141) );
  OAI21_X1 U83258 ( .B1(n80190), .B2(n105437), .A(n96142), .ZN(
        \DLX_Datapath/RegisterFile/N25218 ) );
  AOI22_X1 U83259 ( .A1(n104988), .A2(n110464), .B1(n105435), .B2(n80192), 
        .ZN(n96142) );
  OAI21_X1 U83260 ( .B1(n106190), .B2(n105437), .A(n96143), .ZN(
        \DLX_Datapath/RegisterFile/N25217 ) );
  AOI22_X1 U83261 ( .A1(n104987), .A2(n110246), .B1(n105434), .B2(n81474), 
        .ZN(n96143) );
  OAI21_X1 U83262 ( .B1(n106128), .B2(n105437), .A(n96144), .ZN(
        \DLX_Datapath/RegisterFile/N25216 ) );
  AOI22_X1 U83263 ( .A1(n104988), .A2(n110563), .B1(n105434), .B2(n94523), 
        .ZN(n96144) );
  OAI21_X1 U83264 ( .B1(n106185), .B2(n105437), .A(n96145), .ZN(
        \DLX_Datapath/RegisterFile/N25215 ) );
  AOI22_X1 U83265 ( .A1(n104989), .A2(n110354), .B1(n105434), .B2(n106061), 
        .ZN(n96145) );
  OAI21_X1 U83266 ( .B1(n81345), .B2(n105437), .A(n96146), .ZN(
        \DLX_Datapath/RegisterFile/N25214 ) );
  AOI22_X1 U83267 ( .A1(n104989), .A2(n110029), .B1(n105434), .B2(n81347), 
        .ZN(n96146) );
  OAI21_X1 U83268 ( .B1(n81403), .B2(n105437), .A(n96147), .ZN(
        \DLX_Datapath/RegisterFile/N25213 ) );
  AOI22_X1 U83269 ( .A1(n104987), .A2(n110136), .B1(n105434), .B2(n94527), 
        .ZN(n96147) );
  OAI21_X1 U83270 ( .B1(n106218), .B2(n105437), .A(n96148), .ZN(
        \DLX_Datapath/RegisterFile/N25212 ) );
  AOI22_X1 U83271 ( .A1(n104987), .A2(n109920), .B1(n105434), .B2(n81297), 
        .ZN(n96148) );
  OAI21_X1 U83272 ( .B1(n106108), .B2(n105437), .A(n96149), .ZN(
        \DLX_Datapath/RegisterFile/N25211 ) );
  AOI22_X1 U83273 ( .A1(n104988), .A2(n109802), .B1(n105436), .B2(n94530), 
        .ZN(n96149) );
  OAI21_X1 U83274 ( .B1(n81284), .B2(n105437), .A(n96150), .ZN(
        \DLX_Datapath/RegisterFile/N25210 ) );
  AOI22_X1 U83275 ( .A1(n104989), .A2(n108176), .B1(n105434), .B2(n81286), 
        .ZN(n96150) );
  OAI21_X1 U83276 ( .B1(n106171), .B2(n105437), .A(n96151), .ZN(
        \DLX_Datapath/RegisterFile/N25209 ) );
  AOI22_X1 U83277 ( .A1(n104988), .A2(n108299), .B1(n105434), .B2(n106168), 
        .ZN(n96151) );
  OAI21_X1 U83278 ( .B1(n106236), .B2(n105437), .A(n96152), .ZN(
        \DLX_Datapath/RegisterFile/N25208 ) );
  AOI22_X1 U83279 ( .A1(n104987), .A2(n108410), .B1(n105434), .B2(n81283), 
        .ZN(n96152) );
  OAI21_X1 U83280 ( .B1(n106072), .B2(n105437), .A(n96153), .ZN(
        \DLX_Datapath/RegisterFile/N25207 ) );
  AOI22_X1 U83281 ( .A1(n104988), .A2(n107648), .B1(n105434), .B2(n81453), 
        .ZN(n96153) );
  OAI21_X1 U83282 ( .B1(n106198), .B2(n105437), .A(n96154), .ZN(
        \DLX_Datapath/RegisterFile/N25206 ) );
  AOI22_X1 U83283 ( .A1(n104989), .A2(n109566), .B1(n105435), .B2(n94536), 
        .ZN(n96154) );
  OAI21_X1 U83284 ( .B1(n81278), .B2(n105437), .A(n96155), .ZN(
        \DLX_Datapath/RegisterFile/N25205 ) );
  AOI22_X1 U83285 ( .A1(n104989), .A2(n108527), .B1(n105436), .B2(n106241), 
        .ZN(n96155) );
  OAI21_X1 U83286 ( .B1(n106157), .B2(n96131), .A(n96156), .ZN(
        \DLX_Datapath/RegisterFile/N25204 ) );
  AOI22_X1 U83287 ( .A1(n104989), .A2(n109671), .B1(n105435), .B2(n81351), 
        .ZN(n96156) );
  OAI21_X1 U83288 ( .B1(n106113), .B2(n96131), .A(n96157), .ZN(
        \DLX_Datapath/RegisterFile/N25203 ) );
  AOI22_X1 U83289 ( .A1(n104987), .A2(n109455), .B1(n105436), .B2(n106020), 
        .ZN(n96157) );
  OAI21_X1 U83290 ( .B1(n106007), .B2(n96131), .A(n96158), .ZN(
        \DLX_Datapath/RegisterFile/N25202 ) );
  AOI22_X1 U83291 ( .A1(n104987), .A2(n108992), .B1(n105435), .B2(n94541), 
        .ZN(n96158) );
  OAI21_X1 U83292 ( .B1(n81267), .B2(n105437), .A(n96159), .ZN(
        \DLX_Datapath/RegisterFile/N25201 ) );
  AOI22_X1 U83293 ( .A1(n104988), .A2(n109340), .B1(n105435), .B2(n81269), 
        .ZN(n96159) );
  OAI21_X1 U83294 ( .B1(n106043), .B2(n96131), .A(n96160), .ZN(
        \DLX_Datapath/RegisterFile/N25200 ) );
  AOI22_X1 U83295 ( .A1(n104989), .A2(n109222), .B1(n105436), .B2(n105624), 
        .ZN(n96160) );
  OAI21_X1 U83296 ( .B1(n106048), .B2(n96131), .A(n96161), .ZN(
        \DLX_Datapath/RegisterFile/N25199 ) );
  AOI22_X1 U83297 ( .A1(n104988), .A2(n109114), .B1(n105435), .B2(n94546), 
        .ZN(n96161) );
  OAI21_X1 U83298 ( .B1(n106093), .B2(n96131), .A(n96162), .ZN(
        \DLX_Datapath/RegisterFile/N25198 ) );
  AOI22_X1 U83299 ( .A1(n104987), .A2(n108649), .B1(n105436), .B2(n94548), 
        .ZN(n96162) );
  OAI21_X1 U83300 ( .B1(n106055), .B2(n96131), .A(n96163), .ZN(
        \DLX_Datapath/RegisterFile/N25197 ) );
  AOI22_X1 U83301 ( .A1(n104988), .A2(n108876), .B1(n105436), .B2(n81783), 
        .ZN(n96163) );
  OAI21_X1 U83302 ( .B1(n105219), .B2(n96131), .A(n96164), .ZN(
        \DLX_Datapath/RegisterFile/N25196 ) );
  AOI22_X1 U83303 ( .A1(n104987), .A2(n108764), .B1(n105436), .B2(n80188), 
        .ZN(n96164) );
  OAI21_X1 U83304 ( .B1(n81262), .B2(n105437), .A(n96165), .ZN(
        \DLX_Datapath/RegisterFile/N25195 ) );
  AOI22_X1 U83305 ( .A1(n104989), .A2(n107304), .B1(n105435), .B2(n81265), 
        .ZN(n96165) );
  AOI21_X1 U83307 ( .B1(n96010), .B2(n94398), .A(n96167), .ZN(n96133) );
  NOR2_X1 U83308 ( .A1(n96131), .A2(n105090), .ZN(n96167) );
  NAND2_X1 U83309 ( .A1(n105132), .A2(n94399), .ZN(n96131) );
  OAI21_X1 U83310 ( .B1(n106147), .B2(n96168), .A(n96169), .ZN(
        \DLX_Datapath/RegisterFile/N25194 ) );
  AOI22_X1 U83311 ( .A1(n105432), .A2(n70312), .B1(n104974), .B2(n94559), .ZN(
        n96169) );
  OAI21_X1 U83312 ( .B1(n105970), .B2(n96168), .A(n96172), .ZN(
        \DLX_Datapath/RegisterFile/N25193 ) );
  AOI22_X1 U83313 ( .A1(n105431), .A2(n70454), .B1(n104975), .B2(n94562), .ZN(
        n96172) );
  OAI21_X1 U83314 ( .B1(n81378), .B2(n105433), .A(n96173), .ZN(
        \DLX_Datapath/RegisterFile/N25192 ) );
  AOI22_X1 U83315 ( .A1(n105432), .A2(n69507), .B1(n104974), .B2(n94564), .ZN(
        n96173) );
  OAI21_X1 U83316 ( .B1(n106208), .B2(n105433), .A(n96174), .ZN(
        \DLX_Datapath/RegisterFile/N25191 ) );
  AOI22_X1 U83317 ( .A1(n105431), .A2(n70168), .B1(n104976), .B2(n94566), .ZN(
        n96174) );
  OAI21_X1 U83318 ( .B1(n106204), .B2(n96168), .A(n96175), .ZN(
        \DLX_Datapath/RegisterFile/N25190 ) );
  AOI22_X1 U83319 ( .A1(n105432), .A2(n74014), .B1(n104974), .B2(n94568), .ZN(
        n96175) );
  OAI21_X1 U83320 ( .B1(n106100), .B2(n96168), .A(n96176), .ZN(
        \DLX_Datapath/RegisterFile/N25189 ) );
  AOI22_X1 U83321 ( .A1(n105431), .A2(n70601), .B1(n104975), .B2(n94570), .ZN(
        n96176) );
  OAI21_X1 U83322 ( .B1(n81270), .B2(n105433), .A(n96177), .ZN(
        \DLX_Datapath/RegisterFile/N25188 ) );
  AOI22_X1 U83323 ( .A1(n105432), .A2(n74155), .B1(n104975), .B2(n94572), .ZN(
        n96177) );
  OAI21_X1 U83324 ( .B1(n105992), .B2(n105433), .A(n96178), .ZN(
        \DLX_Datapath/RegisterFile/N25187 ) );
  AOI22_X1 U83325 ( .A1(n105431), .A2(n74295), .B1(n104976), .B2(n94574), .ZN(
        n96178) );
  OAI21_X1 U83326 ( .B1(n80190), .B2(n105433), .A(n96179), .ZN(
        \DLX_Datapath/RegisterFile/N25186 ) );
  AOI22_X1 U83327 ( .A1(n105431), .A2(n73731), .B1(n104975), .B2(n94576), .ZN(
        n96179) );
  OAI21_X1 U83328 ( .B1(n106190), .B2(n105433), .A(n96180), .ZN(
        \DLX_Datapath/RegisterFile/N25185 ) );
  AOI22_X1 U83329 ( .A1(n105430), .A2(n73435), .B1(n104974), .B2(n94578), .ZN(
        n96180) );
  OAI21_X1 U83330 ( .B1(n106128), .B2(n105433), .A(n96181), .ZN(
        \DLX_Datapath/RegisterFile/N25184 ) );
  AOI22_X1 U83331 ( .A1(n105430), .A2(n73872), .B1(n104975), .B2(n94580), .ZN(
        n96181) );
  OAI21_X1 U83332 ( .B1(n106185), .B2(n105433), .A(n96182), .ZN(
        \DLX_Datapath/RegisterFile/N25183 ) );
  AOI22_X1 U83333 ( .A1(n105430), .A2(n73584), .B1(n104976), .B2(n94582), .ZN(
        n96182) );
  OAI21_X1 U83334 ( .B1(n81345), .B2(n105433), .A(n96183), .ZN(
        \DLX_Datapath/RegisterFile/N25182 ) );
  AOI22_X1 U83335 ( .A1(n105430), .A2(n73146), .B1(n104976), .B2(n94584), .ZN(
        n96183) );
  OAI21_X1 U83336 ( .B1(n81403), .B2(n105433), .A(n96184), .ZN(
        \DLX_Datapath/RegisterFile/N25181 ) );
  AOI22_X1 U83337 ( .A1(n105430), .A2(n73288), .B1(n104974), .B2(n94586), .ZN(
        n96184) );
  OAI21_X1 U83338 ( .B1(n81294), .B2(n105433), .A(n96185), .ZN(
        \DLX_Datapath/RegisterFile/N25180 ) );
  AOI22_X1 U83339 ( .A1(n105430), .A2(n73004), .B1(n104974), .B2(n94588), .ZN(
        n96185) );
  OAI21_X1 U83340 ( .B1(n106108), .B2(n105433), .A(n96186), .ZN(
        \DLX_Datapath/RegisterFile/N25179 ) );
  AOI22_X1 U83341 ( .A1(n105430), .A2(n72854), .B1(n104975), .B2(n94590), .ZN(
        n96186) );
  OAI21_X1 U83342 ( .B1(n81284), .B2(n105433), .A(n96187), .ZN(
        \DLX_Datapath/RegisterFile/N25178 ) );
  AOI22_X1 U83343 ( .A1(n105430), .A2(n70750), .B1(n104976), .B2(n94592), .ZN(
        n96187) );
  OAI21_X1 U83344 ( .B1(n106171), .B2(n105433), .A(n96188), .ZN(
        \DLX_Datapath/RegisterFile/N25177 ) );
  AOI22_X1 U83345 ( .A1(n105430), .A2(n70909), .B1(n104975), .B2(n94594), .ZN(
        n96188) );
  OAI21_X1 U83346 ( .B1(n106236), .B2(n105433), .A(n96189), .ZN(
        \DLX_Datapath/RegisterFile/N25176 ) );
  AOI22_X1 U83347 ( .A1(n105430), .A2(n71054), .B1(n104974), .B2(n94596), .ZN(
        n96189) );
  OAI21_X1 U83348 ( .B1(n106072), .B2(n105433), .A(n96190), .ZN(
        \DLX_Datapath/RegisterFile/N25175 ) );
  AOI22_X1 U83349 ( .A1(n105430), .A2(n70015), .B1(n104975), .B2(n94598), .ZN(
        n96190) );
  OAI21_X1 U83350 ( .B1(n106198), .B2(n105433), .A(n96191), .ZN(
        \DLX_Datapath/RegisterFile/N25174 ) );
  AOI22_X1 U83351 ( .A1(n105431), .A2(n72544), .B1(n104976), .B2(n94600), .ZN(
        n96191) );
  OAI21_X1 U83352 ( .B1(n81278), .B2(n105433), .A(n96192), .ZN(
        \DLX_Datapath/RegisterFile/N25173 ) );
  AOI22_X1 U83353 ( .A1(n105432), .A2(n71203), .B1(n104976), .B2(n94602), .ZN(
        n96192) );
  OAI21_X1 U83354 ( .B1(n106157), .B2(n105433), .A(n96193), .ZN(
        \DLX_Datapath/RegisterFile/N25172 ) );
  AOI22_X1 U83355 ( .A1(n105431), .A2(n72686), .B1(n104976), .B2(n94604), .ZN(
        n96193) );
  OAI21_X1 U83356 ( .B1(n106114), .B2(n96168), .A(n96194), .ZN(
        \DLX_Datapath/RegisterFile/N25171 ) );
  AOI22_X1 U83357 ( .A1(n105432), .A2(n72396), .B1(n104974), .B2(n94606), .ZN(
        n96194) );
  OAI21_X1 U83358 ( .B1(n106008), .B2(n105433), .A(n96195), .ZN(
        \DLX_Datapath/RegisterFile/N25170 ) );
  AOI22_X1 U83359 ( .A1(n105431), .A2(n71796), .B1(n104974), .B2(n94608), .ZN(
        n96195) );
  OAI21_X1 U83360 ( .B1(n106262), .B2(n96168), .A(n96196), .ZN(
        \DLX_Datapath/RegisterFile/N25169 ) );
  AOI22_X1 U83361 ( .A1(n105432), .A2(n72245), .B1(n104975), .B2(n94610), .ZN(
        n96196) );
  OAI21_X1 U83362 ( .B1(n106043), .B2(n105433), .A(n96197), .ZN(
        \DLX_Datapath/RegisterFile/N25168 ) );
  AOI22_X1 U83363 ( .A1(n105431), .A2(n72094), .B1(n104976), .B2(n94612), .ZN(
        n96197) );
  OAI21_X1 U83364 ( .B1(n106049), .B2(n96168), .A(n96198), .ZN(
        \DLX_Datapath/RegisterFile/N25167 ) );
  AOI22_X1 U83365 ( .A1(n105432), .A2(n71950), .B1(n104975), .B2(n94614), .ZN(
        n96198) );
  OAI21_X1 U83366 ( .B1(n106095), .B2(n96168), .A(n96199), .ZN(
        \DLX_Datapath/RegisterFile/N25166 ) );
  AOI22_X1 U83367 ( .A1(n105431), .A2(n71352), .B1(n104974), .B2(n94616), .ZN(
        n96199) );
  OAI21_X1 U83368 ( .B1(n106053), .B2(n105433), .A(n96200), .ZN(
        \DLX_Datapath/RegisterFile/N25165 ) );
  AOI22_X1 U83369 ( .A1(n105432), .A2(n71647), .B1(n104975), .B2(n94618), .ZN(
        n96200) );
  OAI21_X1 U83370 ( .B1(n105219), .B2(n105433), .A(n96201), .ZN(
        \DLX_Datapath/RegisterFile/N25164 ) );
  AOI22_X1 U83371 ( .A1(n105432), .A2(n71503), .B1(n104974), .B2(n94620), .ZN(
        n96201) );
  OAI21_X1 U83372 ( .B1(n81262), .B2(n105433), .A(n96202), .ZN(
        \DLX_Datapath/RegisterFile/N25163 ) );
  AOI22_X1 U83373 ( .A1(n105431), .A2(n69612), .B1(n104976), .B2(n94622), .ZN(
        n96202) );
  NOR2_X1 U83376 ( .A1(n96168), .A2(n105090), .ZN(n96203) );
  NAND2_X1 U83377 ( .A1(n94434), .A2(n105131), .ZN(n96168) );
  OAI21_X1 U83378 ( .B1(n106148), .B2(n81619), .A(n96205), .ZN(
        \DLX_Datapath/RegisterFile/N25162 ) );
  AOI22_X1 U83379 ( .A1(n105999), .A2(n107871), .B1(n105996), .B2(n81521), 
        .ZN(n96205) );
  OAI21_X1 U83380 ( .B1(n81619), .B2(n81651), .A(n96206), .ZN(
        \DLX_Datapath/RegisterFile/N25161 ) );
  AOI22_X1 U83381 ( .A1(n105999), .A2(n107968), .B1(n81653), .B2(n105995), 
        .ZN(n96206) );
  OAI21_X1 U83382 ( .B1(n106136), .B2(n81619), .A(n96207), .ZN(
        \DLX_Datapath/RegisterFile/N25160 ) );
  AOI22_X1 U83383 ( .A1(n105999), .A2(n107231), .B1(n105996), .B2(n81380), 
        .ZN(n96207) );
  OAI21_X1 U83384 ( .B1(n106209), .B2(n81619), .A(n96208), .ZN(
        \DLX_Datapath/RegisterFile/N25159 ) );
  AOI22_X1 U83385 ( .A1(n106000), .A2(n107769), .B1(n105997), .B2(n81377), 
        .ZN(n96208) );
  OAI21_X1 U83386 ( .B1(n106204), .B2(n106001), .A(n96209), .ZN(
        \DLX_Datapath/RegisterFile/N25158 ) );
  AOI22_X1 U83387 ( .A1(n105998), .A2(n110672), .B1(n105995), .B2(n81428), 
        .ZN(n96209) );
  OAI21_X1 U83388 ( .B1(n106098), .B2(n106001), .A(n96210), .ZN(
        \DLX_Datapath/RegisterFile/N25157 ) );
  AOI22_X1 U83389 ( .A1(n105998), .A2(n108071), .B1(n105997), .B2(n81410), 
        .ZN(n96210) );
  OAI21_X1 U83390 ( .B1(n81270), .B2(n106001), .A(n96211), .ZN(
        \DLX_Datapath/RegisterFile/N25156 ) );
  AOI22_X1 U83391 ( .A1(n105998), .A2(n110769), .B1(n81700), .B2(n105995), 
        .ZN(n96211) );
  OAI21_X1 U83392 ( .B1(n81619), .B2(n105991), .A(n96212), .ZN(
        \DLX_Datapath/RegisterFile/N25155 ) );
  AOI22_X1 U83393 ( .A1(n105998), .A2(n110870), .B1(n81632), .B2(n105995), 
        .ZN(n96212) );
  OAI21_X1 U83394 ( .B1(n106330), .B2(n106001), .A(n96213), .ZN(
        \DLX_Datapath/RegisterFile/N25154 ) );
  AOI22_X1 U83395 ( .A1(n105998), .A2(n110465), .B1(n105996), .B2(n81414), 
        .ZN(n96213) );
  OAI21_X1 U83396 ( .B1(n106190), .B2(n106001), .A(n96214), .ZN(
        \DLX_Datapath/RegisterFile/N25153 ) );
  AOI22_X1 U83397 ( .A1(n105998), .A2(n110247), .B1(n105997), .B2(n81317), 
        .ZN(n96214) );
  OAI21_X1 U83398 ( .B1(n106130), .B2(n106001), .A(n96215), .ZN(
        \DLX_Datapath/RegisterFile/N25152 ) );
  AOI22_X1 U83399 ( .A1(n105998), .A2(n110564), .B1(n105995), .B2(n81386), 
        .ZN(n96215) );
  OAI21_X1 U83400 ( .B1(n106185), .B2(n106001), .A(n96216), .ZN(
        \DLX_Datapath/RegisterFile/N25151 ) );
  AOI22_X1 U83401 ( .A1(n105998), .A2(n110355), .B1(n105995), .B2(n81320), 
        .ZN(n96216) );
  OAI21_X1 U83402 ( .B1(n106218), .B2(n106001), .A(n96217), .ZN(
        \DLX_Datapath/RegisterFile/N25148 ) );
  AOI22_X1 U83403 ( .A1(n105998), .A2(n109921), .B1(n105995), .B2(n81402), 
        .ZN(n96217) );
  OAI21_X1 U83404 ( .B1(n106108), .B2(n106001), .A(n96218), .ZN(
        \DLX_Datapath/RegisterFile/N25147 ) );
  AOI22_X1 U83405 ( .A1(n105998), .A2(n109803), .B1(n105995), .B2(n81400), 
        .ZN(n96218) );
  OAI21_X1 U83406 ( .B1(n106236), .B2(n106001), .A(n96219), .ZN(
        \DLX_Datapath/RegisterFile/N25144 ) );
  AOI22_X1 U83407 ( .A1(n106000), .A2(n108411), .B1(n105995), .B2(n81322), 
        .ZN(n96219) );
  OAI21_X1 U83408 ( .B1(n106072), .B2(n106001), .A(n96220), .ZN(
        \DLX_Datapath/RegisterFile/N25143 ) );
  AOI22_X1 U83409 ( .A1(n105999), .A2(n107649), .B1(n105995), .B2(n81506), 
        .ZN(n96220) );
  OAI21_X1 U83410 ( .B1(n106197), .B2(n106001), .A(n96221), .ZN(
        \DLX_Datapath/RegisterFile/N25142 ) );
  AOI22_X1 U83411 ( .A1(n105999), .A2(n109567), .B1(n105996), .B2(n81313), 
        .ZN(n96221) );
  OAI21_X1 U83412 ( .B1(n106115), .B2(n106001), .A(n96222), .ZN(
        \DLX_Datapath/RegisterFile/N25139 ) );
  AOI22_X1 U83413 ( .A1(n106000), .A2(n109456), .B1(n105996), .B2(n81396), 
        .ZN(n96222) );
  OAI21_X1 U83414 ( .B1(n106007), .B2(n106001), .A(n96223), .ZN(
        \DLX_Datapath/RegisterFile/N25138 ) );
  AOI22_X1 U83415 ( .A1(n105999), .A2(n108993), .B1(n105997), .B2(n81590), 
        .ZN(n96223) );
  OAI21_X1 U83416 ( .B1(n106259), .B2(n106001), .A(n96224), .ZN(
        \DLX_Datapath/RegisterFile/N25137 ) );
  AOI22_X1 U83417 ( .A1(n106000), .A2(n109341), .B1(n105996), .B2(n81423), 
        .ZN(n96224) );
  OAI21_X1 U83418 ( .B1(n106043), .B2(n106001), .A(n96225), .ZN(
        \DLX_Datapath/RegisterFile/N25136 ) );
  AOI22_X1 U83419 ( .A1(n105999), .A2(n109223), .B1(n105997), .B2(n81511), 
        .ZN(n96225) );
  OAI21_X1 U83420 ( .B1(n106049), .B2(n106001), .A(n96226), .ZN(
        \DLX_Datapath/RegisterFile/N25135 ) );
  AOI22_X1 U83421 ( .A1(n106000), .A2(n109115), .B1(n105996), .B2(n81503), 
        .ZN(n96226) );
  OAI21_X1 U83422 ( .B1(n106096), .B2(n106001), .A(n96227), .ZN(
        \DLX_Datapath/RegisterFile/N25134 ) );
  AOI22_X1 U83423 ( .A1(n105999), .A2(n108650), .B1(n105997), .B2(n81417), 
        .ZN(n96227) );
  OAI21_X1 U83424 ( .B1(n106053), .B2(n106001), .A(n96228), .ZN(
        \DLX_Datapath/RegisterFile/N25133 ) );
  AOI22_X1 U83425 ( .A1(n106000), .A2(n108877), .B1(n105996), .B2(n81500), 
        .ZN(n96228) );
  OAI21_X1 U83426 ( .B1(n105219), .B2(n106001), .A(n96229), .ZN(
        \DLX_Datapath/RegisterFile/N25132 ) );
  AOI22_X1 U83427 ( .A1(n106000), .A2(n108765), .B1(n105997), .B2(n81335), 
        .ZN(n96229) );
  OAI21_X1 U83428 ( .B1(n106269), .B2(n106001), .A(n96230), .ZN(
        \DLX_Datapath/RegisterFile/N25131 ) );
  AOI22_X1 U83429 ( .A1(n105999), .A2(n107305), .B1(n105997), .B2(n81327), 
        .ZN(n96230) );
  NOR2_X1 U83432 ( .A1(n81619), .A2(n105094), .ZN(n96231) );
  AOI21_X1 U83433 ( .B1(n105199), .B2(n96166), .A(n94663), .ZN(n96204) );
  OR2_X1 U83434 ( .A1(n96013), .A2(n95131), .ZN(n96166) );
  NAND2_X1 U83435 ( .A1(n105131), .A2(n95132), .ZN(n81619) );
  OAI21_X1 U83436 ( .B1(n106146), .B2(n105429), .A(n96233), .ZN(
        \DLX_Datapath/RegisterFile/N25130 ) );
  AOI22_X1 U83437 ( .A1(n96234), .A2(n70314), .B1(n105428), .B2(n94667), .ZN(
        n96233) );
  OAI21_X1 U83438 ( .B1(n105971), .B2(n105429), .A(n96236), .ZN(
        \DLX_Datapath/RegisterFile/N25129 ) );
  AOI22_X1 U83439 ( .A1(n104924), .A2(n70456), .B1(n105427), .B2(n94670), .ZN(
        n96236) );
  OAI21_X1 U83440 ( .B1(n106136), .B2(n105429), .A(n96237), .ZN(
        \DLX_Datapath/RegisterFile/N25128 ) );
  AOI22_X1 U83441 ( .A1(n96234), .A2(n69509), .B1(n105428), .B2(n94672), .ZN(
        n96237) );
  OAI21_X1 U83442 ( .B1(n106210), .B2(n105429), .A(n96238), .ZN(
        \DLX_Datapath/RegisterFile/N25127 ) );
  AOI22_X1 U83443 ( .A1(n104925), .A2(n70170), .B1(n105427), .B2(n94674), .ZN(
        n96238) );
  OAI21_X1 U83444 ( .B1(n106204), .B2(n105429), .A(n96239), .ZN(
        \DLX_Datapath/RegisterFile/N25126 ) );
  AOI22_X1 U83445 ( .A1(n96234), .A2(n74016), .B1(n105428), .B2(n94676), .ZN(
        n96239) );
  OAI21_X1 U83446 ( .B1(n106099), .B2(n105429), .A(n96240), .ZN(
        \DLX_Datapath/RegisterFile/N25125 ) );
  AOI22_X1 U83447 ( .A1(n104924), .A2(n70603), .B1(n105427), .B2(n94678), .ZN(
        n96240) );
  OAI21_X1 U83448 ( .B1(n81270), .B2(n105429), .A(n96241), .ZN(
        \DLX_Datapath/RegisterFile/N25124 ) );
  AOI22_X1 U83449 ( .A1(n104924), .A2(n74157), .B1(n105428), .B2(n94680), .ZN(
        n96241) );
  OAI21_X1 U83450 ( .B1(n105992), .B2(n105429), .A(n96242), .ZN(
        \DLX_Datapath/RegisterFile/N25123 ) );
  AOI22_X1 U83451 ( .A1(n104925), .A2(n74297), .B1(n105427), .B2(n94682), .ZN(
        n96242) );
  OAI21_X1 U83452 ( .B1(n80190), .B2(n105429), .A(n96243), .ZN(
        \DLX_Datapath/RegisterFile/N25122 ) );
  AOI22_X1 U83453 ( .A1(n104924), .A2(n73733), .B1(n105427), .B2(n94684), .ZN(
        n96243) );
  OAI21_X1 U83454 ( .B1(n106190), .B2(n105429), .A(n96244), .ZN(
        \DLX_Datapath/RegisterFile/N25121 ) );
  AOI22_X1 U83455 ( .A1(n104924), .A2(n73437), .B1(n105426), .B2(n94686), .ZN(
        n96244) );
  OAI21_X1 U83456 ( .B1(n81383), .B2(n105429), .A(n96245), .ZN(
        \DLX_Datapath/RegisterFile/N25120 ) );
  AOI22_X1 U83457 ( .A1(n104924), .A2(n73874), .B1(n105426), .B2(n94688), .ZN(
        n96245) );
  OAI21_X1 U83458 ( .B1(n106185), .B2(n105429), .A(n96246), .ZN(
        \DLX_Datapath/RegisterFile/N25119 ) );
  AOI22_X1 U83459 ( .A1(n104925), .A2(n73586), .B1(n105426), .B2(n94690), .ZN(
        n96246) );
  OAI21_X1 U83460 ( .B1(n81345), .B2(n105429), .A(n96247), .ZN(
        \DLX_Datapath/RegisterFile/N25118 ) );
  AOI22_X1 U83461 ( .A1(n104925), .A2(n73148), .B1(n105426), .B2(n94692), .ZN(
        n96247) );
  OAI21_X1 U83462 ( .B1(n106105), .B2(n105429), .A(n96248), .ZN(
        \DLX_Datapath/RegisterFile/N25117 ) );
  AOI22_X1 U83463 ( .A1(n104925), .A2(n73290), .B1(n105426), .B2(n94694), .ZN(
        n96248) );
  OAI21_X1 U83464 ( .B1(n81294), .B2(n105429), .A(n96249), .ZN(
        \DLX_Datapath/RegisterFile/N25116 ) );
  AOI22_X1 U83465 ( .A1(n104924), .A2(n73006), .B1(n105426), .B2(n94696), .ZN(
        n96249) );
  OAI21_X1 U83466 ( .B1(n106108), .B2(n105429), .A(n96250), .ZN(
        \DLX_Datapath/RegisterFile/N25115 ) );
  AOI22_X1 U83467 ( .A1(n104924), .A2(n72856), .B1(n105426), .B2(n94698), .ZN(
        n96250) );
  OAI21_X1 U83468 ( .B1(n81284), .B2(n105429), .A(n96251), .ZN(
        \DLX_Datapath/RegisterFile/N25114 ) );
  AOI22_X1 U83469 ( .A1(n104925), .A2(n70752), .B1(n105426), .B2(n94700), .ZN(
        n96251) );
  OAI21_X1 U83470 ( .B1(n106172), .B2(n105429), .A(n96252), .ZN(
        \DLX_Datapath/RegisterFile/N25113 ) );
  AOI22_X1 U83471 ( .A1(n104924), .A2(n70911), .B1(n105426), .B2(n94702), .ZN(
        n96252) );
  OAI21_X1 U83472 ( .B1(n106236), .B2(n105429), .A(n96253), .ZN(
        \DLX_Datapath/RegisterFile/N25112 ) );
  AOI22_X1 U83473 ( .A1(n104924), .A2(n71056), .B1(n105426), .B2(n94704), .ZN(
        n96253) );
  OAI21_X1 U83474 ( .B1(n106072), .B2(n105429), .A(n96254), .ZN(
        \DLX_Datapath/RegisterFile/N25111 ) );
  AOI22_X1 U83475 ( .A1(n104924), .A2(n70017), .B1(n105426), .B2(n94706), .ZN(
        n96254) );
  OAI21_X1 U83476 ( .B1(n106197), .B2(n105429), .A(n96255), .ZN(
        \DLX_Datapath/RegisterFile/N25110 ) );
  AOI22_X1 U83477 ( .A1(n104925), .A2(n72546), .B1(n105427), .B2(n94708), .ZN(
        n96255) );
  OAI21_X1 U83478 ( .B1(n106243), .B2(n105429), .A(n96256), .ZN(
        \DLX_Datapath/RegisterFile/N25109 ) );
  AOI22_X1 U83479 ( .A1(n104925), .A2(n71205), .B1(n105428), .B2(n94710), .ZN(
        n96256) );
  OAI21_X1 U83480 ( .B1(n106157), .B2(n105429), .A(n96257), .ZN(
        \DLX_Datapath/RegisterFile/N25108 ) );
  AOI22_X1 U83481 ( .A1(n104925), .A2(n72688), .B1(n105427), .B2(n94712), .ZN(
        n96257) );
  OAI21_X1 U83482 ( .B1(n106116), .B2(n105429), .A(n96258), .ZN(
        \DLX_Datapath/RegisterFile/N25107 ) );
  AOI22_X1 U83483 ( .A1(n96234), .A2(n72398), .B1(n105428), .B2(n94714), .ZN(
        n96258) );
  OAI21_X1 U83484 ( .B1(n106009), .B2(n105429), .A(n96259), .ZN(
        \DLX_Datapath/RegisterFile/N25106 ) );
  AOI22_X1 U83485 ( .A1(n96234), .A2(n71798), .B1(n105427), .B2(n81259), .ZN(
        n96259) );
  OAI21_X1 U83486 ( .B1(n106260), .B2(n105429), .A(n96260), .ZN(
        \DLX_Datapath/RegisterFile/N25105 ) );
  AOI22_X1 U83487 ( .A1(n104924), .A2(n72247), .B1(n105428), .B2(n94717), .ZN(
        n96260) );
  OAI21_X1 U83488 ( .B1(n106043), .B2(n105429), .A(n96261), .ZN(
        \DLX_Datapath/RegisterFile/N25104 ) );
  AOI22_X1 U83489 ( .A1(n104925), .A2(n72096), .B1(n105427), .B2(n94719), .ZN(
        n96261) );
  OAI21_X1 U83490 ( .B1(n106049), .B2(n105429), .A(n96262), .ZN(
        \DLX_Datapath/RegisterFile/N25103 ) );
  AOI22_X1 U83491 ( .A1(n104924), .A2(n71952), .B1(n105428), .B2(n94721), .ZN(
        n96262) );
  OAI21_X1 U83492 ( .B1(n106094), .B2(n105429), .A(n96263), .ZN(
        \DLX_Datapath/RegisterFile/N25102 ) );
  AOI22_X1 U83493 ( .A1(n96234), .A2(n71354), .B1(n105427), .B2(n94723), .ZN(
        n96263) );
  OAI21_X1 U83494 ( .B1(n106053), .B2(n105429), .A(n96264), .ZN(
        \DLX_Datapath/RegisterFile/N25101 ) );
  AOI22_X1 U83495 ( .A1(n104924), .A2(n71649), .B1(n105428), .B2(n94725), .ZN(
        n96264) );
  OAI21_X1 U83496 ( .B1(n105219), .B2(n105429), .A(n96265), .ZN(
        \DLX_Datapath/RegisterFile/N25100 ) );
  AOI22_X1 U83497 ( .A1(n96234), .A2(n71505), .B1(n105428), .B2(n94727), .ZN(
        n96265) );
  OAI21_X1 U83498 ( .B1(n106267), .B2(n105429), .A(n96266), .ZN(
        \DLX_Datapath/RegisterFile/N25099 ) );
  AOI22_X1 U83499 ( .A1(n104925), .A2(n69614), .B1(n105427), .B2(n94729), .ZN(
        n96266) );
  OR2_X1 U83501 ( .A1(n96268), .A2(n95131), .ZN(n96267) );
  AOI21_X1 U83502 ( .B1(n96269), .B2(n105602), .A(n96268), .ZN(n96234) );
  NOR2_X1 U83503 ( .A1(n96232), .A2(n105091), .ZN(n96268) );
  OAI21_X1 U83504 ( .B1(n106757), .B2(n95131), .A(n105199), .ZN(n96269) );
  NAND2_X1 U83505 ( .A1(n105132), .A2(n94505), .ZN(n96232) );
  OAI21_X1 U83506 ( .B1(n105971), .B2(n105936), .A(n96270), .ZN(
        \DLX_Datapath/RegisterFile/N25097 ) );
  AOI22_X1 U83507 ( .A1(n105934), .A2(n107969), .B1(n94511), .B2(n105931), 
        .ZN(n96270) );
  OAI21_X1 U83508 ( .B1(n106204), .B2(n105936), .A(n96271), .ZN(
        \DLX_Datapath/RegisterFile/N25094 ) );
  AOI22_X1 U83509 ( .A1(n105934), .A2(n110673), .B1(n105930), .B2(n81308), 
        .ZN(n96271) );
  OAI21_X1 U83510 ( .B1(n106100), .B2(n105936), .A(n96272), .ZN(
        \DLX_Datapath/RegisterFile/N25093 ) );
  AOI22_X1 U83511 ( .A1(n105934), .A2(n108072), .B1(n94516), .B2(n105931), 
        .ZN(n96272) );
  OAI21_X1 U83512 ( .B1(n81270), .B2(n105936), .A(n96273), .ZN(
        \DLX_Datapath/RegisterFile/N25092 ) );
  AOI22_X1 U83513 ( .A1(n105934), .A2(n110770), .B1(n105932), .B2(n81272), 
        .ZN(n96273) );
  OAI21_X1 U83514 ( .B1(n105992), .B2(n105936), .A(n96274), .ZN(
        \DLX_Datapath/RegisterFile/N25091 ) );
  AOI22_X1 U83515 ( .A1(n105934), .A2(n110871), .B1(n94519), .B2(n105931), 
        .ZN(n96274) );
  OAI21_X1 U83516 ( .B1(n106333), .B2(n105936), .A(n96275), .ZN(
        \DLX_Datapath/RegisterFile/N25090 ) );
  AOI22_X1 U83517 ( .A1(n105934), .A2(n110466), .B1(n105932), .B2(n80192), 
        .ZN(n96275) );
  OAI21_X1 U83518 ( .B1(n106190), .B2(n105936), .A(n96276), .ZN(
        \DLX_Datapath/RegisterFile/N25089 ) );
  AOI22_X1 U83519 ( .A1(n105934), .A2(n110248), .B1(n105930), .B2(n81474), 
        .ZN(n96276) );
  OAI21_X1 U83520 ( .B1(n81383), .B2(n105936), .A(n96277), .ZN(
        \DLX_Datapath/RegisterFile/N25088 ) );
  AOI22_X1 U83521 ( .A1(n105934), .A2(n110565), .B1(n94523), .B2(n105931), 
        .ZN(n96277) );
  OAI21_X1 U83522 ( .B1(n106185), .B2(n105936), .A(n96278), .ZN(
        \DLX_Datapath/RegisterFile/N25087 ) );
  AOI22_X1 U83523 ( .A1(n105934), .A2(n110356), .B1(n105932), .B2(n106061), 
        .ZN(n96278) );
  OAI21_X1 U83524 ( .B1(n81345), .B2(n105936), .A(n96279), .ZN(
        \DLX_Datapath/RegisterFile/N25086 ) );
  AOI22_X1 U83525 ( .A1(n105934), .A2(n110031), .B1(n105930), .B2(n81347), 
        .ZN(n96279) );
  OAI21_X1 U83526 ( .B1(n106103), .B2(n105936), .A(n96280), .ZN(
        \DLX_Datapath/RegisterFile/N25085 ) );
  AOI22_X1 U83527 ( .A1(n105934), .A2(n110138), .B1(n94527), .B2(n105931), 
        .ZN(n96280) );
  OAI21_X1 U83528 ( .B1(n81294), .B2(n105936), .A(n96281), .ZN(
        \DLX_Datapath/RegisterFile/N25084 ) );
  AOI22_X1 U83529 ( .A1(n105933), .A2(n109922), .B1(n105932), .B2(n81297), 
        .ZN(n96281) );
  OAI21_X1 U83530 ( .B1(n81398), .B2(n105936), .A(n96282), .ZN(
        \DLX_Datapath/RegisterFile/N25083 ) );
  AOI22_X1 U83531 ( .A1(n105933), .A2(n109804), .B1(n94530), .B2(n105931), 
        .ZN(n96282) );
  OAI21_X1 U83532 ( .B1(n106172), .B2(n105936), .A(n96283), .ZN(
        \DLX_Datapath/RegisterFile/N25081 ) );
  AOI22_X1 U83533 ( .A1(n105935), .A2(n108301), .B1(n105930), .B2(n106168), 
        .ZN(n96283) );
  OAI21_X1 U83534 ( .B1(n106072), .B2(n81733), .A(n96284), .ZN(
        \DLX_Datapath/RegisterFile/N25079 ) );
  AOI22_X1 U83535 ( .A1(n105933), .A2(n107650), .B1(n105932), .B2(n81453), 
        .ZN(n96284) );
  OAI21_X1 U83536 ( .B1(n106197), .B2(n81733), .A(n96285), .ZN(
        \DLX_Datapath/RegisterFile/N25078 ) );
  AOI22_X1 U83537 ( .A1(n105935), .A2(n109568), .B1(n94536), .B2(n105931), 
        .ZN(n96285) );
  OAI21_X1 U83538 ( .B1(n106157), .B2(n81733), .A(n96286), .ZN(
        \DLX_Datapath/RegisterFile/N25076 ) );
  AOI22_X1 U83539 ( .A1(n105933), .A2(n109673), .B1(n105930), .B2(n81351), 
        .ZN(n96286) );
  OAI21_X1 U83540 ( .B1(n106008), .B2(n81733), .A(n96287), .ZN(
        \DLX_Datapath/RegisterFile/N25074 ) );
  AOI22_X1 U83541 ( .A1(n105935), .A2(n108994), .B1(n94541), .B2(n105931), 
        .ZN(n96287) );
  OAI21_X1 U83542 ( .B1(n81509), .B2(n105936), .A(n96288), .ZN(
        \DLX_Datapath/RegisterFile/N25072 ) );
  AOI22_X1 U83543 ( .A1(n105933), .A2(n109224), .B1(n105624), .B2(n105930), 
        .ZN(n96288) );
  OAI21_X1 U83544 ( .B1(n106049), .B2(n81733), .A(n96289), .ZN(
        \DLX_Datapath/RegisterFile/N25071 ) );
  AOI22_X1 U83545 ( .A1(n105935), .A2(n109116), .B1(n94546), .B2(n105931), 
        .ZN(n96289) );
  OAI21_X1 U83546 ( .B1(n106095), .B2(n81733), .A(n96290), .ZN(
        \DLX_Datapath/RegisterFile/N25070 ) );
  AOI22_X1 U83547 ( .A1(n105933), .A2(n108651), .B1(n94548), .B2(n105931), 
        .ZN(n96290) );
  OAI21_X1 U83548 ( .B1(n106053), .B2(n81733), .A(n96291), .ZN(
        \DLX_Datapath/RegisterFile/N25069 ) );
  AOI22_X1 U83549 ( .A1(n105935), .A2(n108878), .B1(n81783), .B2(n105932), 
        .ZN(n96291) );
  OAI21_X1 U83550 ( .B1(n106267), .B2(n81733), .A(n96292), .ZN(
        \DLX_Datapath/RegisterFile/N25067 ) );
  AOI22_X1 U83551 ( .A1(n105933), .A2(n107306), .B1(n105930), .B2(n81265), 
        .ZN(n96292) );
  AOI21_X1 U83553 ( .B1(n96010), .B2(n94554), .A(n96294), .ZN(n81735) );
  NOR2_X1 U83554 ( .A1(n81733), .A2(n105090), .ZN(n96294) );
  NAND2_X1 U83555 ( .A1(n105131), .A2(n94555), .ZN(n81733) );
  OAI21_X1 U83556 ( .B1(n81358), .B2(n105425), .A(n96296), .ZN(
        \DLX_Datapath/RegisterFile/N25066 ) );
  AOI22_X1 U83557 ( .A1(n105424), .A2(n70316), .B1(n104959), .B2(n94559), .ZN(
        n96296) );
  OAI21_X1 U83558 ( .B1(n105970), .B2(n105425), .A(n96299), .ZN(
        \DLX_Datapath/RegisterFile/N25065 ) );
  AOI22_X1 U83559 ( .A1(n105423), .A2(n70458), .B1(n104960), .B2(n94562), .ZN(
        n96299) );
  OAI21_X1 U83560 ( .B1(n106136), .B2(n105425), .A(n96300), .ZN(
        \DLX_Datapath/RegisterFile/N25064 ) );
  AOI22_X1 U83561 ( .A1(n105424), .A2(n69511), .B1(n104959), .B2(n94564), .ZN(
        n96300) );
  OAI21_X1 U83562 ( .B1(n106211), .B2(n105425), .A(n96301), .ZN(
        \DLX_Datapath/RegisterFile/N25063 ) );
  AOI22_X1 U83563 ( .A1(n105423), .A2(n70172), .B1(n104961), .B2(n94566), .ZN(
        n96301) );
  OAI21_X1 U83564 ( .B1(n106204), .B2(n105425), .A(n96302), .ZN(
        \DLX_Datapath/RegisterFile/N25062 ) );
  AOI22_X1 U83565 ( .A1(n105424), .A2(n74018), .B1(n104959), .B2(n94568), .ZN(
        n96302) );
  OAI21_X1 U83566 ( .B1(n106098), .B2(n105425), .A(n96303), .ZN(
        \DLX_Datapath/RegisterFile/N25061 ) );
  AOI22_X1 U83567 ( .A1(n105423), .A2(n70605), .B1(n104960), .B2(n94570), .ZN(
        n96303) );
  OAI21_X1 U83568 ( .B1(n81270), .B2(n105425), .A(n96304), .ZN(
        \DLX_Datapath/RegisterFile/N25060 ) );
  AOI22_X1 U83569 ( .A1(n105424), .A2(n74159), .B1(n104960), .B2(n94572), .ZN(
        n96304) );
  OAI21_X1 U83570 ( .B1(n105992), .B2(n105425), .A(n96305), .ZN(
        \DLX_Datapath/RegisterFile/N25059 ) );
  AOI22_X1 U83571 ( .A1(n105423), .A2(n74299), .B1(n104961), .B2(n94574), .ZN(
        n96305) );
  OAI21_X1 U83572 ( .B1(n80190), .B2(n105425), .A(n96306), .ZN(
        \DLX_Datapath/RegisterFile/N25058 ) );
  AOI22_X1 U83573 ( .A1(n105423), .A2(n73735), .B1(n104960), .B2(n94576), .ZN(
        n96306) );
  OAI21_X1 U83574 ( .B1(n106190), .B2(n105425), .A(n96307), .ZN(
        \DLX_Datapath/RegisterFile/N25057 ) );
  AOI22_X1 U83575 ( .A1(n105422), .A2(n73439), .B1(n104959), .B2(n94578), .ZN(
        n96307) );
  OAI21_X1 U83576 ( .B1(n81383), .B2(n105425), .A(n96308), .ZN(
        \DLX_Datapath/RegisterFile/N25056 ) );
  AOI22_X1 U83577 ( .A1(n105422), .A2(n73876), .B1(n104960), .B2(n94580), .ZN(
        n96308) );
  OAI21_X1 U83578 ( .B1(n106185), .B2(n105425), .A(n96309), .ZN(
        \DLX_Datapath/RegisterFile/N25055 ) );
  AOI22_X1 U83579 ( .A1(n105422), .A2(n73588), .B1(n104961), .B2(n94582), .ZN(
        n96309) );
  OAI21_X1 U83580 ( .B1(n81345), .B2(n105425), .A(n96310), .ZN(
        \DLX_Datapath/RegisterFile/N25054 ) );
  AOI22_X1 U83581 ( .A1(n105422), .A2(n73150), .B1(n104961), .B2(n94584), .ZN(
        n96310) );
  OAI21_X1 U83582 ( .B1(n106103), .B2(n105425), .A(n96311), .ZN(
        \DLX_Datapath/RegisterFile/N25053 ) );
  AOI22_X1 U83583 ( .A1(n105422), .A2(n73292), .B1(n104959), .B2(n94586), .ZN(
        n96311) );
  OAI21_X1 U83584 ( .B1(n106221), .B2(n105425), .A(n96312), .ZN(
        \DLX_Datapath/RegisterFile/N25052 ) );
  AOI22_X1 U83585 ( .A1(n105422), .A2(n73008), .B1(n104959), .B2(n94588), .ZN(
        n96312) );
  OAI21_X1 U83586 ( .B1(n106109), .B2(n105425), .A(n96313), .ZN(
        \DLX_Datapath/RegisterFile/N25051 ) );
  AOI22_X1 U83587 ( .A1(n105422), .A2(n72858), .B1(n104960), .B2(n94590), .ZN(
        n96313) );
  OAI21_X1 U83588 ( .B1(n81284), .B2(n105425), .A(n96314), .ZN(
        \DLX_Datapath/RegisterFile/N25050 ) );
  AOI22_X1 U83589 ( .A1(n105422), .A2(n70754), .B1(n104961), .B2(n94592), .ZN(
        n96314) );
  OAI21_X1 U83590 ( .B1(n106170), .B2(n105425), .A(n96315), .ZN(
        \DLX_Datapath/RegisterFile/N25049 ) );
  AOI22_X1 U83591 ( .A1(n105422), .A2(n70913), .B1(n104960), .B2(n94594), .ZN(
        n96315) );
  OAI21_X1 U83592 ( .B1(n106236), .B2(n105425), .A(n96316), .ZN(
        \DLX_Datapath/RegisterFile/N25048 ) );
  AOI22_X1 U83593 ( .A1(n105422), .A2(n71058), .B1(n104959), .B2(n94596), .ZN(
        n96316) );
  OAI21_X1 U83594 ( .B1(n106072), .B2(n105425), .A(n96317), .ZN(
        \DLX_Datapath/RegisterFile/N25047 ) );
  AOI22_X1 U83595 ( .A1(n105422), .A2(n70019), .B1(n104960), .B2(n94598), .ZN(
        n96317) );
  OAI21_X1 U83596 ( .B1(n106197), .B2(n105425), .A(n96318), .ZN(
        \DLX_Datapath/RegisterFile/N25046 ) );
  AOI22_X1 U83597 ( .A1(n105423), .A2(n72548), .B1(n104961), .B2(n94600), .ZN(
        n96318) );
  OAI21_X1 U83598 ( .B1(n81278), .B2(n105425), .A(n96319), .ZN(
        \DLX_Datapath/RegisterFile/N25045 ) );
  AOI22_X1 U83599 ( .A1(n105424), .A2(n71207), .B1(n104961), .B2(n94602), .ZN(
        n96319) );
  OAI21_X1 U83600 ( .B1(n106157), .B2(n96295), .A(n96320), .ZN(
        \DLX_Datapath/RegisterFile/N25044 ) );
  AOI22_X1 U83601 ( .A1(n105423), .A2(n72690), .B1(n104961), .B2(n94604), .ZN(
        n96320) );
  OAI21_X1 U83602 ( .B1(n106113), .B2(n96295), .A(n96321), .ZN(
        \DLX_Datapath/RegisterFile/N25043 ) );
  AOI22_X1 U83603 ( .A1(n105424), .A2(n72400), .B1(n104959), .B2(n94606), .ZN(
        n96321) );
  OAI21_X1 U83604 ( .B1(n106008), .B2(n96295), .A(n96322), .ZN(
        \DLX_Datapath/RegisterFile/N25042 ) );
  AOI22_X1 U83605 ( .A1(n105423), .A2(n71800), .B1(n104959), .B2(n94608), .ZN(
        n96322) );
  OAI21_X1 U83606 ( .B1(n106261), .B2(n96295), .A(n96323), .ZN(
        \DLX_Datapath/RegisterFile/N25041 ) );
  AOI22_X1 U83607 ( .A1(n105424), .A2(n72249), .B1(n104960), .B2(n94610), .ZN(
        n96323) );
  OAI21_X1 U83608 ( .B1(n81509), .B2(n105425), .A(n96324), .ZN(
        \DLX_Datapath/RegisterFile/N25040 ) );
  AOI22_X1 U83609 ( .A1(n105423), .A2(n72098), .B1(n104961), .B2(n94612), .ZN(
        n96324) );
  OAI21_X1 U83610 ( .B1(n106049), .B2(n96295), .A(n96325), .ZN(
        \DLX_Datapath/RegisterFile/N25039 ) );
  AOI22_X1 U83611 ( .A1(n105424), .A2(n71954), .B1(n104960), .B2(n94614), .ZN(
        n96325) );
  OAI21_X1 U83612 ( .B1(n106093), .B2(n96295), .A(n96326), .ZN(
        \DLX_Datapath/RegisterFile/N25038 ) );
  AOI22_X1 U83613 ( .A1(n105423), .A2(n71356), .B1(n104959), .B2(n94616), .ZN(
        n96326) );
  OAI21_X1 U83614 ( .B1(n106053), .B2(n96295), .A(n96327), .ZN(
        \DLX_Datapath/RegisterFile/N25037 ) );
  AOI22_X1 U83615 ( .A1(n105424), .A2(n71651), .B1(n104960), .B2(n94618), .ZN(
        n96327) );
  OAI21_X1 U83616 ( .B1(n105219), .B2(n96295), .A(n96328), .ZN(
        \DLX_Datapath/RegisterFile/N25036 ) );
  AOI22_X1 U83617 ( .A1(n105424), .A2(n71507), .B1(n104959), .B2(n94620), .ZN(
        n96328) );
  OAI21_X1 U83618 ( .B1(n106267), .B2(n96295), .A(n96329), .ZN(
        \DLX_Datapath/RegisterFile/N25035 ) );
  AOI22_X1 U83619 ( .A1(n105423), .A2(n69616), .B1(n104961), .B2(n94622), .ZN(
        n96329) );
  NOR2_X1 U83622 ( .A1(n96295), .A2(n105094), .ZN(n96330) );
  NAND2_X1 U83623 ( .A1(n94625), .A2(n105132), .ZN(n96295) );
  OAI21_X1 U83624 ( .B1(n81634), .B2(n81651), .A(n96332), .ZN(
        \DLX_Datapath/RegisterFile/N25033 ) );
  AOI22_X1 U83625 ( .A1(n105981), .A2(n107970), .B1(n81653), .B2(n105977), 
        .ZN(n96332) );
  OAI21_X1 U83626 ( .B1(n106204), .B2(n105983), .A(n96333), .ZN(
        \DLX_Datapath/RegisterFile/N25030 ) );
  AOI22_X1 U83627 ( .A1(n105980), .A2(n110674), .B1(n105977), .B2(n81428), 
        .ZN(n96333) );
  OAI21_X1 U83628 ( .B1(n106098), .B2(n105983), .A(n96334), .ZN(
        \DLX_Datapath/RegisterFile/N25029 ) );
  AOI22_X1 U83629 ( .A1(n105982), .A2(n108073), .B1(n105978), .B2(n81410), 
        .ZN(n96334) );
  OAI21_X1 U83630 ( .B1(n81270), .B2(n105983), .A(n96335), .ZN(
        \DLX_Datapath/RegisterFile/N25028 ) );
  AOI22_X1 U83631 ( .A1(n105981), .A2(n110771), .B1(n81700), .B2(n105977), 
        .ZN(n96335) );
  OAI21_X1 U83632 ( .B1(n105991), .B2(n105983), .A(n96336), .ZN(
        \DLX_Datapath/RegisterFile/N25027 ) );
  AOI22_X1 U83633 ( .A1(n105982), .A2(n110872), .B1(n105979), .B2(n81632), 
        .ZN(n96336) );
  OAI21_X1 U83634 ( .B1(n80190), .B2(n105983), .A(n96337), .ZN(
        \DLX_Datapath/RegisterFile/N25026 ) );
  AOI22_X1 U83635 ( .A1(n105980), .A2(n110467), .B1(n105978), .B2(n81414), 
        .ZN(n96337) );
  OAI21_X1 U83636 ( .B1(n106190), .B2(n105983), .A(n96338), .ZN(
        \DLX_Datapath/RegisterFile/N25025 ) );
  AOI22_X1 U83637 ( .A1(n105980), .A2(n110249), .B1(n105977), .B2(n81317), 
        .ZN(n96338) );
  OAI21_X1 U83638 ( .B1(n81383), .B2(n105983), .A(n96339), .ZN(
        \DLX_Datapath/RegisterFile/N25024 ) );
  AOI22_X1 U83639 ( .A1(n105980), .A2(n110566), .B1(n105977), .B2(n81386), 
        .ZN(n96339) );
  OAI21_X1 U83640 ( .B1(n106185), .B2(n105983), .A(n96340), .ZN(
        \DLX_Datapath/RegisterFile/N25023 ) );
  AOI22_X1 U83641 ( .A1(n105980), .A2(n110357), .B1(n105977), .B2(n81320), 
        .ZN(n96340) );
  OAI21_X1 U83642 ( .B1(n81345), .B2(n105983), .A(n96341), .ZN(
        \DLX_Datapath/RegisterFile/N25022 ) );
  AOI22_X1 U83643 ( .A1(n105980), .A2(n110032), .B1(n105977), .B2(n81604), 
        .ZN(n96341) );
  OAI21_X1 U83644 ( .B1(n106103), .B2(n105983), .A(n96342), .ZN(
        \DLX_Datapath/RegisterFile/N25021 ) );
  AOI22_X1 U83645 ( .A1(n105980), .A2(n110139), .B1(n105977), .B2(n81405), 
        .ZN(n96342) );
  OAI21_X1 U83646 ( .B1(n81294), .B2(n105983), .A(n96343), .ZN(
        \DLX_Datapath/RegisterFile/N25020 ) );
  AOI22_X1 U83647 ( .A1(n105980), .A2(n109923), .B1(n105977), .B2(n81402), 
        .ZN(n96343) );
  OAI21_X1 U83648 ( .B1(n106109), .B2(n105983), .A(n96344), .ZN(
        \DLX_Datapath/RegisterFile/N25019 ) );
  AOI22_X1 U83649 ( .A1(n105981), .A2(n109805), .B1(n105978), .B2(n81400), 
        .ZN(n96344) );
  OAI21_X1 U83650 ( .B1(n106072), .B2(n105983), .A(n96345), .ZN(
        \DLX_Datapath/RegisterFile/N25015 ) );
  AOI22_X1 U83651 ( .A1(n105981), .A2(n107651), .B1(n105978), .B2(n81506), 
        .ZN(n96345) );
  OAI21_X1 U83652 ( .B1(n106197), .B2(n105983), .A(n96346), .ZN(
        \DLX_Datapath/RegisterFile/N25014 ) );
  AOI22_X1 U83653 ( .A1(n105981), .A2(n109569), .B1(n105978), .B2(n81313), 
        .ZN(n96346) );
  OAI21_X1 U83654 ( .B1(n106157), .B2(n105983), .A(n96347), .ZN(
        \DLX_Datapath/RegisterFile/N25012 ) );
  AOI22_X1 U83655 ( .A1(n105982), .A2(n109674), .B1(n105979), .B2(n81425), 
        .ZN(n96347) );
  OAI21_X1 U83656 ( .B1(n106114), .B2(n105983), .A(n96348), .ZN(
        \DLX_Datapath/RegisterFile/N25011 ) );
  AOI22_X1 U83657 ( .A1(n105981), .A2(n109458), .B1(n105978), .B2(n81396), 
        .ZN(n96348) );
  OAI21_X1 U83658 ( .B1(n106008), .B2(n105983), .A(n96349), .ZN(
        \DLX_Datapath/RegisterFile/N25010 ) );
  AOI22_X1 U83659 ( .A1(n105982), .A2(n108995), .B1(n105979), .B2(n81590), 
        .ZN(n96349) );
  OAI21_X1 U83660 ( .B1(n106262), .B2(n105983), .A(n96350), .ZN(
        \DLX_Datapath/RegisterFile/N25009 ) );
  AOI22_X1 U83661 ( .A1(n105982), .A2(n109343), .B1(n105979), .B2(n81423), 
        .ZN(n96350) );
  OAI21_X1 U83662 ( .B1(n106044), .B2(n105983), .A(n96351), .ZN(
        \DLX_Datapath/RegisterFile/N25008 ) );
  AOI22_X1 U83663 ( .A1(n105981), .A2(n109225), .B1(n105978), .B2(n81511), 
        .ZN(n96351) );
  OAI21_X1 U83664 ( .B1(n106049), .B2(n105983), .A(n96352), .ZN(
        \DLX_Datapath/RegisterFile/N25007 ) );
  AOI22_X1 U83665 ( .A1(n105982), .A2(n109117), .B1(n105979), .B2(n81503), 
        .ZN(n96352) );
  OAI21_X1 U83666 ( .B1(n106267), .B2(n81634), .A(n96353), .ZN(
        \DLX_Datapath/RegisterFile/N25003 ) );
  AOI22_X1 U83667 ( .A1(n105982), .A2(n107307), .B1(n105979), .B2(n81327), 
        .ZN(n96353) );
  NOR2_X1 U83670 ( .A1(n81634), .A2(n105090), .ZN(n96354) );
  AOI21_X1 U83671 ( .B1(n105199), .B2(n96293), .A(n105601), .ZN(n96331) );
  OR2_X1 U83672 ( .A1(n96013), .A2(n86230), .ZN(n96293) );
  NAND2_X1 U83673 ( .A1(n105132), .A2(n94664), .ZN(n81634) );
  OAI21_X1 U83674 ( .B1(n81358), .B2(n105420), .A(n96356), .ZN(
        \DLX_Datapath/RegisterFile/N25002 ) );
  AOI22_X1 U83675 ( .A1(n104836), .A2(n94667), .B1(n105419), .B2(n107873), 
        .ZN(n96356) );
  OAI21_X1 U83676 ( .B1(n105971), .B2(n105421), .A(n96359), .ZN(
        \DLX_Datapath/RegisterFile/N25001 ) );
  AOI22_X1 U83677 ( .A1(n104836), .A2(n94670), .B1(n105418), .B2(n107971), 
        .ZN(n96359) );
  OAI21_X1 U83678 ( .B1(n106136), .B2(n105420), .A(n96360), .ZN(
        \DLX_Datapath/RegisterFile/N25000 ) );
  AOI22_X1 U83679 ( .A1(n104836), .A2(n94672), .B1(n96358), .B2(n107234), .ZN(
        n96360) );
  OAI21_X1 U83680 ( .B1(n106210), .B2(n105421), .A(n96361), .ZN(
        \DLX_Datapath/RegisterFile/N24999 ) );
  AOI22_X1 U83681 ( .A1(n104836), .A2(n94674), .B1(n96358), .B2(n107772), .ZN(
        n96361) );
  OAI21_X1 U83682 ( .B1(n106204), .B2(n105420), .A(n96362), .ZN(
        \DLX_Datapath/RegisterFile/N24998 ) );
  AOI22_X1 U83683 ( .A1(n104837), .A2(n94676), .B1(n96358), .B2(n110675), .ZN(
        n96362) );
  OAI21_X1 U83684 ( .B1(n106098), .B2(n105420), .A(n96363), .ZN(
        \DLX_Datapath/RegisterFile/N24997 ) );
  AOI22_X1 U83685 ( .A1(n104838), .A2(n94678), .B1(n96358), .B2(n108074), .ZN(
        n96363) );
  OAI21_X1 U83686 ( .B1(n106254), .B2(n105421), .A(n96364), .ZN(
        \DLX_Datapath/RegisterFile/N24996 ) );
  AOI22_X1 U83687 ( .A1(n104837), .A2(n94680), .B1(n96358), .B2(n110772), .ZN(
        n96364) );
  OAI21_X1 U83688 ( .B1(n105990), .B2(n105420), .A(n96365), .ZN(
        \DLX_Datapath/RegisterFile/N24995 ) );
  AOI22_X1 U83689 ( .A1(n104838), .A2(n94682), .B1(n96358), .B2(n110873), .ZN(
        n96365) );
  OAI21_X1 U83690 ( .B1(n106333), .B2(n105420), .A(n96366), .ZN(
        \DLX_Datapath/RegisterFile/N24994 ) );
  AOI22_X1 U83691 ( .A1(n104838), .A2(n94684), .B1(n105419), .B2(n110468), 
        .ZN(n96366) );
  OAI21_X1 U83692 ( .B1(n106190), .B2(n105421), .A(n96367), .ZN(
        \DLX_Datapath/RegisterFile/N24993 ) );
  AOI22_X1 U83693 ( .A1(n104837), .A2(n94686), .B1(n105419), .B2(n110250), 
        .ZN(n96367) );
  AOI22_X1 U83695 ( .A1(n104836), .A2(n94688), .B1(n105419), .B2(n110567), 
        .ZN(n96368) );
  OAI21_X1 U83696 ( .B1(n106185), .B2(n105420), .A(n96369), .ZN(
        \DLX_Datapath/RegisterFile/N24991 ) );
  AOI22_X1 U83697 ( .A1(n104838), .A2(n94690), .B1(n105419), .B2(n110358), 
        .ZN(n96369) );
  OAI21_X1 U83698 ( .B1(n81345), .B2(n105420), .A(n96370), .ZN(
        \DLX_Datapath/RegisterFile/N24990 ) );
  AOI22_X1 U83699 ( .A1(n104836), .A2(n94692), .B1(n105419), .B2(n110033), 
        .ZN(n96370) );
  OAI21_X1 U83700 ( .B1(n106103), .B2(n105420), .A(n96371), .ZN(
        \DLX_Datapath/RegisterFile/N24989 ) );
  AOI22_X1 U83701 ( .A1(n104837), .A2(n94694), .B1(n105419), .B2(n110140), 
        .ZN(n96371) );
  OAI21_X1 U83702 ( .B1(n106218), .B2(n105421), .A(n96372), .ZN(
        \DLX_Datapath/RegisterFile/N24988 ) );
  AOI22_X1 U83703 ( .A1(n104838), .A2(n94696), .B1(n105419), .B2(n109924), 
        .ZN(n96372) );
  OAI21_X1 U83704 ( .B1(n81398), .B2(n105420), .A(n96373), .ZN(
        \DLX_Datapath/RegisterFile/N24987 ) );
  AOI22_X1 U83705 ( .A1(n104837), .A2(n94698), .B1(n105419), .B2(n109806), 
        .ZN(n96373) );
  OAI21_X1 U83706 ( .B1(n106233), .B2(n105420), .A(n96374), .ZN(
        \DLX_Datapath/RegisterFile/N24986 ) );
  AOI22_X1 U83707 ( .A1(n104838), .A2(n94700), .B1(n105419), .B2(n108180), 
        .ZN(n96374) );
  OAI21_X1 U83708 ( .B1(n106170), .B2(n105421), .A(n96375), .ZN(
        \DLX_Datapath/RegisterFile/N24985 ) );
  AOI22_X1 U83709 ( .A1(n104838), .A2(n94702), .B1(n105419), .B2(n108303), 
        .ZN(n96375) );
  OAI21_X1 U83710 ( .B1(n106236), .B2(n105420), .A(n96376), .ZN(
        \DLX_Datapath/RegisterFile/N24984 ) );
  AOI22_X1 U83711 ( .A1(n104836), .A2(n94704), .B1(n105419), .B2(n108414), 
        .ZN(n96376) );
  OAI21_X1 U83712 ( .B1(n106071), .B2(n105420), .A(n96377), .ZN(
        \DLX_Datapath/RegisterFile/N24983 ) );
  AOI22_X1 U83713 ( .A1(n104836), .A2(n94706), .B1(n105419), .B2(n107652), 
        .ZN(n96377) );
  OAI21_X1 U83714 ( .B1(n106197), .B2(n105421), .A(n96378), .ZN(
        \DLX_Datapath/RegisterFile/N24982 ) );
  AOI22_X1 U83715 ( .A1(n104836), .A2(n94708), .B1(n105418), .B2(n109570), 
        .ZN(n96378) );
  OAI21_X1 U83716 ( .B1(n106244), .B2(n105421), .A(n96379), .ZN(
        \DLX_Datapath/RegisterFile/N24981 ) );
  AOI22_X1 U83717 ( .A1(n104837), .A2(n94710), .B1(n105418), .B2(n108531), 
        .ZN(n96379) );
  OAI21_X1 U83718 ( .B1(n106157), .B2(n105420), .A(n96380), .ZN(
        \DLX_Datapath/RegisterFile/N24980 ) );
  AOI22_X1 U83719 ( .A1(n104838), .A2(n94712), .B1(n105418), .B2(n109675), 
        .ZN(n96380) );
  OAI21_X1 U83720 ( .B1(n106113), .B2(n105421), .A(n96381), .ZN(
        \DLX_Datapath/RegisterFile/N24979 ) );
  AOI22_X1 U83721 ( .A1(n104838), .A2(n94714), .B1(n105418), .B2(n109459), 
        .ZN(n96381) );
  OAI21_X1 U83722 ( .B1(n106008), .B2(n105421), .A(n96382), .ZN(
        \DLX_Datapath/RegisterFile/N24978 ) );
  AOI22_X1 U83723 ( .A1(n104836), .A2(n81259), .B1(n105418), .B2(n108996), 
        .ZN(n96382) );
  OAI21_X1 U83724 ( .B1(n106262), .B2(n105420), .A(n96383), .ZN(
        \DLX_Datapath/RegisterFile/N24977 ) );
  AOI22_X1 U83725 ( .A1(n104836), .A2(n94717), .B1(n105418), .B2(n109344), 
        .ZN(n96383) );
  OAI21_X1 U83726 ( .B1(n106045), .B2(n105420), .A(n96384), .ZN(
        \DLX_Datapath/RegisterFile/N24976 ) );
  AOI22_X1 U83727 ( .A1(n104836), .A2(n94719), .B1(n105418), .B2(n109226), 
        .ZN(n96384) );
  OAI21_X1 U83728 ( .B1(n106049), .B2(n105421), .A(n96385), .ZN(
        \DLX_Datapath/RegisterFile/N24975 ) );
  AOI22_X1 U83729 ( .A1(n104837), .A2(n94721), .B1(n105418), .B2(n109118), 
        .ZN(n96385) );
  OAI21_X1 U83730 ( .B1(n81415), .B2(n105420), .A(n96386), .ZN(
        \DLX_Datapath/RegisterFile/N24974 ) );
  AOI22_X1 U83731 ( .A1(n104838), .A2(n94723), .B1(n105418), .B2(n108653), 
        .ZN(n96386) );
  OAI21_X1 U83732 ( .B1(n106053), .B2(n105420), .A(n96387), .ZN(
        \DLX_Datapath/RegisterFile/N24973 ) );
  AOI22_X1 U83733 ( .A1(n104837), .A2(n94725), .B1(n105418), .B2(n108880), 
        .ZN(n96387) );
  OAI21_X1 U83734 ( .B1(n105219), .B2(n105421), .A(n96388), .ZN(
        \DLX_Datapath/RegisterFile/N24972 ) );
  AOI22_X1 U83735 ( .A1(n104837), .A2(n94727), .B1(n105418), .B2(n108768), 
        .ZN(n96388) );
  OAI21_X1 U83736 ( .B1(n106267), .B2(n105421), .A(n96389), .ZN(
        \DLX_Datapath/RegisterFile/N24971 ) );
  AOI22_X1 U83737 ( .A1(n104838), .A2(n94729), .B1(n105418), .B2(n107308), 
        .ZN(n96389) );
  AOI21_X1 U83738 ( .B1(n96390), .B2(n105602), .A(n96391), .ZN(n96358) );
  OAI21_X1 U83739 ( .B1(n106757), .B2(n86230), .A(n105206), .ZN(n96390) );
  NOR2_X1 U83740 ( .A1(n96392), .A2(n106757), .ZN(n96357) );
  OR2_X1 U83741 ( .A1(n96391), .A2(n86230), .ZN(n96392) );
  NOR2_X1 U83742 ( .A1(n96355), .A2(n105094), .ZN(n96391) );
  NAND2_X1 U83743 ( .A1(n94734), .A2(n105131), .ZN(n96355) );
  OAI21_X1 U83744 ( .B1(n105971), .B2(n105929), .A(n96393), .ZN(
        \DLX_Datapath/RegisterFile/N24969 ) );
  AOI22_X1 U83745 ( .A1(n70461), .A2(n105927), .B1(n94511), .B2(n105924), .ZN(
        n96393) );
  OAI21_X1 U83746 ( .B1(n106136), .B2(n105929), .A(n96394), .ZN(
        \DLX_Datapath/RegisterFile/N24968 ) );
  AOI22_X1 U83747 ( .A1(n69514), .A2(n105927), .B1(n105923), .B2(n81539), .ZN(
        n96394) );
  OAI21_X1 U83748 ( .B1(n106204), .B2(n105929), .A(n96395), .ZN(
        \DLX_Datapath/RegisterFile/N24966 ) );
  AOI22_X1 U83749 ( .A1(n74021), .A2(n105927), .B1(n105925), .B2(n81308), .ZN(
        n96395) );
  OAI21_X1 U83750 ( .B1(n106098), .B2(n105929), .A(n96396), .ZN(
        \DLX_Datapath/RegisterFile/N24965 ) );
  AOI22_X1 U83751 ( .A1(n105928), .A2(n108075), .B1(n94516), .B2(n105924), 
        .ZN(n96396) );
  OAI21_X1 U83752 ( .B1(n105992), .B2(n105929), .A(n96397), .ZN(
        \DLX_Datapath/RegisterFile/N24963 ) );
  AOI22_X1 U83753 ( .A1(n74302), .A2(n105927), .B1(n94519), .B2(n105924), .ZN(
        n96397) );
  OAI21_X1 U83754 ( .B1(n106333), .B2(n105929), .A(n96398), .ZN(
        \DLX_Datapath/RegisterFile/N24962 ) );
  AOI22_X1 U83755 ( .A1(n73738), .A2(n105927), .B1(n105925), .B2(n80192), .ZN(
        n96398) );
  OAI21_X1 U83756 ( .B1(n106190), .B2(n105929), .A(n96399), .ZN(
        \DLX_Datapath/RegisterFile/N24961 ) );
  AOI22_X1 U83757 ( .A1(n73442), .A2(n105927), .B1(n105923), .B2(n81474), .ZN(
        n96399) );
  OAI21_X1 U83758 ( .B1(n81383), .B2(n105929), .A(n96400), .ZN(
        \DLX_Datapath/RegisterFile/N24960 ) );
  AOI22_X1 U83759 ( .A1(n73879), .A2(n105927), .B1(n94523), .B2(n105924), .ZN(
        n96400) );
  OAI21_X1 U83760 ( .B1(n81318), .B2(n105929), .A(n96401), .ZN(
        \DLX_Datapath/RegisterFile/N24959 ) );
  AOI22_X1 U83761 ( .A1(n73591), .A2(n105927), .B1(n105925), .B2(n106061), 
        .ZN(n96401) );
  OAI21_X1 U83762 ( .B1(n81345), .B2(n105929), .A(n96402), .ZN(
        \DLX_Datapath/RegisterFile/N24958 ) );
  AOI22_X1 U83763 ( .A1(n105926), .A2(n110034), .B1(n105923), .B2(n81347), 
        .ZN(n96402) );
  OAI21_X1 U83764 ( .B1(n106103), .B2(n105929), .A(n96403), .ZN(
        \DLX_Datapath/RegisterFile/N24957 ) );
  AOI22_X1 U83765 ( .A1(n105928), .A2(n110141), .B1(n94527), .B2(n105924), 
        .ZN(n96403) );
  OAI21_X1 U83766 ( .B1(n81294), .B2(n105929), .A(n96404), .ZN(
        \DLX_Datapath/RegisterFile/N24956 ) );
  AOI22_X1 U83767 ( .A1(n105927), .A2(n109925), .B1(n105925), .B2(n81297), 
        .ZN(n96404) );
  OAI21_X1 U83768 ( .B1(n106110), .B2(n81745), .A(n96405), .ZN(
        \DLX_Datapath/RegisterFile/N24955 ) );
  AOI22_X1 U83769 ( .A1(n105928), .A2(n109807), .B1(n94530), .B2(n105924), 
        .ZN(n96405) );
  OAI21_X1 U83770 ( .B1(n106170), .B2(n81745), .A(n96406), .ZN(
        \DLX_Datapath/RegisterFile/N24953 ) );
  AOI22_X1 U83771 ( .A1(n105926), .A2(n108304), .B1(n105923), .B2(n106168), 
        .ZN(n96406) );
  OAI21_X1 U83772 ( .B1(n106070), .B2(n105929), .A(n96407), .ZN(
        \DLX_Datapath/RegisterFile/N24951 ) );
  AOI22_X1 U83773 ( .A1(n105926), .A2(n107653), .B1(n105925), .B2(n81453), 
        .ZN(n96407) );
  OAI21_X1 U83774 ( .B1(n106197), .B2(n81745), .A(n96408), .ZN(
        \DLX_Datapath/RegisterFile/N24950 ) );
  AOI22_X1 U83775 ( .A1(n105926), .A2(n109571), .B1(n94536), .B2(n105924), 
        .ZN(n96408) );
  OAI21_X1 U83776 ( .B1(n106157), .B2(n105929), .A(n96409), .ZN(
        \DLX_Datapath/RegisterFile/N24948 ) );
  AOI22_X1 U83777 ( .A1(n105928), .A2(n109676), .B1(n105923), .B2(n81351), 
        .ZN(n96409) );
  OAI21_X1 U83778 ( .B1(n106008), .B2(n81745), .A(n96410), .ZN(
        \DLX_Datapath/RegisterFile/N24946 ) );
  AOI22_X1 U83779 ( .A1(n105928), .A2(n108997), .B1(n94541), .B2(n105924), 
        .ZN(n96410) );
  OAI21_X1 U83780 ( .B1(n81509), .B2(n105929), .A(n96411), .ZN(
        \DLX_Datapath/RegisterFile/N24944 ) );
  AOI22_X1 U83781 ( .A1(n105926), .A2(n109227), .B1(n105624), .B2(n105923), 
        .ZN(n96411) );
  OAI21_X1 U83782 ( .B1(n106049), .B2(n81745), .A(n96412), .ZN(
        \DLX_Datapath/RegisterFile/N24943 ) );
  AOI22_X1 U83783 ( .A1(n105928), .A2(n109119), .B1(n94546), .B2(n105924), 
        .ZN(n96412) );
  OAI21_X1 U83784 ( .B1(n106095), .B2(n81745), .A(n96413), .ZN(
        \DLX_Datapath/RegisterFile/N24942 ) );
  AOI22_X1 U83785 ( .A1(n105926), .A2(n108654), .B1(n94548), .B2(n105924), 
        .ZN(n96413) );
  OAI21_X1 U83786 ( .B1(n106053), .B2(n81745), .A(n96414), .ZN(
        \DLX_Datapath/RegisterFile/N24941 ) );
  AOI22_X1 U83787 ( .A1(n105928), .A2(n108881), .B1(n81783), .B2(n105925), 
        .ZN(n96414) );
  OAI21_X1 U83788 ( .B1(n106267), .B2(n81745), .A(n96415), .ZN(
        \DLX_Datapath/RegisterFile/N24939 ) );
  AOI22_X1 U83789 ( .A1(n105928), .A2(n107309), .B1(n105925), .B2(n81265), 
        .ZN(n96415) );
  NOR2_X1 U83792 ( .A1(n81745), .A2(n105090), .ZN(n96417) );
  NAND2_X1 U83793 ( .A1(n96013), .A2(n105199), .ZN(n96010) );
  NAND2_X1 U83794 ( .A1(n105131), .A2(n94772), .ZN(n81745) );
  OAI21_X1 U83795 ( .B1(n81358), .B2(n105417), .A(n96419), .ZN(
        \DLX_Datapath/RegisterFile/N24938 ) );
  AOI22_X1 U83796 ( .A1(n105416), .A2(n70320), .B1(n104932), .B2(n94559), .ZN(
        n96419) );
  OAI21_X1 U83797 ( .B1(n105971), .B2(n105417), .A(n96422), .ZN(
        \DLX_Datapath/RegisterFile/N24937 ) );
  AOI22_X1 U83798 ( .A1(n105415), .A2(n70462), .B1(n104933), .B2(n94562), .ZN(
        n96422) );
  OAI21_X1 U83799 ( .B1(n106136), .B2(n105417), .A(n96423), .ZN(
        \DLX_Datapath/RegisterFile/N24936 ) );
  AOI22_X1 U83800 ( .A1(n105416), .A2(n69515), .B1(n104932), .B2(n94564), .ZN(
        n96423) );
  OAI21_X1 U83801 ( .B1(n106208), .B2(n105417), .A(n96424), .ZN(
        \DLX_Datapath/RegisterFile/N24935 ) );
  AOI22_X1 U83802 ( .A1(n105415), .A2(n70176), .B1(n104934), .B2(n94566), .ZN(
        n96424) );
  OAI21_X1 U83803 ( .B1(n106204), .B2(n105417), .A(n96425), .ZN(
        \DLX_Datapath/RegisterFile/N24934 ) );
  AOI22_X1 U83804 ( .A1(n105416), .A2(n74022), .B1(n104932), .B2(n94568), .ZN(
        n96425) );
  OAI21_X1 U83805 ( .B1(n106098), .B2(n105417), .A(n96426), .ZN(
        \DLX_Datapath/RegisterFile/N24933 ) );
  AOI22_X1 U83806 ( .A1(n105415), .A2(n70609), .B1(n104933), .B2(n94570), .ZN(
        n96426) );
  OAI21_X1 U83807 ( .B1(n81270), .B2(n105417), .A(n96427), .ZN(
        \DLX_Datapath/RegisterFile/N24932 ) );
  AOI22_X1 U83808 ( .A1(n105416), .A2(n74163), .B1(n104933), .B2(n94572), .ZN(
        n96427) );
  OAI21_X1 U83809 ( .B1(n105992), .B2(n105417), .A(n96428), .ZN(
        \DLX_Datapath/RegisterFile/N24931 ) );
  AOI22_X1 U83810 ( .A1(n105415), .A2(n74303), .B1(n104934), .B2(n94574), .ZN(
        n96428) );
  OAI21_X1 U83811 ( .B1(n106333), .B2(n105417), .A(n96429), .ZN(
        \DLX_Datapath/RegisterFile/N24930 ) );
  AOI22_X1 U83812 ( .A1(n105415), .A2(n73739), .B1(n104933), .B2(n94576), .ZN(
        n96429) );
  OAI21_X1 U83813 ( .B1(n106190), .B2(n105417), .A(n96430), .ZN(
        \DLX_Datapath/RegisterFile/N24929 ) );
  AOI22_X1 U83814 ( .A1(n105414), .A2(n73443), .B1(n104932), .B2(n94578), .ZN(
        n96430) );
  OAI21_X1 U83815 ( .B1(n81383), .B2(n105417), .A(n96431), .ZN(
        \DLX_Datapath/RegisterFile/N24928 ) );
  AOI22_X1 U83816 ( .A1(n105414), .A2(n73880), .B1(n104933), .B2(n94580), .ZN(
        n96431) );
  OAI21_X1 U83817 ( .B1(n81318), .B2(n105417), .A(n96432), .ZN(
        \DLX_Datapath/RegisterFile/N24927 ) );
  AOI22_X1 U83818 ( .A1(n105414), .A2(n73592), .B1(n104934), .B2(n94582), .ZN(
        n96432) );
  OAI21_X1 U83819 ( .B1(n81345), .B2(n105417), .A(n96433), .ZN(
        \DLX_Datapath/RegisterFile/N24926 ) );
  AOI22_X1 U83820 ( .A1(n105414), .A2(n73154), .B1(n104934), .B2(n94584), .ZN(
        n96433) );
  OAI21_X1 U83821 ( .B1(n106103), .B2(n105417), .A(n96434), .ZN(
        \DLX_Datapath/RegisterFile/N24925 ) );
  AOI22_X1 U83822 ( .A1(n105414), .A2(n73296), .B1(n104932), .B2(n94586), .ZN(
        n96434) );
  OAI21_X1 U83823 ( .B1(n81294), .B2(n105417), .A(n96435), .ZN(
        \DLX_Datapath/RegisterFile/N24924 ) );
  AOI22_X1 U83824 ( .A1(n105414), .A2(n73012), .B1(n104932), .B2(n94588), .ZN(
        n96435) );
  OAI21_X1 U83825 ( .B1(n106108), .B2(n105417), .A(n96436), .ZN(
        \DLX_Datapath/RegisterFile/N24923 ) );
  AOI22_X1 U83826 ( .A1(n105414), .A2(n72862), .B1(n104933), .B2(n94590), .ZN(
        n96436) );
  OAI21_X1 U83827 ( .B1(n106231), .B2(n105417), .A(n96437), .ZN(
        \DLX_Datapath/RegisterFile/N24922 ) );
  AOI22_X1 U83828 ( .A1(n105414), .A2(n70758), .B1(n104934), .B2(n94592), .ZN(
        n96437) );
  OAI21_X1 U83829 ( .B1(n106170), .B2(n105417), .A(n96438), .ZN(
        \DLX_Datapath/RegisterFile/N24921 ) );
  AOI22_X1 U83830 ( .A1(n105414), .A2(n70917), .B1(n104933), .B2(n94594), .ZN(
        n96438) );
  OAI21_X1 U83831 ( .B1(n106236), .B2(n105417), .A(n96439), .ZN(
        \DLX_Datapath/RegisterFile/N24920 ) );
  AOI22_X1 U83832 ( .A1(n105414), .A2(n71062), .B1(n104932), .B2(n94596), .ZN(
        n96439) );
  OAI21_X1 U83833 ( .B1(n106071), .B2(n105417), .A(n96440), .ZN(
        \DLX_Datapath/RegisterFile/N24919 ) );
  AOI22_X1 U83834 ( .A1(n105414), .A2(n70023), .B1(n104933), .B2(n94598), .ZN(
        n96440) );
  OAI21_X1 U83835 ( .B1(n106197), .B2(n105417), .A(n96441), .ZN(
        \DLX_Datapath/RegisterFile/N24918 ) );
  AOI22_X1 U83836 ( .A1(n105415), .A2(n72552), .B1(n104934), .B2(n94600), .ZN(
        n96441) );
  OAI21_X1 U83837 ( .B1(n81278), .B2(n105417), .A(n96442), .ZN(
        \DLX_Datapath/RegisterFile/N24917 ) );
  AOI22_X1 U83838 ( .A1(n105416), .A2(n71211), .B1(n104934), .B2(n94602), .ZN(
        n96442) );
  OAI21_X1 U83839 ( .B1(n106157), .B2(n96418), .A(n96443), .ZN(
        \DLX_Datapath/RegisterFile/N24916 ) );
  AOI22_X1 U83840 ( .A1(n105415), .A2(n72694), .B1(n104934), .B2(n94604), .ZN(
        n96443) );
  OAI21_X1 U83841 ( .B1(n106115), .B2(n96418), .A(n96444), .ZN(
        \DLX_Datapath/RegisterFile/N24915 ) );
  AOI22_X1 U83842 ( .A1(n105416), .A2(n72404), .B1(n104932), .B2(n94606), .ZN(
        n96444) );
  OAI21_X1 U83843 ( .B1(n106008), .B2(n96418), .A(n96445), .ZN(
        \DLX_Datapath/RegisterFile/N24914 ) );
  AOI22_X1 U83844 ( .A1(n105415), .A2(n71804), .B1(n104932), .B2(n94608), .ZN(
        n96445) );
  OAI21_X1 U83845 ( .B1(n106259), .B2(n96418), .A(n96446), .ZN(
        \DLX_Datapath/RegisterFile/N24913 ) );
  AOI22_X1 U83846 ( .A1(n105416), .A2(n72253), .B1(n104933), .B2(n94610), .ZN(
        n96446) );
  OAI21_X1 U83847 ( .B1(n81509), .B2(n105417), .A(n96447), .ZN(
        \DLX_Datapath/RegisterFile/N24912 ) );
  AOI22_X1 U83848 ( .A1(n105415), .A2(n72102), .B1(n104934), .B2(n94612), .ZN(
        n96447) );
  OAI21_X1 U83849 ( .B1(n106049), .B2(n96418), .A(n96448), .ZN(
        \DLX_Datapath/RegisterFile/N24911 ) );
  AOI22_X1 U83850 ( .A1(n105416), .A2(n71958), .B1(n104933), .B2(n94614), .ZN(
        n96448) );
  OAI21_X1 U83851 ( .B1(n106096), .B2(n96418), .A(n96449), .ZN(
        \DLX_Datapath/RegisterFile/N24910 ) );
  AOI22_X1 U83852 ( .A1(n105415), .A2(n71360), .B1(n104932), .B2(n94616), .ZN(
        n96449) );
  OAI21_X1 U83853 ( .B1(n106053), .B2(n96418), .A(n96450), .ZN(
        \DLX_Datapath/RegisterFile/N24909 ) );
  AOI22_X1 U83854 ( .A1(n105416), .A2(n71655), .B1(n104933), .B2(n94618), .ZN(
        n96450) );
  OAI21_X1 U83855 ( .B1(n105219), .B2(n105417), .A(n96451), .ZN(
        \DLX_Datapath/RegisterFile/N24908 ) );
  AOI22_X1 U83856 ( .A1(n105416), .A2(n71511), .B1(n104932), .B2(n94620), .ZN(
        n96451) );
  OAI21_X1 U83857 ( .B1(n106267), .B2(n96418), .A(n96452), .ZN(
        \DLX_Datapath/RegisterFile/N24907 ) );
  AOI22_X1 U83858 ( .A1(n105415), .A2(n69620), .B1(n104934), .B2(n94622), .ZN(
        n96452) );
  NOR2_X1 U83861 ( .A1(n96418), .A2(n105090), .ZN(n96453) );
  NAND2_X1 U83862 ( .A1(n105132), .A2(n94810), .ZN(n96418) );
  OAI21_X1 U83863 ( .B1(n106147), .B2(n81628), .A(n96455), .ZN(
        \DLX_Datapath/RegisterFile/N24906 ) );
  AOI22_X1 U83864 ( .A1(n105987), .A2(n81521), .B1(n70321), .B2(n105984), .ZN(
        n96455) );
  OAI21_X1 U83865 ( .B1(n81628), .B2(n81651), .A(n96456), .ZN(
        \DLX_Datapath/RegisterFile/N24905 ) );
  AOI22_X1 U83866 ( .A1(n81653), .A2(n105988), .B1(n70463), .B2(n105984), .ZN(
        n96456) );
  OAI21_X1 U83867 ( .B1(n106136), .B2(n81628), .A(n96457), .ZN(
        \DLX_Datapath/RegisterFile/N24904 ) );
  AOI22_X1 U83868 ( .A1(n105989), .A2(n81380), .B1(n105985), .B2(n107235), 
        .ZN(n96457) );
  OAI21_X1 U83869 ( .B1(n81299), .B2(n105994), .A(n96458), .ZN(
        \DLX_Datapath/RegisterFile/N24903 ) );
  AOI22_X1 U83870 ( .A1(n105987), .A2(n81377), .B1(n105986), .B2(n107774), 
        .ZN(n96458) );
  OAI21_X1 U83871 ( .B1(n106204), .B2(n81628), .A(n96459), .ZN(
        \DLX_Datapath/RegisterFile/N24902 ) );
  AOI22_X1 U83872 ( .A1(n105989), .A2(n81428), .B1(n105985), .B2(n110676), 
        .ZN(n96459) );
  OAI21_X1 U83873 ( .B1(n106098), .B2(n81628), .A(n96460), .ZN(
        \DLX_Datapath/RegisterFile/N24901 ) );
  AOI22_X1 U83874 ( .A1(n105987), .A2(n81410), .B1(n105986), .B2(n108076), 
        .ZN(n96460) );
  OAI21_X1 U83875 ( .B1(n81270), .B2(n105994), .A(n96461), .ZN(
        \DLX_Datapath/RegisterFile/N24900 ) );
  AOI22_X1 U83876 ( .A1(n81700), .A2(n105988), .B1(n105985), .B2(n110773), 
        .ZN(n96461) );
  OAI21_X1 U83877 ( .B1(n106333), .B2(n105994), .A(n96462), .ZN(
        \DLX_Datapath/RegisterFile/N24898 ) );
  AOI22_X1 U83878 ( .A1(n105988), .A2(n81414), .B1(n105984), .B2(n110469), 
        .ZN(n96462) );
  OAI21_X1 U83879 ( .B1(n106190), .B2(n81628), .A(n96463), .ZN(
        \DLX_Datapath/RegisterFile/N24897 ) );
  AOI22_X1 U83880 ( .A1(n105987), .A2(n81317), .B1(n105985), .B2(n110251), 
        .ZN(n96463) );
  OAI21_X1 U83881 ( .B1(n81383), .B2(n105994), .A(n96464), .ZN(
        \DLX_Datapath/RegisterFile/N24896 ) );
  AOI22_X1 U83882 ( .A1(n105987), .A2(n81386), .B1(n105985), .B2(n110568), 
        .ZN(n96464) );
  OAI21_X1 U83883 ( .B1(n81318), .B2(n105994), .A(n96465), .ZN(
        \DLX_Datapath/RegisterFile/N24895 ) );
  AOI22_X1 U83884 ( .A1(n105988), .A2(n81320), .B1(n105984), .B2(n110359), 
        .ZN(n96465) );
  OAI21_X1 U83885 ( .B1(n106162), .B2(n105994), .A(n96466), .ZN(
        \DLX_Datapath/RegisterFile/N24894 ) );
  AOI22_X1 U83886 ( .A1(n105989), .A2(n81604), .B1(n105986), .B2(n110035), 
        .ZN(n96466) );
  OAI21_X1 U83887 ( .B1(n106103), .B2(n105994), .A(n96467), .ZN(
        \DLX_Datapath/RegisterFile/N24893 ) );
  AOI22_X1 U83888 ( .A1(n105987), .A2(n81405), .B1(n105985), .B2(n110142), 
        .ZN(n96467) );
  OAI21_X1 U83889 ( .B1(n106220), .B2(n105994), .A(n96468), .ZN(
        \DLX_Datapath/RegisterFile/N24892 ) );
  AOI22_X1 U83890 ( .A1(n105989), .A2(n81402), .B1(n105986), .B2(n109926), 
        .ZN(n96468) );
  OAI21_X1 U83891 ( .B1(n106108), .B2(n105994), .A(n96469), .ZN(
        \DLX_Datapath/RegisterFile/N24891 ) );
  AOI22_X1 U83892 ( .A1(n105988), .A2(n81400), .B1(n105984), .B2(n109808), 
        .ZN(n96469) );
  OAI21_X1 U83893 ( .B1(n106231), .B2(n105994), .A(n96470), .ZN(
        \DLX_Datapath/RegisterFile/N24890 ) );
  AOI22_X1 U83894 ( .A1(n105989), .A2(n81332), .B1(n105986), .B2(n108182), 
        .ZN(n96470) );
  OAI21_X1 U83895 ( .B1(n106170), .B2(n105994), .A(n96471), .ZN(
        \DLX_Datapath/RegisterFile/N24889 ) );
  AOI22_X1 U83896 ( .A1(n105988), .A2(n81373), .B1(n105984), .B2(n108305), 
        .ZN(n96471) );
  OAI21_X1 U83897 ( .B1(n81281), .B2(n105994), .A(n96472), .ZN(
        \DLX_Datapath/RegisterFile/N24888 ) );
  AOI22_X1 U83898 ( .A1(n105988), .A2(n81322), .B1(n105984), .B2(n108416), 
        .ZN(n96472) );
  OAI21_X1 U83899 ( .B1(n106071), .B2(n105994), .A(n96473), .ZN(
        \DLX_Datapath/RegisterFile/N24887 ) );
  AOI22_X1 U83900 ( .A1(n105988), .A2(n81506), .B1(n105984), .B2(n107654), 
        .ZN(n96473) );
  OAI21_X1 U83901 ( .B1(n106197), .B2(n105994), .A(n96474), .ZN(
        \DLX_Datapath/RegisterFile/N24886 ) );
  AOI22_X1 U83902 ( .A1(n105988), .A2(n81313), .B1(n105984), .B2(n109572), 
        .ZN(n96474) );
  OAI21_X1 U83903 ( .B1(n81278), .B2(n105994), .A(n96475), .ZN(
        \DLX_Datapath/RegisterFile/N24885 ) );
  AOI22_X1 U83904 ( .A1(n105988), .A2(n81330), .B1(n105984), .B2(n108533), 
        .ZN(n96475) );
  OAI21_X1 U83905 ( .B1(n106157), .B2(n105994), .A(n96476), .ZN(
        \DLX_Datapath/RegisterFile/N24884 ) );
  AOI22_X1 U83906 ( .A1(n105989), .A2(n81425), .B1(n105986), .B2(n109677), 
        .ZN(n96476) );
  OAI21_X1 U83907 ( .B1(n106116), .B2(n105994), .A(n96477), .ZN(
        \DLX_Datapath/RegisterFile/N24883 ) );
  AOI22_X1 U83908 ( .A1(n105989), .A2(n81396), .B1(n105986), .B2(n109461), 
        .ZN(n96477) );
  OAI21_X1 U83909 ( .B1(n106008), .B2(n105994), .A(n96478), .ZN(
        \DLX_Datapath/RegisterFile/N24882 ) );
  AOI22_X1 U83910 ( .A1(n105987), .A2(n81590), .B1(n105985), .B2(n108998), 
        .ZN(n96478) );
  OAI21_X1 U83911 ( .B1(n106260), .B2(n105994), .A(n96479), .ZN(
        \DLX_Datapath/RegisterFile/N24881 ) );
  AOI22_X1 U83912 ( .A1(n105987), .A2(n81423), .B1(n105985), .B2(n109346), 
        .ZN(n96479) );
  OAI21_X1 U83913 ( .B1(n106045), .B2(n105994), .A(n96480), .ZN(
        \DLX_Datapath/RegisterFile/N24880 ) );
  AOI22_X1 U83914 ( .A1(n105989), .A2(n81511), .B1(n105986), .B2(n109228), 
        .ZN(n96480) );
  OAI21_X1 U83915 ( .B1(n106049), .B2(n105994), .A(n96481), .ZN(
        \DLX_Datapath/RegisterFile/N24879 ) );
  AOI22_X1 U83916 ( .A1(n105987), .A2(n81503), .B1(n105985), .B2(n109120), 
        .ZN(n96481) );
  OAI21_X1 U83917 ( .B1(n81415), .B2(n105994), .A(n96482), .ZN(
        \DLX_Datapath/RegisterFile/N24878 ) );
  AOI22_X1 U83918 ( .A1(n105989), .A2(n81417), .B1(n105986), .B2(n108655), 
        .ZN(n96482) );
  OAI21_X1 U83919 ( .B1(n106053), .B2(n105994), .A(n96483), .ZN(
        \DLX_Datapath/RegisterFile/N24877 ) );
  AOI22_X1 U83920 ( .A1(n105987), .A2(n81500), .B1(n105985), .B2(n108882), 
        .ZN(n96483) );
  OAI21_X1 U83921 ( .B1(n105219), .B2(n105994), .A(n96484), .ZN(
        \DLX_Datapath/RegisterFile/N24876 ) );
  AOI22_X1 U83922 ( .A1(n105989), .A2(n81335), .B1(n105986), .B2(n108770), 
        .ZN(n96484) );
  OAI21_X1 U83923 ( .B1(n106267), .B2(n81628), .A(n96485), .ZN(
        \DLX_Datapath/RegisterFile/N24875 ) );
  AOI22_X1 U83924 ( .A1(n105989), .A2(n81327), .B1(n105986), .B2(n107310), 
        .ZN(n96485) );
  AOI21_X1 U83926 ( .B1(n105205), .B2(n96416), .A(n105601), .ZN(n96454) );
  NOR2_X1 U83928 ( .A1(n81628), .A2(n105090), .ZN(n96486) );
  OR2_X1 U83929 ( .A1(n96013), .A2(n94848), .ZN(n96416) );
  NAND2_X1 U83930 ( .A1(n96487), .A2(n94850), .ZN(n96013) );
  AND2_X2 U83931 ( .A1(n96488), .A2(n96489), .ZN(n94850) );
  NOR2_X1 U83932 ( .A1(n107028), .A2(n106763), .ZN(n96487) );
  NAND2_X1 U83933 ( .A1(n105131), .A2(n94853), .ZN(n81628) );
  OAI21_X1 U83934 ( .B1(n106147), .B2(n105413), .A(n96491), .ZN(
        \DLX_Datapath/RegisterFile/N24874 ) );
  AOI22_X1 U83935 ( .A1(n105412), .A2(n94667), .B1(n96493), .B2(n107875), .ZN(
        n96491) );
  OAI21_X1 U83936 ( .B1(n105971), .B2(n105413), .A(n96494), .ZN(
        \DLX_Datapath/RegisterFile/N24873 ) );
  AOI22_X1 U83937 ( .A1(n105411), .A2(n94670), .B1(n104967), .B2(n107972), 
        .ZN(n96494) );
  OAI21_X1 U83938 ( .B1(n106136), .B2(n105413), .A(n96495), .ZN(
        \DLX_Datapath/RegisterFile/N24872 ) );
  AOI22_X1 U83939 ( .A1(n105412), .A2(n94672), .B1(n96493), .B2(n107236), .ZN(
        n96495) );
  OAI21_X1 U83940 ( .B1(n81299), .B2(n105413), .A(n96496), .ZN(
        \DLX_Datapath/RegisterFile/N24871 ) );
  AOI22_X1 U83941 ( .A1(n105411), .A2(n94674), .B1(n104968), .B2(n107775), 
        .ZN(n96496) );
  OAI21_X1 U83942 ( .B1(n81306), .B2(n105413), .A(n96497), .ZN(
        \DLX_Datapath/RegisterFile/N24870 ) );
  AOI22_X1 U83943 ( .A1(n105412), .A2(n94676), .B1(n104967), .B2(n110677), 
        .ZN(n96497) );
  OAI21_X1 U83944 ( .B1(n106098), .B2(n105413), .A(n96498), .ZN(
        \DLX_Datapath/RegisterFile/N24869 ) );
  AOI22_X1 U83945 ( .A1(n105411), .A2(n94678), .B1(n104967), .B2(n108077), 
        .ZN(n96498) );
  OAI21_X1 U83946 ( .B1(n106256), .B2(n105413), .A(n96499), .ZN(
        \DLX_Datapath/RegisterFile/N24868 ) );
  AOI22_X1 U83947 ( .A1(n105412), .A2(n94680), .B1(n104967), .B2(n110774), 
        .ZN(n96499) );
  OAI21_X1 U83948 ( .B1(n105992), .B2(n105413), .A(n96500), .ZN(
        \DLX_Datapath/RegisterFile/N24867 ) );
  AOI22_X1 U83949 ( .A1(n105411), .A2(n94682), .B1(n104968), .B2(n110875), 
        .ZN(n96500) );
  OAI21_X1 U83950 ( .B1(n106333), .B2(n105413), .A(n96501), .ZN(
        \DLX_Datapath/RegisterFile/N24866 ) );
  AOI22_X1 U83951 ( .A1(n105411), .A2(n94684), .B1(n104967), .B2(n110470), 
        .ZN(n96501) );
  OAI21_X1 U83952 ( .B1(n106190), .B2(n105413), .A(n96502), .ZN(
        \DLX_Datapath/RegisterFile/N24865 ) );
  AOI22_X1 U83953 ( .A1(n105410), .A2(n94686), .B1(n96493), .B2(n110252), .ZN(
        n96502) );
  OAI21_X1 U83954 ( .B1(n81383), .B2(n105413), .A(n96503), .ZN(
        \DLX_Datapath/RegisterFile/N24864 ) );
  AOI22_X1 U83955 ( .A1(n105410), .A2(n94688), .B1(n104967), .B2(n110569), 
        .ZN(n96503) );
  OAI21_X1 U83956 ( .B1(n106187), .B2(n105413), .A(n96504), .ZN(
        \DLX_Datapath/RegisterFile/N24863 ) );
  AOI22_X1 U83957 ( .A1(n105410), .A2(n94690), .B1(n104968), .B2(n110360), 
        .ZN(n96504) );
  OAI21_X1 U83958 ( .B1(n106162), .B2(n105413), .A(n96505), .ZN(
        \DLX_Datapath/RegisterFile/N24862 ) );
  AOI22_X1 U83959 ( .A1(n105410), .A2(n94692), .B1(n104968), .B2(n110036), 
        .ZN(n96505) );
  OAI21_X1 U83960 ( .B1(n106103), .B2(n105413), .A(n96506), .ZN(
        \DLX_Datapath/RegisterFile/N24861 ) );
  AOI22_X1 U83961 ( .A1(n105410), .A2(n94694), .B1(n104967), .B2(n110143), 
        .ZN(n96506) );
  OAI21_X1 U83962 ( .B1(n81294), .B2(n105413), .A(n96507), .ZN(
        \DLX_Datapath/RegisterFile/N24860 ) );
  AOI22_X1 U83963 ( .A1(n105410), .A2(n94696), .B1(n104968), .B2(n109927), 
        .ZN(n96507) );
  OAI21_X1 U83964 ( .B1(n106111), .B2(n105413), .A(n96508), .ZN(
        \DLX_Datapath/RegisterFile/N24859 ) );
  AOI22_X1 U83965 ( .A1(n105410), .A2(n94698), .B1(n104967), .B2(n109809), 
        .ZN(n96508) );
  OAI21_X1 U83966 ( .B1(n106231), .B2(n105413), .A(n96509), .ZN(
        \DLX_Datapath/RegisterFile/N24858 ) );
  AOI22_X1 U83967 ( .A1(n105410), .A2(n94700), .B1(n104968), .B2(n108183), 
        .ZN(n96509) );
  OAI21_X1 U83968 ( .B1(n106170), .B2(n105413), .A(n96510), .ZN(
        \DLX_Datapath/RegisterFile/N24857 ) );
  AOI22_X1 U83969 ( .A1(n105410), .A2(n94702), .B1(n104967), .B2(n108306), 
        .ZN(n96510) );
  OAI21_X1 U83970 ( .B1(n106238), .B2(n105413), .A(n96511), .ZN(
        \DLX_Datapath/RegisterFile/N24856 ) );
  AOI22_X1 U83971 ( .A1(n105410), .A2(n94704), .B1(n96493), .B2(n108417), .ZN(
        n96511) );
  OAI21_X1 U83972 ( .B1(n106071), .B2(n105413), .A(n96512), .ZN(
        \DLX_Datapath/RegisterFile/N24855 ) );
  AOI22_X1 U83973 ( .A1(n105410), .A2(n94706), .B1(n104967), .B2(n107655), 
        .ZN(n96512) );
  OAI21_X1 U83974 ( .B1(n106197), .B2(n105413), .A(n96513), .ZN(
        \DLX_Datapath/RegisterFile/N24854 ) );
  AOI22_X1 U83975 ( .A1(n105411), .A2(n94708), .B1(n104968), .B2(n109573), 
        .ZN(n96513) );
  OAI21_X1 U83976 ( .B1(n81278), .B2(n105413), .A(n96514), .ZN(
        \DLX_Datapath/RegisterFile/N24853 ) );
  AOI22_X1 U83977 ( .A1(n105411), .A2(n94710), .B1(n104968), .B2(n108534), 
        .ZN(n96514) );
  OAI21_X1 U83978 ( .B1(n106157), .B2(n105413), .A(n96515), .ZN(
        \DLX_Datapath/RegisterFile/N24852 ) );
  AOI22_X1 U83979 ( .A1(n105412), .A2(n94712), .B1(n104968), .B2(n109678), 
        .ZN(n96515) );
  OAI21_X1 U83980 ( .B1(n106115), .B2(n105413), .A(n96516), .ZN(
        \DLX_Datapath/RegisterFile/N24851 ) );
  AOI22_X1 U83981 ( .A1(n105411), .A2(n94714), .B1(n96493), .B2(n109462), .ZN(
        n96516) );
  OAI21_X1 U83982 ( .B1(n106008), .B2(n105413), .A(n96517), .ZN(
        \DLX_Datapath/RegisterFile/N24850 ) );
  AOI22_X1 U83983 ( .A1(n105412), .A2(n81259), .B1(n96493), .B2(n108999), .ZN(
        n96517) );
  OAI21_X1 U83984 ( .B1(n106259), .B2(n105413), .A(n96518), .ZN(
        \DLX_Datapath/RegisterFile/N24849 ) );
  AOI22_X1 U83985 ( .A1(n105411), .A2(n94717), .B1(n104967), .B2(n109347), 
        .ZN(n96518) );
  OAI21_X1 U83986 ( .B1(n106043), .B2(n105413), .A(n96519), .ZN(
        \DLX_Datapath/RegisterFile/N24848 ) );
  AOI22_X1 U83987 ( .A1(n105412), .A2(n94719), .B1(n104968), .B2(n109229), 
        .ZN(n96519) );
  OAI21_X1 U83988 ( .B1(n106049), .B2(n105413), .A(n96520), .ZN(
        \DLX_Datapath/RegisterFile/N24847 ) );
  AOI22_X1 U83989 ( .A1(n105411), .A2(n94721), .B1(n104967), .B2(n109121), 
        .ZN(n96520) );
  OAI21_X1 U83990 ( .B1(n81415), .B2(n105413), .A(n96521), .ZN(
        \DLX_Datapath/RegisterFile/N24846 ) );
  AOI22_X1 U83991 ( .A1(n105412), .A2(n94723), .B1(n104967), .B2(n108656), 
        .ZN(n96521) );
  OAI21_X1 U83992 ( .B1(n106053), .B2(n105413), .A(n96522), .ZN(
        \DLX_Datapath/RegisterFile/N24845 ) );
  AOI22_X1 U83993 ( .A1(n105411), .A2(n94725), .B1(n104967), .B2(n108883), 
        .ZN(n96522) );
  OAI21_X1 U83994 ( .B1(n105219), .B2(n105413), .A(n96523), .ZN(
        \DLX_Datapath/RegisterFile/N24844 ) );
  AOI22_X1 U83995 ( .A1(n105412), .A2(n94727), .B1(n96493), .B2(n108771), .ZN(
        n96523) );
  OAI21_X1 U83996 ( .B1(n106267), .B2(n105413), .A(n96524), .ZN(
        \DLX_Datapath/RegisterFile/N24843 ) );
  AOI22_X1 U83997 ( .A1(n105412), .A2(n94729), .B1(n104968), .B2(n107311), 
        .ZN(n96524) );
  AOI21_X1 U83998 ( .B1(n96525), .B2(n105602), .A(n96526), .ZN(n96493) );
  OAI21_X1 U83999 ( .B1(n106757), .B2(n94848), .A(n107022), .ZN(n96525) );
  NOR2_X1 U84001 ( .A1(n96528), .A2(n106763), .ZN(n96130) );
  NAND2_X1 U84002 ( .A1(n94852), .A2(n59515), .ZN(n96528) );
  OR2_X1 U84003 ( .A1(n96526), .A2(n94848), .ZN(n96527) );
  NOR2_X1 U84004 ( .A1(n104503), .A2(n105091), .ZN(n96526) );
  NOR2_X1 U84006 ( .A1(n94894), .A2(n96529), .ZN(n96014) );
  NAND2_X1 U84007 ( .A1(n96530), .A2(n96531), .ZN(n94894) );
  OAI21_X1 U84008 ( .B1(n106147), .B2(n106028), .A(n96532), .ZN(
        \DLX_Datapath/RegisterFile/N24842 ) );
  AOI22_X1 U84009 ( .A1(n106027), .A2(n107876), .B1(n104789), .B2(n81360), 
        .ZN(n96532) );
  OAI21_X1 U84010 ( .B1(n106028), .B2(n81651), .A(n96533), .ZN(
        \DLX_Datapath/RegisterFile/N24841 ) );
  AOI22_X1 U84011 ( .A1(n106026), .A2(n107973), .B1(n94511), .B2(n104789), 
        .ZN(n96533) );
  OAI21_X1 U84012 ( .B1(n106136), .B2(n106028), .A(n96534), .ZN(
        \DLX_Datapath/RegisterFile/N24840 ) );
  AOI22_X1 U84013 ( .A1(n106026), .A2(n107237), .B1(n81557), .B2(n81539), .ZN(
        n96534) );
  OAI21_X1 U84014 ( .B1(n81306), .B2(n106028), .A(n96535), .ZN(
        \DLX_Datapath/RegisterFile/N24838 ) );
  AOI22_X1 U84015 ( .A1(n106026), .A2(n110678), .B1(n104789), .B2(n81308), 
        .ZN(n96535) );
  OAI21_X1 U84016 ( .B1(n106098), .B2(n106028), .A(n96536), .ZN(
        \DLX_Datapath/RegisterFile/N24837 ) );
  AOI22_X1 U84017 ( .A1(n81556), .A2(n108078), .B1(n94516), .B2(n104789), .ZN(
        n96536) );
  OAI21_X1 U84018 ( .B1(n81270), .B2(n106028), .A(n96537), .ZN(
        \DLX_Datapath/RegisterFile/N24836 ) );
  AOI22_X1 U84019 ( .A1(n106026), .A2(n110775), .B1(n104789), .B2(n81272), 
        .ZN(n96537) );
  OAI21_X1 U84020 ( .B1(n106028), .B2(n105992), .A(n96538), .ZN(
        \DLX_Datapath/RegisterFile/N24835 ) );
  AOI22_X1 U84021 ( .A1(n106026), .A2(n110876), .B1(n94519), .B2(n81557), .ZN(
        n96538) );
  OAI21_X1 U84022 ( .B1(n106333), .B2(n106028), .A(n96539), .ZN(
        \DLX_Datapath/RegisterFile/N24834 ) );
  AOI22_X1 U84023 ( .A1(n106026), .A2(n110471), .B1(n104790), .B2(n80192), 
        .ZN(n96539) );
  OAI21_X1 U84024 ( .B1(n81315), .B2(n106028), .A(n96540), .ZN(
        \DLX_Datapath/RegisterFile/N24833 ) );
  AOI22_X1 U84025 ( .A1(n106026), .A2(n110253), .B1(n81557), .B2(n81474), .ZN(
        n96540) );
  OAI21_X1 U84026 ( .B1(n81383), .B2(n106028), .A(n96541), .ZN(
        \DLX_Datapath/RegisterFile/N24832 ) );
  AOI22_X1 U84027 ( .A1(n106026), .A2(n110570), .B1(n94523), .B2(n81557), .ZN(
        n96541) );
  OAI21_X1 U84028 ( .B1(n106103), .B2(n106028), .A(n96542), .ZN(
        \DLX_Datapath/RegisterFile/N24829 ) );
  AOI22_X1 U84029 ( .A1(n81556), .A2(n110144), .B1(n94527), .B2(n104790), .ZN(
        n96542) );
  OAI21_X1 U84030 ( .B1(n106221), .B2(n106028), .A(n96543), .ZN(
        \DLX_Datapath/RegisterFile/N24828 ) );
  AOI22_X1 U84031 ( .A1(n106026), .A2(n109928), .B1(n81557), .B2(n81297), .ZN(
        n96543) );
  OAI21_X1 U84032 ( .B1(n81398), .B2(n106028), .A(n96544), .ZN(
        \DLX_Datapath/RegisterFile/N24827 ) );
  AOI22_X1 U84033 ( .A1(n81556), .A2(n109810), .B1(n94530), .B2(n104790), .ZN(
        n96544) );
  OAI21_X1 U84034 ( .B1(n106170), .B2(n106028), .A(n96545), .ZN(
        \DLX_Datapath/RegisterFile/N24825 ) );
  AOI22_X1 U84035 ( .A1(n106026), .A2(n108307), .B1(n81557), .B2(n106168), 
        .ZN(n96545) );
  OAI21_X1 U84036 ( .B1(n106071), .B2(n106028), .A(n96546), .ZN(
        \DLX_Datapath/RegisterFile/N24823 ) );
  AOI22_X1 U84037 ( .A1(n106026), .A2(n107656), .B1(n104790), .B2(n81453), 
        .ZN(n96546) );
  OAI21_X1 U84038 ( .B1(n106197), .B2(n106028), .A(n96547), .ZN(
        \DLX_Datapath/RegisterFile/N24822 ) );
  AOI22_X1 U84039 ( .A1(n106026), .A2(n109574), .B1(n94536), .B2(n81557), .ZN(
        n96547) );
  OAI21_X1 U84040 ( .B1(n106157), .B2(n106028), .A(n96548), .ZN(
        \DLX_Datapath/RegisterFile/N24820 ) );
  AOI22_X1 U84041 ( .A1(n106026), .A2(n109679), .B1(n81557), .B2(n81351), .ZN(
        n96548) );
  OAI21_X1 U84042 ( .B1(n106116), .B2(n106028), .A(n96549), .ZN(
        \DLX_Datapath/RegisterFile/N24819 ) );
  AOI22_X1 U84043 ( .A1(n106026), .A2(n109463), .B1(n106021), .B2(n104789), 
        .ZN(n96549) );
  OAI21_X1 U84044 ( .B1(n106008), .B2(n106028), .A(n96550), .ZN(
        \DLX_Datapath/RegisterFile/N24818 ) );
  AOI22_X1 U84045 ( .A1(n106026), .A2(n109000), .B1(n94541), .B2(n104790), 
        .ZN(n96550) );
  OAI21_X1 U84046 ( .B1(n106046), .B2(n106028), .A(n96551), .ZN(
        \DLX_Datapath/RegisterFile/N24816 ) );
  AOI22_X1 U84047 ( .A1(n106026), .A2(n109230), .B1(n105625), .B2(n104789), 
        .ZN(n96551) );
  OAI21_X1 U84048 ( .B1(n106049), .B2(n106028), .A(n96552), .ZN(
        \DLX_Datapath/RegisterFile/N24815 ) );
  AOI22_X1 U84049 ( .A1(n106026), .A2(n109122), .B1(n94546), .B2(n104789), 
        .ZN(n96552) );
  OAI21_X1 U84050 ( .B1(n81415), .B2(n106028), .A(n96553), .ZN(
        \DLX_Datapath/RegisterFile/N24814 ) );
  AOI22_X1 U84051 ( .A1(n106026), .A2(n108657), .B1(n94548), .B2(n104790), 
        .ZN(n96553) );
  OAI21_X1 U84052 ( .B1(n106053), .B2(n106028), .A(n96554), .ZN(
        \DLX_Datapath/RegisterFile/N24813 ) );
  AOI22_X1 U84053 ( .A1(n106026), .A2(n108884), .B1(n81783), .B2(n104790), 
        .ZN(n96554) );
  OAI21_X1 U84054 ( .B1(n105219), .B2(n106028), .A(n96555), .ZN(
        \DLX_Datapath/RegisterFile/N24812 ) );
  AOI22_X1 U84055 ( .A1(n106026), .A2(n108772), .B1(n81557), .B2(n80188), .ZN(
        n96555) );
  OAI21_X1 U84056 ( .B1(n106267), .B2(n106028), .A(n96556), .ZN(
        \DLX_Datapath/RegisterFile/N24811 ) );
  AOI22_X1 U84057 ( .A1(n106026), .A2(n107312), .B1(n104789), .B2(n81265), 
        .ZN(n96556) );
  NOR2_X1 U84058 ( .A1(n96557), .A2(n96558), .ZN(n81557) );
  OR2_X1 U84059 ( .A1(n96559), .A2(n94999), .ZN(n96557) );
  AOI21_X1 U84060 ( .B1(n96560), .B2(n94258), .A(n96559), .ZN(n81556) );
  NOR2_X1 U84061 ( .A1(n81554), .A2(n105090), .ZN(n96559) );
  NAND2_X1 U84062 ( .A1(n105130), .A2(n94934), .ZN(n81554) );
  OAI21_X1 U84063 ( .B1(n106147), .B2(n96562), .A(n96563), .ZN(
        \DLX_Datapath/RegisterFile/N24810 ) );
  AOI22_X1 U84064 ( .A1(n96564), .A2(n70324), .B1(n104733), .B2(n94559), .ZN(
        n96563) );
  OAI21_X1 U84065 ( .B1(n105971), .B2(n96562), .A(n96566), .ZN(
        \DLX_Datapath/RegisterFile/N24809 ) );
  AOI22_X1 U84066 ( .A1(n96564), .A2(n70466), .B1(n96565), .B2(n94562), .ZN(
        n96566) );
  OAI21_X1 U84067 ( .B1(n106136), .B2(n96562), .A(n96567), .ZN(
        \DLX_Datapath/RegisterFile/N24808 ) );
  AOI22_X1 U84068 ( .A1(n96564), .A2(n69519), .B1(n104733), .B2(n94564), .ZN(
        n96567) );
  OAI21_X1 U84069 ( .B1(n106211), .B2(n96562), .A(n96568), .ZN(
        \DLX_Datapath/RegisterFile/N24807 ) );
  AOI22_X1 U84070 ( .A1(n96564), .A2(n70180), .B1(n96565), .B2(n94566), .ZN(
        n96568) );
  OAI21_X1 U84071 ( .B1(n106203), .B2(n96562), .A(n96569), .ZN(
        \DLX_Datapath/RegisterFile/N24806 ) );
  AOI22_X1 U84072 ( .A1(n96564), .A2(n74026), .B1(n104733), .B2(n94568), .ZN(
        n96569) );
  OAI21_X1 U84073 ( .B1(n106098), .B2(n96562), .A(n96570), .ZN(
        \DLX_Datapath/RegisterFile/N24805 ) );
  AOI22_X1 U84074 ( .A1(n96564), .A2(n70613), .B1(n96565), .B2(n94570), .ZN(
        n96570) );
  OAI21_X1 U84075 ( .B1(n106257), .B2(n105409), .A(n96571), .ZN(
        \DLX_Datapath/RegisterFile/N24804 ) );
  AOI22_X1 U84076 ( .A1(n96564), .A2(n74167), .B1(n104733), .B2(n94572), .ZN(
        n96571) );
  OAI21_X1 U84077 ( .B1(n105992), .B2(n105409), .A(n96572), .ZN(
        \DLX_Datapath/RegisterFile/N24803 ) );
  AOI22_X1 U84078 ( .A1(n96564), .A2(n74307), .B1(n96565), .B2(n94574), .ZN(
        n96572) );
  OAI21_X1 U84079 ( .B1(n106333), .B2(n105409), .A(n96573), .ZN(
        \DLX_Datapath/RegisterFile/N24802 ) );
  AOI22_X1 U84080 ( .A1(n96564), .A2(n73743), .B1(n96565), .B2(n94576), .ZN(
        n96573) );
  OAI21_X1 U84081 ( .B1(n106193), .B2(n105409), .A(n96574), .ZN(
        \DLX_Datapath/RegisterFile/N24801 ) );
  AOI22_X1 U84082 ( .A1(n96564), .A2(n73447), .B1(n104733), .B2(n94578), .ZN(
        n96574) );
  OAI21_X1 U84083 ( .B1(n106130), .B2(n105409), .A(n96575), .ZN(
        \DLX_Datapath/RegisterFile/N24800 ) );
  AOI22_X1 U84084 ( .A1(n96564), .A2(n73884), .B1(n96565), .B2(n94580), .ZN(
        n96575) );
  OAI21_X1 U84085 ( .B1(n106188), .B2(n105409), .A(n96576), .ZN(
        \DLX_Datapath/RegisterFile/N24799 ) );
  AOI22_X1 U84086 ( .A1(n96564), .A2(n73596), .B1(n104733), .B2(n94582), .ZN(
        n96576) );
  OAI21_X1 U84087 ( .B1(n106162), .B2(n105409), .A(n96577), .ZN(
        \DLX_Datapath/RegisterFile/N24798 ) );
  AOI22_X1 U84088 ( .A1(n96564), .A2(n73158), .B1(n96565), .B2(n94584), .ZN(
        n96577) );
  OAI21_X1 U84089 ( .B1(n106103), .B2(n105409), .A(n96578), .ZN(
        \DLX_Datapath/RegisterFile/N24797 ) );
  AOI22_X1 U84090 ( .A1(n96564), .A2(n73300), .B1(n104733), .B2(n94586), .ZN(
        n96578) );
  OAI21_X1 U84091 ( .B1(n106219), .B2(n105409), .A(n96579), .ZN(
        \DLX_Datapath/RegisterFile/N24796 ) );
  AOI22_X1 U84092 ( .A1(n96564), .A2(n73016), .B1(n104733), .B2(n94588), .ZN(
        n96579) );
  OAI21_X1 U84093 ( .B1(n106110), .B2(n105409), .A(n96580), .ZN(
        \DLX_Datapath/RegisterFile/N24795 ) );
  AOI22_X1 U84094 ( .A1(n96564), .A2(n72866), .B1(n96565), .B2(n94590), .ZN(
        n96580) );
  OAI21_X1 U84095 ( .B1(n106231), .B2(n105409), .A(n96581), .ZN(
        \DLX_Datapath/RegisterFile/N24794 ) );
  AOI22_X1 U84096 ( .A1(n96564), .A2(n70762), .B1(n104733), .B2(n94592), .ZN(
        n96581) );
  OAI21_X1 U84097 ( .B1(n106170), .B2(n105409), .A(n96582), .ZN(
        \DLX_Datapath/RegisterFile/N24793 ) );
  AOI22_X1 U84098 ( .A1(n96564), .A2(n70921), .B1(n96565), .B2(n94594), .ZN(
        n96582) );
  OAI21_X1 U84099 ( .B1(n81281), .B2(n105409), .A(n96583), .ZN(
        \DLX_Datapath/RegisterFile/N24792 ) );
  AOI22_X1 U84100 ( .A1(n96564), .A2(n71066), .B1(n96565), .B2(n94596), .ZN(
        n96583) );
  OAI21_X1 U84101 ( .B1(n106071), .B2(n105409), .A(n96584), .ZN(
        \DLX_Datapath/RegisterFile/N24791 ) );
  AOI22_X1 U84102 ( .A1(n96564), .A2(n70027), .B1(n104733), .B2(n94598), .ZN(
        n96584) );
  OAI21_X1 U84103 ( .B1(n106197), .B2(n105409), .A(n96585), .ZN(
        \DLX_Datapath/RegisterFile/N24790 ) );
  AOI22_X1 U84104 ( .A1(n96564), .A2(n72556), .B1(n96565), .B2(n94600), .ZN(
        n96585) );
  OAI21_X1 U84105 ( .B1(n81278), .B2(n105409), .A(n96586), .ZN(
        \DLX_Datapath/RegisterFile/N24789 ) );
  AOI22_X1 U84106 ( .A1(n96564), .A2(n71215), .B1(n104733), .B2(n94602), .ZN(
        n96586) );
  OAI21_X1 U84107 ( .B1(n106158), .B2(n105409), .A(n96587), .ZN(
        \DLX_Datapath/RegisterFile/N24788 ) );
  AOI22_X1 U84108 ( .A1(n96564), .A2(n72698), .B1(n104733), .B2(n94604), .ZN(
        n96587) );
  OAI21_X1 U84109 ( .B1(n106114), .B2(n105409), .A(n96588), .ZN(
        \DLX_Datapath/RegisterFile/N24787 ) );
  AOI22_X1 U84110 ( .A1(n96564), .A2(n72408), .B1(n96565), .B2(n94606), .ZN(
        n96588) );
  OAI21_X1 U84111 ( .B1(n106008), .B2(n105409), .A(n96589), .ZN(
        \DLX_Datapath/RegisterFile/N24786 ) );
  AOI22_X1 U84112 ( .A1(n96564), .A2(n71808), .B1(n104733), .B2(n94608), .ZN(
        n96589) );
  OAI21_X1 U84113 ( .B1(n106260), .B2(n105409), .A(n96590), .ZN(
        \DLX_Datapath/RegisterFile/N24785 ) );
  AOI22_X1 U84114 ( .A1(n96564), .A2(n72257), .B1(n104733), .B2(n94610), .ZN(
        n96590) );
  OAI21_X1 U84115 ( .B1(n81509), .B2(n105409), .A(n96591), .ZN(
        \DLX_Datapath/RegisterFile/N24784 ) );
  AOI22_X1 U84116 ( .A1(n96564), .A2(n72106), .B1(n96565), .B2(n94612), .ZN(
        n96591) );
  OAI21_X1 U84117 ( .B1(n81501), .B2(n105409), .A(n96592), .ZN(
        \DLX_Datapath/RegisterFile/N24783 ) );
  AOI22_X1 U84118 ( .A1(n96564), .A2(n71962), .B1(n104733), .B2(n94614), .ZN(
        n96592) );
  OAI21_X1 U84119 ( .B1(n106093), .B2(n105409), .A(n96593), .ZN(
        \DLX_Datapath/RegisterFile/N24782 ) );
  AOI22_X1 U84120 ( .A1(n96564), .A2(n71364), .B1(n96565), .B2(n94616), .ZN(
        n96593) );
  OAI21_X1 U84121 ( .B1(n106053), .B2(n105409), .A(n96594), .ZN(
        \DLX_Datapath/RegisterFile/N24781 ) );
  AOI22_X1 U84122 ( .A1(n96564), .A2(n71659), .B1(n96565), .B2(n94618), .ZN(
        n96594) );
  OAI21_X1 U84123 ( .B1(n105219), .B2(n105409), .A(n96595), .ZN(
        \DLX_Datapath/RegisterFile/N24780 ) );
  AOI22_X1 U84124 ( .A1(n96564), .A2(n71515), .B1(n96565), .B2(n94620), .ZN(
        n96595) );
  OAI21_X1 U84125 ( .B1(n106267), .B2(n105409), .A(n96596), .ZN(
        \DLX_Datapath/RegisterFile/N24779 ) );
  AOI22_X1 U84126 ( .A1(n96564), .A2(n69624), .B1(n104733), .B2(n94622), .ZN(
        n96596) );
  AND2_X2 U84127 ( .A1(n96597), .A2(n96598), .ZN(n96565) );
  AND2_X2 U84128 ( .A1(n96598), .A2(n96599), .ZN(n96564) );
  OR2_X1 U84129 ( .A1(n96562), .A2(n105089), .ZN(n96598) );
  NAND2_X1 U84130 ( .A1(n94296), .A2(n105130), .ZN(n96562) );
  OAI21_X1 U84131 ( .B1(n106147), .B2(n106006), .A(n96600), .ZN(
        \DLX_Datapath/RegisterFile/N24778 ) );
  AOI22_X1 U84132 ( .A1(n106004), .A2(n81521), .B1(n104943), .B2(n107877), 
        .ZN(n96600) );
  OAI21_X1 U84133 ( .B1(n81594), .B2(n81651), .A(n96601), .ZN(
        \DLX_Datapath/RegisterFile/N24777 ) );
  AOI22_X1 U84134 ( .A1(n81653), .A2(n106003), .B1(n104945), .B2(n107974), 
        .ZN(n96601) );
  OAI21_X1 U84135 ( .B1(n106136), .B2(n81594), .A(n96602), .ZN(
        \DLX_Datapath/RegisterFile/N24776 ) );
  AOI22_X1 U84136 ( .A1(n106003), .A2(n81380), .B1(n104942), .B2(n107238), 
        .ZN(n96602) );
  OAI21_X1 U84137 ( .B1(n106206), .B2(n106006), .A(n96603), .ZN(
        \DLX_Datapath/RegisterFile/N24774 ) );
  AOI22_X1 U84138 ( .A1(n106003), .A2(n81428), .B1(n104942), .B2(n110679), 
        .ZN(n96603) );
  OAI21_X1 U84139 ( .B1(n106098), .B2(n106006), .A(n96604), .ZN(
        \DLX_Datapath/RegisterFile/N24773 ) );
  AOI22_X1 U84140 ( .A1(n106003), .A2(n81410), .B1(n104945), .B2(n108079), 
        .ZN(n96604) );
  OAI21_X1 U84141 ( .B1(n106255), .B2(n106006), .A(n96605), .ZN(
        \DLX_Datapath/RegisterFile/N24772 ) );
  AOI22_X1 U84142 ( .A1(n81700), .A2(n106003), .B1(n104946), .B2(n110776), 
        .ZN(n96605) );
  OAI21_X1 U84143 ( .B1(n81594), .B2(n105990), .A(n96606), .ZN(
        \DLX_Datapath/RegisterFile/N24771 ) );
  AOI22_X1 U84144 ( .A1(n81632), .A2(n106003), .B1(n104944), .B2(n110877), 
        .ZN(n96606) );
  OAI21_X1 U84145 ( .B1(n106333), .B2(n106006), .A(n96607), .ZN(
        \DLX_Datapath/RegisterFile/N24770 ) );
  AOI22_X1 U84146 ( .A1(n106003), .A2(n81414), .B1(n73744), .B2(n104946), .ZN(
        n96607) );
  OAI21_X1 U84147 ( .B1(n106193), .B2(n106006), .A(n96608), .ZN(
        \DLX_Datapath/RegisterFile/N24769 ) );
  AOI22_X1 U84148 ( .A1(n106005), .A2(n81317), .B1(n73448), .B2(n104942), .ZN(
        n96608) );
  AOI22_X1 U84150 ( .A1(n106004), .A2(n81386), .B1(n73885), .B2(n104944), .ZN(
        n96609) );
  OAI21_X1 U84151 ( .B1(n106188), .B2(n106006), .A(n96610), .ZN(
        \DLX_Datapath/RegisterFile/N24767 ) );
  AOI22_X1 U84152 ( .A1(n106005), .A2(n81320), .B1(n73597), .B2(n104943), .ZN(
        n96610) );
  OAI21_X1 U84153 ( .B1(n106103), .B2(n106006), .A(n96611), .ZN(
        \DLX_Datapath/RegisterFile/N24765 ) );
  AOI22_X1 U84154 ( .A1(n106004), .A2(n81405), .B1(n73301), .B2(n104945), .ZN(
        n96611) );
  OAI21_X1 U84155 ( .B1(n106221), .B2(n106006), .A(n96612), .ZN(
        \DLX_Datapath/RegisterFile/N24764 ) );
  AOI22_X1 U84156 ( .A1(n106005), .A2(n81402), .B1(n73017), .B2(n104943), .ZN(
        n96612) );
  OAI21_X1 U84157 ( .B1(n81398), .B2(n106006), .A(n96613), .ZN(
        \DLX_Datapath/RegisterFile/N24763 ) );
  AOI22_X1 U84158 ( .A1(n106003), .A2(n81400), .B1(n104944), .B2(n109811), 
        .ZN(n96613) );
  OAI21_X1 U84159 ( .B1(n106071), .B2(n106006), .A(n96614), .ZN(
        \DLX_Datapath/RegisterFile/N24759 ) );
  AOI22_X1 U84160 ( .A1(n106005), .A2(n81506), .B1(n104946), .B2(n107657), 
        .ZN(n96614) );
  OAI21_X1 U84161 ( .B1(n106200), .B2(n106006), .A(n96615), .ZN(
        \DLX_Datapath/RegisterFile/N24758 ) );
  AOI22_X1 U84162 ( .A1(n106005), .A2(n81313), .B1(n104943), .B2(n109575), 
        .ZN(n96615) );
  OAI21_X1 U84163 ( .B1(n106008), .B2(n106006), .A(n96616), .ZN(
        \DLX_Datapath/RegisterFile/N24754 ) );
  AOI22_X1 U84164 ( .A1(n106005), .A2(n81590), .B1(n104943), .B2(n109001), 
        .ZN(n96616) );
  OAI21_X1 U84165 ( .B1(n81267), .B2(n106006), .A(n96617), .ZN(
        \DLX_Datapath/RegisterFile/N24753 ) );
  AOI22_X1 U84166 ( .A1(n106005), .A2(n81423), .B1(n104941), .B2(n109349), 
        .ZN(n96617) );
  OAI21_X1 U84167 ( .B1(n106045), .B2(n106006), .A(n96618), .ZN(
        \DLX_Datapath/RegisterFile/N24752 ) );
  AOI22_X1 U84168 ( .A1(n106004), .A2(n81511), .B1(n104942), .B2(n109231), 
        .ZN(n96618) );
  OAI21_X1 U84169 ( .B1(n106050), .B2(n106006), .A(n96619), .ZN(
        \DLX_Datapath/RegisterFile/N24751 ) );
  AOI22_X1 U84170 ( .A1(n106004), .A2(n81503), .B1(n104941), .B2(n109123), 
        .ZN(n96619) );
  OAI21_X1 U84171 ( .B1(n106054), .B2(n106006), .A(n96620), .ZN(
        \DLX_Datapath/RegisterFile/N24749 ) );
  AOI22_X1 U84172 ( .A1(n106004), .A2(n81500), .B1(n104942), .B2(n108885), 
        .ZN(n96620) );
  OAI21_X1 U84173 ( .B1(n106267), .B2(n106006), .A(n96621), .ZN(
        \DLX_Datapath/RegisterFile/N24747 ) );
  AOI22_X1 U84174 ( .A1(n106004), .A2(n81327), .B1(n104943), .B2(n107313), 
        .ZN(n96621) );
  AND2_X2 U84175 ( .A1(n96599), .A2(n96622), .ZN(n81597) );
  AND2_X2 U84176 ( .A1(n96597), .A2(n96622), .ZN(n81596) );
  OR2_X1 U84177 ( .A1(n81594), .A2(n105089), .ZN(n96622) );
  NAND2_X1 U84178 ( .A1(n105129), .A2(n94331), .ZN(n81594) );
  OAI21_X1 U84179 ( .B1(n106147), .B2(n105408), .A(n96624), .ZN(
        \DLX_Datapath/RegisterFile/N24746 ) );
  AOI22_X1 U84180 ( .A1(n96625), .A2(n94667), .B1(n96626), .B2(n70326), .ZN(
        n96624) );
  OAI21_X1 U84181 ( .B1(n105971), .B2(n105408), .A(n96627), .ZN(
        \DLX_Datapath/RegisterFile/N24745 ) );
  AOI22_X1 U84182 ( .A1(n96625), .A2(n94670), .B1(n96626), .B2(n70468), .ZN(
        n96627) );
  OAI21_X1 U84183 ( .B1(n106136), .B2(n105408), .A(n96628), .ZN(
        \DLX_Datapath/RegisterFile/N24744 ) );
  AOI22_X1 U84184 ( .A1(n96625), .A2(n94672), .B1(n96626), .B2(n69521), .ZN(
        n96628) );
  OAI21_X1 U84185 ( .B1(n81299), .B2(n105408), .A(n96629), .ZN(
        \DLX_Datapath/RegisterFile/N24743 ) );
  AOI22_X1 U84186 ( .A1(n96625), .A2(n94674), .B1(n96626), .B2(n70182), .ZN(
        n96629) );
  OAI21_X1 U84187 ( .B1(n81306), .B2(n105408), .A(n96630), .ZN(
        \DLX_Datapath/RegisterFile/N24742 ) );
  AOI22_X1 U84188 ( .A1(n96625), .A2(n94676), .B1(n96626), .B2(n74028), .ZN(
        n96630) );
  OAI21_X1 U84189 ( .B1(n106098), .B2(n105408), .A(n96631), .ZN(
        \DLX_Datapath/RegisterFile/N24741 ) );
  AOI22_X1 U84190 ( .A1(n96625), .A2(n94678), .B1(n96626), .B2(n70615), .ZN(
        n96631) );
  OAI21_X1 U84191 ( .B1(n81270), .B2(n105408), .A(n96632), .ZN(
        \DLX_Datapath/RegisterFile/N24740 ) );
  AOI22_X1 U84192 ( .A1(n96625), .A2(n94680), .B1(n96626), .B2(n74169), .ZN(
        n96632) );
  OAI21_X1 U84193 ( .B1(n105992), .B2(n105408), .A(n96633), .ZN(
        \DLX_Datapath/RegisterFile/N24739 ) );
  AOI22_X1 U84194 ( .A1(n96625), .A2(n94682), .B1(n96626), .B2(n74309), .ZN(
        n96633) );
  OAI21_X1 U84195 ( .B1(n106333), .B2(n105408), .A(n96634), .ZN(
        \DLX_Datapath/RegisterFile/N24738 ) );
  AOI22_X1 U84196 ( .A1(n96625), .A2(n94684), .B1(n96626), .B2(n73745), .ZN(
        n96634) );
  OAI21_X1 U84197 ( .B1(n81315), .B2(n105408), .A(n96635), .ZN(
        \DLX_Datapath/RegisterFile/N24737 ) );
  AOI22_X1 U84198 ( .A1(n96625), .A2(n94686), .B1(n96626), .B2(n73449), .ZN(
        n96635) );
  OAI21_X1 U84199 ( .B1(n106129), .B2(n105408), .A(n96636), .ZN(
        \DLX_Datapath/RegisterFile/N24736 ) );
  AOI22_X1 U84200 ( .A1(n96625), .A2(n94688), .B1(n96626), .B2(n73886), .ZN(
        n96636) );
  OAI21_X1 U84201 ( .B1(n81318), .B2(n105408), .A(n96637), .ZN(
        \DLX_Datapath/RegisterFile/N24735 ) );
  AOI22_X1 U84202 ( .A1(n96625), .A2(n94690), .B1(n96626), .B2(n73598), .ZN(
        n96637) );
  OAI21_X1 U84203 ( .B1(n106162), .B2(n105408), .A(n96638), .ZN(
        \DLX_Datapath/RegisterFile/N24734 ) );
  AOI22_X1 U84204 ( .A1(n96625), .A2(n94692), .B1(n96626), .B2(n73160), .ZN(
        n96638) );
  OAI21_X1 U84205 ( .B1(n106103), .B2(n105408), .A(n96639), .ZN(
        \DLX_Datapath/RegisterFile/N24733 ) );
  AOI22_X1 U84206 ( .A1(n96625), .A2(n94694), .B1(n96626), .B2(n73302), .ZN(
        n96639) );
  OAI21_X1 U84207 ( .B1(n106221), .B2(n105408), .A(n96640), .ZN(
        \DLX_Datapath/RegisterFile/N24732 ) );
  AOI22_X1 U84208 ( .A1(n96625), .A2(n94696), .B1(n96626), .B2(n73018), .ZN(
        n96640) );
  OAI21_X1 U84209 ( .B1(n106111), .B2(n105408), .A(n96641), .ZN(
        \DLX_Datapath/RegisterFile/N24731 ) );
  AOI22_X1 U84210 ( .A1(n96625), .A2(n94698), .B1(n96626), .B2(n72868), .ZN(
        n96641) );
  OAI21_X1 U84211 ( .B1(n106231), .B2(n105408), .A(n96642), .ZN(
        \DLX_Datapath/RegisterFile/N24730 ) );
  AOI22_X1 U84212 ( .A1(n96625), .A2(n94700), .B1(n96626), .B2(n70764), .ZN(
        n96642) );
  OAI21_X1 U84213 ( .B1(n106170), .B2(n105408), .A(n96643), .ZN(
        \DLX_Datapath/RegisterFile/N24729 ) );
  AOI22_X1 U84214 ( .A1(n96625), .A2(n94702), .B1(n96626), .B2(n70923), .ZN(
        n96643) );
  OAI21_X1 U84215 ( .B1(n81281), .B2(n105408), .A(n96644), .ZN(
        \DLX_Datapath/RegisterFile/N24728 ) );
  AOI22_X1 U84216 ( .A1(n96625), .A2(n94704), .B1(n96626), .B2(n71068), .ZN(
        n96644) );
  OAI21_X1 U84217 ( .B1(n106071), .B2(n105408), .A(n96645), .ZN(
        \DLX_Datapath/RegisterFile/N24727 ) );
  AOI22_X1 U84218 ( .A1(n96625), .A2(n94706), .B1(n96626), .B2(n70029), .ZN(
        n96645) );
  OAI21_X1 U84219 ( .B1(n81310), .B2(n105408), .A(n96646), .ZN(
        \DLX_Datapath/RegisterFile/N24726 ) );
  AOI22_X1 U84220 ( .A1(n96625), .A2(n94708), .B1(n96626), .B2(n72558), .ZN(
        n96646) );
  OAI21_X1 U84221 ( .B1(n81278), .B2(n105408), .A(n96647), .ZN(
        \DLX_Datapath/RegisterFile/N24725 ) );
  AOI22_X1 U84222 ( .A1(n96625), .A2(n94710), .B1(n96626), .B2(n71217), .ZN(
        n96647) );
  OAI21_X1 U84223 ( .B1(n106158), .B2(n105408), .A(n96648), .ZN(
        \DLX_Datapath/RegisterFile/N24724 ) );
  AOI22_X1 U84224 ( .A1(n96625), .A2(n94712), .B1(n96626), .B2(n72700), .ZN(
        n96648) );
  OAI21_X1 U84225 ( .B1(n106114), .B2(n105408), .A(n96649), .ZN(
        \DLX_Datapath/RegisterFile/N24723 ) );
  AOI22_X1 U84226 ( .A1(n96625), .A2(n94714), .B1(n96626), .B2(n72410), .ZN(
        n96649) );
  OAI21_X1 U84227 ( .B1(n106008), .B2(n105408), .A(n96650), .ZN(
        \DLX_Datapath/RegisterFile/N24722 ) );
  AOI22_X1 U84228 ( .A1(n96625), .A2(n81259), .B1(n96626), .B2(n71810), .ZN(
        n96650) );
  OAI21_X1 U84229 ( .B1(n106261), .B2(n105408), .A(n96651), .ZN(
        \DLX_Datapath/RegisterFile/N24721 ) );
  AOI22_X1 U84230 ( .A1(n96625), .A2(n94717), .B1(n96626), .B2(n72259), .ZN(
        n96651) );
  OAI21_X1 U84231 ( .B1(n106046), .B2(n105408), .A(n96652), .ZN(
        \DLX_Datapath/RegisterFile/N24720 ) );
  AOI22_X1 U84232 ( .A1(n96625), .A2(n94719), .B1(n96626), .B2(n72108), .ZN(
        n96652) );
  OAI21_X1 U84233 ( .B1(n81501), .B2(n105408), .A(n96653), .ZN(
        \DLX_Datapath/RegisterFile/N24719 ) );
  AOI22_X1 U84234 ( .A1(n96625), .A2(n94721), .B1(n96626), .B2(n71964), .ZN(
        n96653) );
  OAI21_X1 U84235 ( .B1(n106093), .B2(n105408), .A(n96654), .ZN(
        \DLX_Datapath/RegisterFile/N24718 ) );
  AOI22_X1 U84236 ( .A1(n96625), .A2(n94723), .B1(n96626), .B2(n71366), .ZN(
        n96654) );
  OAI21_X1 U84237 ( .B1(n106054), .B2(n105408), .A(n96655), .ZN(
        \DLX_Datapath/RegisterFile/N24717 ) );
  AOI22_X1 U84238 ( .A1(n96625), .A2(n94725), .B1(n96626), .B2(n71661), .ZN(
        n96655) );
  OAI21_X1 U84239 ( .B1(n105218), .B2(n105408), .A(n96656), .ZN(
        \DLX_Datapath/RegisterFile/N24716 ) );
  AOI22_X1 U84240 ( .A1(n96625), .A2(n94727), .B1(n96626), .B2(n71517), .ZN(
        n96656) );
  OAI21_X1 U84241 ( .B1(n81262), .B2(n105408), .A(n96657), .ZN(
        \DLX_Datapath/RegisterFile/N24715 ) );
  AOI22_X1 U84242 ( .A1(n96625), .A2(n94729), .B1(n96626), .B2(n69626), .ZN(
        n96657) );
  AND2_X2 U84243 ( .A1(n96599), .A2(n96658), .ZN(n96626) );
  OAI21_X1 U84244 ( .B1(n94366), .B2(n96597), .A(n105602), .ZN(n96599) );
  AND2_X2 U84245 ( .A1(n96597), .A2(n96658), .ZN(n96625) );
  OR2_X1 U84246 ( .A1(n96623), .A2(n105091), .ZN(n96658) );
  NOR2_X1 U84247 ( .A1(n96558), .A2(n94999), .ZN(n96597) );
  NAND2_X1 U84248 ( .A1(n94367), .A2(n105129), .ZN(n96623) );
  OAI21_X1 U84249 ( .B1(n106025), .B2(n81651), .A(n96659), .ZN(
        \DLX_Datapath/RegisterFile/N24713 ) );
  AOI22_X1 U84250 ( .A1(n106024), .A2(n107975), .B1(n94511), .B2(n106017), 
        .ZN(n96659) );
  OAI21_X1 U84251 ( .B1(n106137), .B2(n106025), .A(n96660), .ZN(
        \DLX_Datapath/RegisterFile/N24712 ) );
  AOI22_X1 U84252 ( .A1(n106023), .A2(n107239), .B1(n81568), .B2(n81539), .ZN(
        n96660) );
  OAI21_X1 U84253 ( .B1(n106098), .B2(n106025), .A(n96661), .ZN(
        \DLX_Datapath/RegisterFile/N24709 ) );
  AOI22_X1 U84254 ( .A1(n106023), .A2(n108080), .B1(n94516), .B2(n106017), 
        .ZN(n96661) );
  OAI21_X1 U84255 ( .B1(n106025), .B2(n105992), .A(n96662), .ZN(
        \DLX_Datapath/RegisterFile/N24707 ) );
  AOI22_X1 U84256 ( .A1(n106023), .A2(n110878), .B1(n94519), .B2(n106017), 
        .ZN(n96662) );
  OAI21_X1 U84257 ( .B1(n106333), .B2(n106025), .A(n96663), .ZN(
        \DLX_Datapath/RegisterFile/N24706 ) );
  AOI22_X1 U84258 ( .A1(n106023), .A2(n110472), .B1(n81568), .B2(n80192), .ZN(
        n96663) );
  OAI21_X1 U84259 ( .B1(n106129), .B2(n106025), .A(n96664), .ZN(
        \DLX_Datapath/RegisterFile/N24704 ) );
  AOI22_X1 U84260 ( .A1(n106023), .A2(n110571), .B1(n94523), .B2(n106017), 
        .ZN(n96664) );
  OAI21_X1 U84261 ( .B1(n106104), .B2(n106025), .A(n96665), .ZN(
        \DLX_Datapath/RegisterFile/N24701 ) );
  AOI22_X1 U84262 ( .A1(n106023), .A2(n110145), .B1(n94527), .B2(n106017), 
        .ZN(n96665) );
  OAI21_X1 U84263 ( .B1(n106219), .B2(n106025), .A(n96666), .ZN(
        \DLX_Datapath/RegisterFile/N24700 ) );
  AOI22_X1 U84264 ( .A1(n106023), .A2(n109929), .B1(n81568), .B2(n81297), .ZN(
        n96666) );
  OAI21_X1 U84265 ( .B1(n81398), .B2(n106025), .A(n96667), .ZN(
        \DLX_Datapath/RegisterFile/N24699 ) );
  AOI22_X1 U84266 ( .A1(n106024), .A2(n109812), .B1(n94530), .B2(n106017), 
        .ZN(n96667) );
  OAI21_X1 U84267 ( .B1(n106170), .B2(n106025), .A(n96668), .ZN(
        \DLX_Datapath/RegisterFile/N24697 ) );
  AOI22_X1 U84268 ( .A1(n106022), .A2(n108309), .B1(n81568), .B2(n106168), 
        .ZN(n96668) );
  OAI21_X1 U84269 ( .B1(n106235), .B2(n81564), .A(n96669), .ZN(
        \DLX_Datapath/RegisterFile/N24696 ) );
  AOI22_X1 U84270 ( .A1(n106024), .A2(n108420), .B1(n106018), .B2(n81283), 
        .ZN(n96669) );
  OAI21_X1 U84271 ( .B1(n106071), .B2(n81564), .A(n96670), .ZN(
        \DLX_Datapath/RegisterFile/N24695 ) );
  AOI22_X1 U84272 ( .A1(n106022), .A2(n107658), .B1(n81568), .B2(n81453), .ZN(
        n96670) );
  OAI21_X1 U84273 ( .B1(n106197), .B2(n81564), .A(n96671), .ZN(
        \DLX_Datapath/RegisterFile/N24694 ) );
  AOI22_X1 U84274 ( .A1(n106024), .A2(n109576), .B1(n94536), .B2(n106017), 
        .ZN(n96671) );
  OAI21_X1 U84275 ( .B1(n81588), .B2(n106025), .A(n96672), .ZN(
        \DLX_Datapath/RegisterFile/N24690 ) );
  AOI22_X1 U84276 ( .A1(n106022), .A2(n109002), .B1(n94541), .B2(n106017), 
        .ZN(n96672) );
  OAI21_X1 U84277 ( .B1(n106259), .B2(n81564), .A(n96673), .ZN(
        \DLX_Datapath/RegisterFile/N24689 ) );
  AOI22_X1 U84278 ( .A1(n106024), .A2(n109350), .B1(n81568), .B2(n81269), .ZN(
        n96673) );
  OAI21_X1 U84279 ( .B1(n106043), .B2(n81564), .A(n96674), .ZN(
        \DLX_Datapath/RegisterFile/N24688 ) );
  AOI22_X1 U84280 ( .A1(n106022), .A2(n109232), .B1(n105624), .B2(n106017), 
        .ZN(n96674) );
  OAI21_X1 U84281 ( .B1(n106048), .B2(n81564), .A(n96675), .ZN(
        \DLX_Datapath/RegisterFile/N24687 ) );
  AOI22_X1 U84282 ( .A1(n106024), .A2(n109124), .B1(n94546), .B2(n106017), 
        .ZN(n96675) );
  OAI21_X1 U84283 ( .B1(n106093), .B2(n106025), .A(n96676), .ZN(
        \DLX_Datapath/RegisterFile/N24686 ) );
  AOI22_X1 U84284 ( .A1(n106022), .A2(n108659), .B1(n94548), .B2(n106017), 
        .ZN(n96676) );
  OAI21_X1 U84285 ( .B1(n106054), .B2(n106025), .A(n96677), .ZN(
        \DLX_Datapath/RegisterFile/N24685 ) );
  AOI22_X1 U84286 ( .A1(n106024), .A2(n108886), .B1(n81783), .B2(n106017), 
        .ZN(n96677) );
  OAI21_X1 U84287 ( .B1(n106269), .B2(n106025), .A(n96678), .ZN(
        \DLX_Datapath/RegisterFile/N24683 ) );
  AOI22_X1 U84288 ( .A1(n106022), .A2(n107314), .B1(n106018), .B2(n81265), 
        .ZN(n96678) );
  NOR2_X1 U84289 ( .A1(n96679), .A2(n104690), .ZN(n81568) );
  AOI21_X1 U84290 ( .B1(n96560), .B2(n94398), .A(n96680), .ZN(n81566) );
  NOR2_X1 U84291 ( .A1(n81564), .A2(n105094), .ZN(n96680) );
  NAND2_X1 U84292 ( .A1(n105130), .A2(n94399), .ZN(n81564) );
  OAI21_X1 U84293 ( .B1(n106147), .B2(n105407), .A(n96682), .ZN(
        \DLX_Datapath/RegisterFile/N24682 ) );
  AOI22_X1 U84294 ( .A1(n105406), .A2(n107879), .B1(n105404), .B2(n94559), 
        .ZN(n96682) );
  OAI21_X1 U84295 ( .B1(n105971), .B2(n105407), .A(n96685), .ZN(
        \DLX_Datapath/RegisterFile/N24681 ) );
  AOI22_X1 U84296 ( .A1(n105406), .A2(n70470), .B1(n105403), .B2(n94562), .ZN(
        n96685) );
  OAI21_X1 U84297 ( .B1(n106138), .B2(n96681), .A(n96686), .ZN(
        \DLX_Datapath/RegisterFile/N24680 ) );
  AOI22_X1 U84298 ( .A1(n105406), .A2(n107240), .B1(n105404), .B2(n94564), 
        .ZN(n96686) );
  OAI21_X1 U84299 ( .B1(n106211), .B2(n96681), .A(n96687), .ZN(
        \DLX_Datapath/RegisterFile/N24679 ) );
  AOI22_X1 U84300 ( .A1(n105406), .A2(n107779), .B1(n105403), .B2(n94566), 
        .ZN(n96687) );
  OAI21_X1 U84301 ( .B1(n106206), .B2(n96681), .A(n96688), .ZN(
        \DLX_Datapath/RegisterFile/N24678 ) );
  AOI22_X1 U84302 ( .A1(n105406), .A2(n110681), .B1(n105404), .B2(n94568), 
        .ZN(n96688) );
  OAI21_X1 U84303 ( .B1(n106099), .B2(n96681), .A(n96689), .ZN(
        \DLX_Datapath/RegisterFile/N24677 ) );
  AOI22_X1 U84304 ( .A1(n105406), .A2(n108081), .B1(n105403), .B2(n94570), 
        .ZN(n96689) );
  OAI21_X1 U84305 ( .B1(n106254), .B2(n96681), .A(n96690), .ZN(
        \DLX_Datapath/RegisterFile/N24676 ) );
  AOI22_X1 U84306 ( .A1(n105406), .A2(n110778), .B1(n105404), .B2(n94572), 
        .ZN(n96690) );
  OAI21_X1 U84307 ( .B1(n105992), .B2(n105407), .A(n96691), .ZN(
        \DLX_Datapath/RegisterFile/N24675 ) );
  AOI22_X1 U84308 ( .A1(n105406), .A2(n110879), .B1(n105403), .B2(n94574), 
        .ZN(n96691) );
  OAI21_X1 U84309 ( .B1(n106333), .B2(n96681), .A(n96692), .ZN(
        \DLX_Datapath/RegisterFile/N24674 ) );
  AOI22_X1 U84310 ( .A1(n105405), .A2(n110473), .B1(n105403), .B2(n94576), 
        .ZN(n96692) );
  OAI21_X1 U84311 ( .B1(n106192), .B2(n105407), .A(n96693), .ZN(
        \DLX_Datapath/RegisterFile/N24673 ) );
  AOI22_X1 U84312 ( .A1(n96683), .A2(n110255), .B1(n105402), .B2(n94578), .ZN(
        n96693) );
  OAI21_X1 U84313 ( .B1(n106129), .B2(n105407), .A(n96694), .ZN(
        \DLX_Datapath/RegisterFile/N24672 ) );
  AOI22_X1 U84314 ( .A1(n105406), .A2(n110572), .B1(n105402), .B2(n94580), 
        .ZN(n96694) );
  OAI21_X1 U84315 ( .B1(n81318), .B2(n105407), .A(n96695), .ZN(
        \DLX_Datapath/RegisterFile/N24671 ) );
  AOI22_X1 U84316 ( .A1(n105406), .A2(n110363), .B1(n105402), .B2(n94582), 
        .ZN(n96695) );
  OAI21_X1 U84317 ( .B1(n106162), .B2(n105407), .A(n96696), .ZN(
        \DLX_Datapath/RegisterFile/N24670 ) );
  AOI22_X1 U84318 ( .A1(n96683), .A2(n110039), .B1(n105402), .B2(n94584), .ZN(
        n96696) );
  OAI21_X1 U84319 ( .B1(n106104), .B2(n105407), .A(n96697), .ZN(
        \DLX_Datapath/RegisterFile/N24669 ) );
  AOI22_X1 U84320 ( .A1(n96683), .A2(n110146), .B1(n105402), .B2(n94586), .ZN(
        n96697) );
  OAI21_X1 U84321 ( .B1(n106218), .B2(n105407), .A(n96698), .ZN(
        \DLX_Datapath/RegisterFile/N24668 ) );
  AOI22_X1 U84322 ( .A1(n105406), .A2(n109930), .B1(n105402), .B2(n94588), 
        .ZN(n96698) );
  OAI21_X1 U84323 ( .B1(n106109), .B2(n105407), .A(n96699), .ZN(
        \DLX_Datapath/RegisterFile/N24667 ) );
  AOI22_X1 U84324 ( .A1(n96683), .A2(n109813), .B1(n105402), .B2(n94590), .ZN(
        n96699) );
  OAI21_X1 U84325 ( .B1(n106231), .B2(n105407), .A(n96700), .ZN(
        \DLX_Datapath/RegisterFile/N24666 ) );
  AOI22_X1 U84326 ( .A1(n105406), .A2(n108187), .B1(n105402), .B2(n94592), 
        .ZN(n96700) );
  OAI21_X1 U84327 ( .B1(n106170), .B2(n105407), .A(n96701), .ZN(
        \DLX_Datapath/RegisterFile/N24665 ) );
  AOI22_X1 U84328 ( .A1(n96683), .A2(n108310), .B1(n105402), .B2(n94594), .ZN(
        n96701) );
  OAI21_X1 U84329 ( .B1(n106237), .B2(n105407), .A(n96702), .ZN(
        \DLX_Datapath/RegisterFile/N24664 ) );
  AOI22_X1 U84330 ( .A1(n105406), .A2(n108421), .B1(n105402), .B2(n94596), 
        .ZN(n96702) );
  OAI21_X1 U84331 ( .B1(n106071), .B2(n105407), .A(n96703), .ZN(
        \DLX_Datapath/RegisterFile/N24663 ) );
  AOI22_X1 U84332 ( .A1(n96683), .A2(n107659), .B1(n105402), .B2(n94598), .ZN(
        n96703) );
  OAI21_X1 U84333 ( .B1(n106198), .B2(n105407), .A(n96704), .ZN(
        \DLX_Datapath/RegisterFile/N24662 ) );
  AOI22_X1 U84334 ( .A1(n105405), .A2(n109577), .B1(n105403), .B2(n94600), 
        .ZN(n96704) );
  OAI21_X1 U84335 ( .B1(n81278), .B2(n105407), .A(n96705), .ZN(
        \DLX_Datapath/RegisterFile/N24661 ) );
  AOI22_X1 U84336 ( .A1(n105405), .A2(n108538), .B1(n105404), .B2(n94602), 
        .ZN(n96705) );
  OAI21_X1 U84337 ( .B1(n106158), .B2(n105407), .A(n96706), .ZN(
        \DLX_Datapath/RegisterFile/N24660 ) );
  AOI22_X1 U84338 ( .A1(n105405), .A2(n109682), .B1(n105403), .B2(n94604), 
        .ZN(n96706) );
  OAI21_X1 U84339 ( .B1(n106114), .B2(n105407), .A(n96707), .ZN(
        \DLX_Datapath/RegisterFile/N24659 ) );
  AOI22_X1 U84340 ( .A1(n105405), .A2(n109466), .B1(n105404), .B2(n94606), 
        .ZN(n96707) );
  OAI21_X1 U84341 ( .B1(n81588), .B2(n105407), .A(n96708), .ZN(
        \DLX_Datapath/RegisterFile/N24658 ) );
  AOI22_X1 U84342 ( .A1(n105405), .A2(n109003), .B1(n105403), .B2(n94608), 
        .ZN(n96708) );
  OAI21_X1 U84343 ( .B1(n81267), .B2(n105407), .A(n96709), .ZN(
        \DLX_Datapath/RegisterFile/N24657 ) );
  AOI22_X1 U84344 ( .A1(n105405), .A2(n109351), .B1(n105404), .B2(n94610), 
        .ZN(n96709) );
  OAI21_X1 U84345 ( .B1(n106045), .B2(n105407), .A(n96710), .ZN(
        \DLX_Datapath/RegisterFile/N24656 ) );
  AOI22_X1 U84346 ( .A1(n105405), .A2(n109233), .B1(n105403), .B2(n94612), 
        .ZN(n96710) );
  OAI21_X1 U84347 ( .B1(n81501), .B2(n105407), .A(n96711), .ZN(
        \DLX_Datapath/RegisterFile/N24655 ) );
  AOI22_X1 U84348 ( .A1(n105405), .A2(n109125), .B1(n105404), .B2(n94614), 
        .ZN(n96711) );
  OAI21_X1 U84349 ( .B1(n106093), .B2(n105407), .A(n96712), .ZN(
        \DLX_Datapath/RegisterFile/N24654 ) );
  AOI22_X1 U84350 ( .A1(n105405), .A2(n108660), .B1(n105403), .B2(n94616), 
        .ZN(n96712) );
  OAI21_X1 U84351 ( .B1(n106054), .B2(n105407), .A(n96713), .ZN(
        \DLX_Datapath/RegisterFile/N24653 ) );
  AOI22_X1 U84352 ( .A1(n105405), .A2(n108887), .B1(n105404), .B2(n94618), 
        .ZN(n96713) );
  OAI21_X1 U84353 ( .B1(n105218), .B2(n105407), .A(n96714), .ZN(
        \DLX_Datapath/RegisterFile/N24652 ) );
  AOI22_X1 U84354 ( .A1(n105405), .A2(n108775), .B1(n105404), .B2(n94620), 
        .ZN(n96714) );
  OAI21_X1 U84355 ( .B1(n81262), .B2(n105407), .A(n96715), .ZN(
        \DLX_Datapath/RegisterFile/N24651 ) );
  AOI22_X1 U84356 ( .A1(n105405), .A2(n107315), .B1(n105403), .B2(n94622), 
        .ZN(n96715) );
  NOR2_X1 U84357 ( .A1(n96679), .A2(n96716), .ZN(n96684) );
  NOR2_X1 U84358 ( .A1(n96716), .A2(n96717), .ZN(n96683) );
  NOR2_X1 U84359 ( .A1(n96681), .A2(n105090), .ZN(n96716) );
  NAND2_X1 U84360 ( .A1(n94434), .A2(n105130), .ZN(n96681) );
  OAI21_X1 U84361 ( .B1(n106147), .B2(n106015), .A(n96718), .ZN(
        \DLX_Datapath/RegisterFile/N24650 ) );
  AOI22_X1 U84362 ( .A1(n104855), .A2(n81521), .B1(n70329), .B2(n81583), .ZN(
        n96718) );
  OAI21_X1 U84363 ( .B1(n106015), .B2(n81651), .A(n96719), .ZN(
        \DLX_Datapath/RegisterFile/N24649 ) );
  AOI22_X1 U84364 ( .A1(n81653), .A2(n104854), .B1(n70471), .B2(n106014), .ZN(
        n96719) );
  OAI21_X1 U84365 ( .B1(n106135), .B2(n106015), .A(n96720), .ZN(
        \DLX_Datapath/RegisterFile/N24648 ) );
  AOI22_X1 U84366 ( .A1(n104855), .A2(n81380), .B1(n69524), .B2(n106013), .ZN(
        n96720) );
  OAI21_X1 U84367 ( .B1(n106211), .B2(n106015), .A(n96721), .ZN(
        \DLX_Datapath/RegisterFile/N24647 ) );
  AOI22_X1 U84368 ( .A1(n104855), .A2(n81377), .B1(n70185), .B2(n106013), .ZN(
        n96721) );
  OAI21_X1 U84369 ( .B1(n106206), .B2(n106015), .A(n96722), .ZN(
        \DLX_Datapath/RegisterFile/N24646 ) );
  AOI22_X1 U84370 ( .A1(n104855), .A2(n81428), .B1(n74031), .B2(n106013), .ZN(
        n96722) );
  OAI21_X1 U84371 ( .B1(n106099), .B2(n106015), .A(n96723), .ZN(
        \DLX_Datapath/RegisterFile/N24645 ) );
  AOI22_X1 U84372 ( .A1(n104854), .A2(n81410), .B1(n70618), .B2(n106013), .ZN(
        n96723) );
  OAI21_X1 U84373 ( .B1(n106254), .B2(n106015), .A(n96724), .ZN(
        \DLX_Datapath/RegisterFile/N24644 ) );
  AOI22_X1 U84374 ( .A1(n81700), .A2(n104855), .B1(n74172), .B2(n106014), .ZN(
        n96724) );
  OAI21_X1 U84375 ( .B1(n106016), .B2(n105990), .A(n96725), .ZN(
        \DLX_Datapath/RegisterFile/N24643 ) );
  AOI22_X1 U84376 ( .A1(n81632), .A2(n104855), .B1(n74312), .B2(n106013), .ZN(
        n96725) );
  OAI21_X1 U84377 ( .B1(n106333), .B2(n106015), .A(n96726), .ZN(
        \DLX_Datapath/RegisterFile/N24642 ) );
  AOI22_X1 U84378 ( .A1(n104854), .A2(n81414), .B1(n73748), .B2(n106013), .ZN(
        n96726) );
  OAI21_X1 U84379 ( .B1(n106190), .B2(n106015), .A(n96727), .ZN(
        \DLX_Datapath/RegisterFile/N24641 ) );
  AOI22_X1 U84380 ( .A1(n81582), .A2(n81317), .B1(n73452), .B2(n106013), .ZN(
        n96727) );
  OAI21_X1 U84381 ( .B1(n106129), .B2(n106015), .A(n96728), .ZN(
        \DLX_Datapath/RegisterFile/N24640 ) );
  AOI22_X1 U84382 ( .A1(n104854), .A2(n81386), .B1(n73889), .B2(n106013), .ZN(
        n96728) );
  OAI21_X1 U84383 ( .B1(n106185), .B2(n106015), .A(n96729), .ZN(
        \DLX_Datapath/RegisterFile/N24639 ) );
  AOI22_X1 U84384 ( .A1(n81582), .A2(n81320), .B1(n73601), .B2(n106013), .ZN(
        n96729) );
  OAI21_X1 U84385 ( .B1(n106162), .B2(n106015), .A(n96730), .ZN(
        \DLX_Datapath/RegisterFile/N24638 ) );
  AOI22_X1 U84386 ( .A1(n81604), .A2(n104854), .B1(n73163), .B2(n81583), .ZN(
        n96730) );
  OAI21_X1 U84387 ( .B1(n106104), .B2(n106016), .A(n96731), .ZN(
        \DLX_Datapath/RegisterFile/N24637 ) );
  AOI22_X1 U84388 ( .A1(n104854), .A2(n81405), .B1(n73305), .B2(n81583), .ZN(
        n96731) );
  OAI21_X1 U84389 ( .B1(n106220), .B2(n106016), .A(n96732), .ZN(
        \DLX_Datapath/RegisterFile/N24636 ) );
  AOI22_X1 U84390 ( .A1(n104854), .A2(n81402), .B1(n73021), .B2(n106014), .ZN(
        n96732) );
  OAI21_X1 U84391 ( .B1(n106109), .B2(n106016), .A(n96733), .ZN(
        \DLX_Datapath/RegisterFile/N24635 ) );
  AOI22_X1 U84392 ( .A1(n104854), .A2(n81400), .B1(n72871), .B2(n81583), .ZN(
        n96733) );
  OAI21_X1 U84393 ( .B1(n106237), .B2(n106016), .A(n96734), .ZN(
        \DLX_Datapath/RegisterFile/N24632 ) );
  AOI22_X1 U84394 ( .A1(n104854), .A2(n81322), .B1(n71071), .B2(n106014), .ZN(
        n96734) );
  OAI21_X1 U84395 ( .B1(n106071), .B2(n106016), .A(n96735), .ZN(
        \DLX_Datapath/RegisterFile/N24631 ) );
  AOI22_X1 U84396 ( .A1(n81582), .A2(n81506), .B1(n70032), .B2(n81583), .ZN(
        n96735) );
  OAI21_X1 U84397 ( .B1(n106199), .B2(n106016), .A(n96736), .ZN(
        \DLX_Datapath/RegisterFile/N24630 ) );
  AOI22_X1 U84398 ( .A1(n81582), .A2(n81313), .B1(n72561), .B2(n106014), .ZN(
        n96736) );
  OAI21_X1 U84399 ( .B1(n106158), .B2(n106016), .A(n96737), .ZN(
        \DLX_Datapath/RegisterFile/N24628 ) );
  AOI22_X1 U84400 ( .A1(n81582), .A2(n81425), .B1(n72703), .B2(n81583), .ZN(
        n96737) );
  OAI21_X1 U84401 ( .B1(n106262), .B2(n106016), .A(n96738), .ZN(
        \DLX_Datapath/RegisterFile/N24625 ) );
  AOI22_X1 U84402 ( .A1(n104855), .A2(n81423), .B1(n72262), .B2(n106014), .ZN(
        n96738) );
  OAI21_X1 U84403 ( .B1(n106046), .B2(n106016), .A(n96739), .ZN(
        \DLX_Datapath/RegisterFile/N24624 ) );
  AOI22_X1 U84404 ( .A1(n104855), .A2(n81511), .B1(n72111), .B2(n81583), .ZN(
        n96739) );
  OAI21_X1 U84405 ( .B1(n106266), .B2(n106016), .A(n96740), .ZN(
        \DLX_Datapath/RegisterFile/N24619 ) );
  AOI22_X1 U84406 ( .A1(n104855), .A2(n81327), .B1(n69629), .B2(n106014), .ZN(
        n96740) );
  NOR2_X1 U84407 ( .A1(n96741), .A2(n96717), .ZN(n81583) );
  NOR2_X1 U84408 ( .A1(n96679), .A2(n96741), .ZN(n81582) );
  NOR2_X1 U84409 ( .A1(n81580), .A2(n105091), .ZN(n96741) );
  NAND2_X1 U84410 ( .A1(n105129), .A2(n95132), .ZN(n81580) );
  OAI21_X1 U84411 ( .B1(n106147), .B2(n105401), .A(n96743), .ZN(
        \DLX_Datapath/RegisterFile/N24618 ) );
  AOI22_X1 U84412 ( .A1(n104873), .A2(n94667), .B1(n105399), .B2(n70330), .ZN(
        n96743) );
  OAI21_X1 U84413 ( .B1(n105971), .B2(n105401), .A(n96746), .ZN(
        \DLX_Datapath/RegisterFile/N24617 ) );
  AOI22_X1 U84414 ( .A1(n104872), .A2(n94670), .B1(n105398), .B2(n70472), .ZN(
        n96746) );
  OAI21_X1 U84415 ( .B1(n106137), .B2(n105401), .A(n96747), .ZN(
        \DLX_Datapath/RegisterFile/N24616 ) );
  AOI22_X1 U84416 ( .A1(n104872), .A2(n94672), .B1(n105399), .B2(n107241), 
        .ZN(n96747) );
  OAI21_X1 U84417 ( .B1(n106211), .B2(n105401), .A(n96748), .ZN(
        \DLX_Datapath/RegisterFile/N24615 ) );
  AOI22_X1 U84418 ( .A1(n104872), .A2(n94674), .B1(n105398), .B2(n107780), 
        .ZN(n96748) );
  OAI21_X1 U84419 ( .B1(n81306), .B2(n105401), .A(n96749), .ZN(
        \DLX_Datapath/RegisterFile/N24614 ) );
  AOI22_X1 U84420 ( .A1(n104873), .A2(n94676), .B1(n105399), .B2(n74032), .ZN(
        n96749) );
  OAI21_X1 U84421 ( .B1(n106099), .B2(n105401), .A(n96750), .ZN(
        \DLX_Datapath/RegisterFile/N24613 ) );
  AOI22_X1 U84422 ( .A1(n104872), .A2(n94678), .B1(n105398), .B2(n70619), .ZN(
        n96750) );
  OAI21_X1 U84423 ( .B1(n106255), .B2(n105401), .A(n96751), .ZN(
        \DLX_Datapath/RegisterFile/N24612 ) );
  AOI22_X1 U84424 ( .A1(n96744), .A2(n94680), .B1(n105399), .B2(n110779), .ZN(
        n96751) );
  OAI21_X1 U84425 ( .B1(n105992), .B2(n105401), .A(n96752), .ZN(
        \DLX_Datapath/RegisterFile/N24611 ) );
  AOI22_X1 U84426 ( .A1(n104872), .A2(n94682), .B1(n105398), .B2(n110880), 
        .ZN(n96752) );
  OAI21_X1 U84427 ( .B1(n106333), .B2(n105401), .A(n96753), .ZN(
        \DLX_Datapath/RegisterFile/N24610 ) );
  AOI22_X1 U84428 ( .A1(n104872), .A2(n94684), .B1(n105398), .B2(n110474), 
        .ZN(n96753) );
  OAI21_X1 U84429 ( .B1(n106191), .B2(n105400), .A(n96754), .ZN(
        \DLX_Datapath/RegisterFile/N24609 ) );
  AOI22_X1 U84430 ( .A1(n104873), .A2(n94686), .B1(n105398), .B2(n110256), 
        .ZN(n96754) );
  OAI21_X1 U84431 ( .B1(n106129), .B2(n105400), .A(n96755), .ZN(
        \DLX_Datapath/RegisterFile/N24608 ) );
  AOI22_X1 U84432 ( .A1(n104872), .A2(n94688), .B1(n105398), .B2(n110573), 
        .ZN(n96755) );
  OAI21_X1 U84433 ( .B1(n81318), .B2(n105400), .A(n96756), .ZN(
        \DLX_Datapath/RegisterFile/N24607 ) );
  AOI22_X1 U84434 ( .A1(n104872), .A2(n94690), .B1(n105398), .B2(n110364), 
        .ZN(n96756) );
  OAI21_X1 U84435 ( .B1(n106162), .B2(n105400), .A(n96757), .ZN(
        \DLX_Datapath/RegisterFile/N24606 ) );
  AOI22_X1 U84436 ( .A1(n96744), .A2(n94692), .B1(n96745), .B2(n110040), .ZN(
        n96757) );
  OAI21_X1 U84437 ( .B1(n106104), .B2(n105400), .A(n96758), .ZN(
        \DLX_Datapath/RegisterFile/N24605 ) );
  AOI22_X1 U84438 ( .A1(n104873), .A2(n94694), .B1(n96745), .B2(n110147), .ZN(
        n96758) );
  OAI21_X1 U84439 ( .B1(n106219), .B2(n105400), .A(n96759), .ZN(
        \DLX_Datapath/RegisterFile/N24604 ) );
  AOI22_X1 U84440 ( .A1(n96744), .A2(n94696), .B1(n96745), .B2(n109931), .ZN(
        n96759) );
  OAI21_X1 U84441 ( .B1(n106109), .B2(n105400), .A(n96760), .ZN(
        \DLX_Datapath/RegisterFile/N24603 ) );
  AOI22_X1 U84442 ( .A1(n104872), .A2(n94698), .B1(n96745), .B2(n109814), .ZN(
        n96760) );
  OAI21_X1 U84443 ( .B1(n106231), .B2(n105400), .A(n96761), .ZN(
        \DLX_Datapath/RegisterFile/N24602 ) );
  AOI22_X1 U84444 ( .A1(n104872), .A2(n94700), .B1(n105399), .B2(n108188), 
        .ZN(n96761) );
  OAI21_X1 U84445 ( .B1(n106170), .B2(n105400), .A(n96762), .ZN(
        \DLX_Datapath/RegisterFile/N24601 ) );
  AOI22_X1 U84446 ( .A1(n104873), .A2(n94702), .B1(n96745), .B2(n108311), .ZN(
        n96762) );
  OAI21_X1 U84447 ( .B1(n106236), .B2(n105400), .A(n96763), .ZN(
        \DLX_Datapath/RegisterFile/N24600 ) );
  AOI22_X1 U84448 ( .A1(n104873), .A2(n94704), .B1(n96745), .B2(n108422), .ZN(
        n96763) );
  OAI21_X1 U84449 ( .B1(n106070), .B2(n105400), .A(n96764), .ZN(
        \DLX_Datapath/RegisterFile/N24599 ) );
  AOI22_X1 U84450 ( .A1(n96744), .A2(n94706), .B1(n96745), .B2(n107660), .ZN(
        n96764) );
  OAI21_X1 U84451 ( .B1(n106197), .B2(n105400), .A(n96765), .ZN(
        \DLX_Datapath/RegisterFile/N24598 ) );
  AOI22_X1 U84452 ( .A1(n96744), .A2(n94708), .B1(n105398), .B2(n109578), .ZN(
        n96765) );
  OAI21_X1 U84453 ( .B1(n81278), .B2(n105401), .A(n96766), .ZN(
        \DLX_Datapath/RegisterFile/N24597 ) );
  AOI22_X1 U84454 ( .A1(n104872), .A2(n94710), .B1(n105399), .B2(n108539), 
        .ZN(n96766) );
  OAI21_X1 U84455 ( .B1(n106158), .B2(n105401), .A(n96767), .ZN(
        \DLX_Datapath/RegisterFile/N24596 ) );
  AOI22_X1 U84456 ( .A1(n96744), .A2(n94712), .B1(n105398), .B2(n109683), .ZN(
        n96767) );
  OAI21_X1 U84457 ( .B1(n106114), .B2(n105400), .A(n96768), .ZN(
        \DLX_Datapath/RegisterFile/N24595 ) );
  AOI22_X1 U84458 ( .A1(n104872), .A2(n94714), .B1(n105399), .B2(n109467), 
        .ZN(n96768) );
  OAI21_X1 U84459 ( .B1(n81588), .B2(n105401), .A(n96769), .ZN(
        \DLX_Datapath/RegisterFile/N24594 ) );
  AOI22_X1 U84460 ( .A1(n104873), .A2(n81259), .B1(n105398), .B2(n109004), 
        .ZN(n96769) );
  OAI21_X1 U84461 ( .B1(n81267), .B2(n105401), .A(n96770), .ZN(
        \DLX_Datapath/RegisterFile/N24593 ) );
  AOI22_X1 U84462 ( .A1(n104873), .A2(n94717), .B1(n105399), .B2(n109352), 
        .ZN(n96770) );
  OAI21_X1 U84463 ( .B1(n106043), .B2(n105400), .A(n96771), .ZN(
        \DLX_Datapath/RegisterFile/N24592 ) );
  AOI22_X1 U84464 ( .A1(n96744), .A2(n94719), .B1(n105398), .B2(n109234), .ZN(
        n96771) );
  OAI21_X1 U84465 ( .B1(n106051), .B2(n105401), .A(n96772), .ZN(
        \DLX_Datapath/RegisterFile/N24591 ) );
  AOI22_X1 U84466 ( .A1(n104873), .A2(n94721), .B1(n105399), .B2(n109126), 
        .ZN(n96772) );
  OAI21_X1 U84467 ( .B1(n106093), .B2(n105400), .A(n96773), .ZN(
        \DLX_Datapath/RegisterFile/N24590 ) );
  AOI22_X1 U84468 ( .A1(n104872), .A2(n94723), .B1(n105398), .B2(n108661), 
        .ZN(n96773) );
  OAI21_X1 U84469 ( .B1(n106054), .B2(n105401), .A(n96774), .ZN(
        \DLX_Datapath/RegisterFile/N24589 ) );
  AOI22_X1 U84470 ( .A1(n104873), .A2(n94725), .B1(n105399), .B2(n108888), 
        .ZN(n96774) );
  OAI21_X1 U84471 ( .B1(n105218), .B2(n105401), .A(n96775), .ZN(
        \DLX_Datapath/RegisterFile/N24588 ) );
  AOI22_X1 U84472 ( .A1(n104873), .A2(n94727), .B1(n105399), .B2(n108776), 
        .ZN(n96775) );
  OAI21_X1 U84473 ( .B1(n81262), .B2(n105400), .A(n96776), .ZN(
        \DLX_Datapath/RegisterFile/N24587 ) );
  AOI22_X1 U84474 ( .A1(n104872), .A2(n94729), .B1(n105398), .B2(n107316), 
        .ZN(n96776) );
  NOR2_X1 U84475 ( .A1(n96717), .A2(n96777), .ZN(n96745) );
  AOI21_X1 U84476 ( .B1(n105205), .B2(n96679), .A(n94663), .ZN(n96717) );
  NOR2_X1 U84477 ( .A1(n96679), .A2(n96777), .ZN(n96744) );
  NOR2_X1 U84478 ( .A1(n96742), .A2(n105094), .ZN(n96777) );
  OR2_X1 U84479 ( .A1(n96558), .A2(n95131), .ZN(n96679) );
  NAND2_X1 U84480 ( .A1(n105130), .A2(n94505), .ZN(n96742) );
  OAI21_X1 U84481 ( .B1(n106147), .B2(n106038), .A(n96778), .ZN(
        \DLX_Datapath/RegisterFile/N24586 ) );
  AOI22_X1 U84482 ( .A1(n106035), .A2(n81360), .B1(n70331), .B2(n106034), .ZN(
        n96778) );
  OAI21_X1 U84483 ( .B1(n106037), .B2(n81651), .A(n96779), .ZN(
        \DLX_Datapath/RegisterFile/N24585 ) );
  AOI22_X1 U84484 ( .A1(n94511), .A2(n81528), .B1(n70473), .B2(n106034), .ZN(
        n96779) );
  OAI21_X1 U84485 ( .B1(n106210), .B2(n106038), .A(n96780), .ZN(
        \DLX_Datapath/RegisterFile/N24583 ) );
  AOI22_X1 U84486 ( .A1(n106035), .A2(n81301), .B1(n70187), .B2(n81529), .ZN(
        n96780) );
  OAI21_X1 U84487 ( .B1(n106099), .B2(n106038), .A(n96781), .ZN(
        \DLX_Datapath/RegisterFile/N24581 ) );
  AOI22_X1 U84488 ( .A1(n94516), .A2(n106035), .B1(n70620), .B2(n81529), .ZN(
        n96781) );
  OAI21_X1 U84489 ( .B1(n81270), .B2(n106038), .A(n96782), .ZN(
        \DLX_Datapath/RegisterFile/N24580 ) );
  AOI22_X1 U84490 ( .A1(n106035), .A2(n81272), .B1(n74174), .B2(n106034), .ZN(
        n96782) );
  OAI21_X1 U84491 ( .B1(n106037), .B2(n105991), .A(n96783), .ZN(
        \DLX_Datapath/RegisterFile/N24579 ) );
  AOI22_X1 U84492 ( .A1(n94519), .A2(n106036), .B1(n74314), .B2(n81529), .ZN(
        n96783) );
  OAI21_X1 U84493 ( .B1(n106332), .B2(n106038), .A(n96784), .ZN(
        \DLX_Datapath/RegisterFile/N24578 ) );
  AOI22_X1 U84494 ( .A1(n106036), .A2(n80192), .B1(n73750), .B2(n106033), .ZN(
        n96784) );
  OAI21_X1 U84495 ( .B1(n106129), .B2(n106038), .A(n96785), .ZN(
        \DLX_Datapath/RegisterFile/N24576 ) );
  AOI22_X1 U84496 ( .A1(n94523), .A2(n81528), .B1(n73891), .B2(n81529), .ZN(
        n96785) );
  OAI21_X1 U84497 ( .B1(n106104), .B2(n106038), .A(n96786), .ZN(
        \DLX_Datapath/RegisterFile/N24573 ) );
  AOI22_X1 U84498 ( .A1(n94527), .A2(n81528), .B1(n73307), .B2(n81529), .ZN(
        n96786) );
  OAI21_X1 U84499 ( .B1(n106218), .B2(n106038), .A(n96787), .ZN(
        \DLX_Datapath/RegisterFile/N24572 ) );
  AOI22_X1 U84500 ( .A1(n106036), .A2(n81297), .B1(n73023), .B2(n81529), .ZN(
        n96787) );
  OAI21_X1 U84501 ( .B1(n106109), .B2(n106038), .A(n96788), .ZN(
        \DLX_Datapath/RegisterFile/N24571 ) );
  AOI22_X1 U84502 ( .A1(n94530), .A2(n81528), .B1(n72873), .B2(n81529), .ZN(
        n96788) );
  OAI21_X1 U84503 ( .B1(n106170), .B2(n106038), .A(n96789), .ZN(
        \DLX_Datapath/RegisterFile/N24569 ) );
  AOI22_X1 U84504 ( .A1(n106036), .A2(n106167), .B1(n70928), .B2(n106033), 
        .ZN(n96789) );
  OAI21_X1 U84505 ( .B1(n106070), .B2(n106038), .A(n96790), .ZN(
        \DLX_Datapath/RegisterFile/N24567 ) );
  AOI22_X1 U84506 ( .A1(n106035), .A2(n81453), .B1(n70034), .B2(n106033), .ZN(
        n96790) );
  OAI21_X1 U84507 ( .B1(n81310), .B2(n106037), .A(n96791), .ZN(
        \DLX_Datapath/RegisterFile/N24566 ) );
  AOI22_X1 U84508 ( .A1(n94536), .A2(n81528), .B1(n72563), .B2(n106034), .ZN(
        n96791) );
  OAI21_X1 U84509 ( .B1(n106158), .B2(n106037), .A(n96792), .ZN(
        \DLX_Datapath/RegisterFile/N24564 ) );
  AOI22_X1 U84510 ( .A1(n106036), .A2(n81351), .B1(n72705), .B2(n106034), .ZN(
        n96792) );
  OAI21_X1 U84511 ( .B1(n106114), .B2(n106038), .A(n96793), .ZN(
        \DLX_Datapath/RegisterFile/N24563 ) );
  AOI22_X1 U84512 ( .A1(n106019), .A2(n81528), .B1(n72415), .B2(n106033), .ZN(
        n96793) );
  OAI21_X1 U84513 ( .B1(n81588), .B2(n106038), .A(n96794), .ZN(
        \DLX_Datapath/RegisterFile/N24562 ) );
  AOI22_X1 U84514 ( .A1(n94541), .A2(n81528), .B1(n71815), .B2(n106034), .ZN(
        n96794) );
  OAI21_X1 U84515 ( .B1(n106044), .B2(n106037), .A(n96795), .ZN(
        \DLX_Datapath/RegisterFile/N24560 ) );
  AOI22_X1 U84516 ( .A1(n105624), .A2(n106036), .B1(n72113), .B2(n106033), 
        .ZN(n96795) );
  OAI21_X1 U84517 ( .B1(n81501), .B2(n106037), .A(n96796), .ZN(
        \DLX_Datapath/RegisterFile/N24559 ) );
  AOI22_X1 U84518 ( .A1(n94546), .A2(n106035), .B1(n71969), .B2(n106034), .ZN(
        n96796) );
  OAI21_X1 U84519 ( .B1(n106093), .B2(n106038), .A(n96797), .ZN(
        \DLX_Datapath/RegisterFile/N24558 ) );
  AOI22_X1 U84520 ( .A1(n94548), .A2(n106036), .B1(n71371), .B2(n106033), .ZN(
        n96797) );
  OAI21_X1 U84521 ( .B1(n106054), .B2(n106037), .A(n96798), .ZN(
        \DLX_Datapath/RegisterFile/N24557 ) );
  AOI22_X1 U84522 ( .A1(n105911), .A2(n106035), .B1(n71666), .B2(n106034), 
        .ZN(n96798) );
  OAI21_X1 U84523 ( .B1(n81262), .B2(n106037), .A(n96799), .ZN(
        \DLX_Datapath/RegisterFile/N24555 ) );
  AOI22_X1 U84524 ( .A1(n106036), .A2(n81265), .B1(n69631), .B2(n106033), .ZN(
        n96799) );
  AOI21_X1 U84525 ( .B1(n96560), .B2(n94554), .A(n96800), .ZN(n81529) );
  NOR2_X1 U84526 ( .A1(n96801), .A2(n96800), .ZN(n81528) );
  NOR2_X1 U84527 ( .A1(n81526), .A2(n105091), .ZN(n96800) );
  NAND2_X1 U84528 ( .A1(n105129), .A2(n94555), .ZN(n81526) );
  OAI21_X1 U84529 ( .B1(n106147), .B2(n105396), .A(n96803), .ZN(
        \DLX_Datapath/RegisterFile/N24554 ) );
  AOI22_X1 U84530 ( .A1(n105395), .A2(n94559), .B1(n96805), .B2(n107880), .ZN(
        n96803) );
  OAI21_X1 U84531 ( .B1(n105971), .B2(n105397), .A(n96806), .ZN(
        \DLX_Datapath/RegisterFile/N24553 ) );
  AOI22_X1 U84532 ( .A1(n96804), .A2(n94562), .B1(n105393), .B2(n70474), .ZN(
        n96806) );
  OAI21_X1 U84533 ( .B1(n106138), .B2(n105396), .A(n96807), .ZN(
        \DLX_Datapath/RegisterFile/N24552 ) );
  AOI22_X1 U84534 ( .A1(n105395), .A2(n94564), .B1(n96805), .B2(n107242), .ZN(
        n96807) );
  OAI21_X1 U84535 ( .B1(n81299), .B2(n105396), .A(n96808), .ZN(
        \DLX_Datapath/RegisterFile/N24551 ) );
  AOI22_X1 U84536 ( .A1(n96804), .A2(n94566), .B1(n105393), .B2(n107781), .ZN(
        n96808) );
  OAI21_X1 U84537 ( .B1(n81306), .B2(n105396), .A(n96809), .ZN(
        \DLX_Datapath/RegisterFile/N24550 ) );
  AOI22_X1 U84538 ( .A1(n105395), .A2(n94568), .B1(n96805), .B2(n110682), .ZN(
        n96809) );
  OAI21_X1 U84539 ( .B1(n106099), .B2(n105397), .A(n96810), .ZN(
        \DLX_Datapath/RegisterFile/N24549 ) );
  AOI22_X1 U84540 ( .A1(n105394), .A2(n94570), .B1(n105393), .B2(n108082), 
        .ZN(n96810) );
  OAI21_X1 U84541 ( .B1(n81270), .B2(n105397), .A(n96811), .ZN(
        \DLX_Datapath/RegisterFile/N24548 ) );
  AOI22_X1 U84542 ( .A1(n105395), .A2(n94572), .B1(n96805), .B2(n110780), .ZN(
        n96811) );
  OAI21_X1 U84543 ( .B1(n105992), .B2(n105396), .A(n96812), .ZN(
        \DLX_Datapath/RegisterFile/N24547 ) );
  AOI22_X1 U84544 ( .A1(n96804), .A2(n94574), .B1(n105393), .B2(n110881), .ZN(
        n96812) );
  OAI21_X1 U84545 ( .B1(n106332), .B2(n105397), .A(n96813), .ZN(
        \DLX_Datapath/RegisterFile/N24546 ) );
  AOI22_X1 U84546 ( .A1(n96804), .A2(n94576), .B1(n105393), .B2(n110475), .ZN(
        n96813) );
  OAI21_X1 U84547 ( .B1(n81315), .B2(n105397), .A(n96814), .ZN(
        \DLX_Datapath/RegisterFile/N24545 ) );
  AOI22_X1 U84548 ( .A1(n105394), .A2(n94578), .B1(n105392), .B2(n110257), 
        .ZN(n96814) );
  OAI21_X1 U84549 ( .B1(n106129), .B2(n105397), .A(n96815), .ZN(
        \DLX_Datapath/RegisterFile/N24544 ) );
  AOI22_X1 U84550 ( .A1(n105394), .A2(n94580), .B1(n105392), .B2(n110574), 
        .ZN(n96815) );
  OAI21_X1 U84551 ( .B1(n106186), .B2(n105397), .A(n96816), .ZN(
        \DLX_Datapath/RegisterFile/N24543 ) );
  AOI22_X1 U84552 ( .A1(n105394), .A2(n94582), .B1(n105392), .B2(n110365), 
        .ZN(n96816) );
  OAI21_X1 U84553 ( .B1(n106162), .B2(n105397), .A(n96817), .ZN(
        \DLX_Datapath/RegisterFile/N24542 ) );
  AOI22_X1 U84554 ( .A1(n105394), .A2(n94584), .B1(n105392), .B2(n110041), 
        .ZN(n96817) );
  OAI21_X1 U84555 ( .B1(n106104), .B2(n105397), .A(n96818), .ZN(
        \DLX_Datapath/RegisterFile/N24541 ) );
  AOI22_X1 U84556 ( .A1(n105394), .A2(n94586), .B1(n105392), .B2(n110148), 
        .ZN(n96818) );
  OAI21_X1 U84557 ( .B1(n106220), .B2(n105397), .A(n96819), .ZN(
        \DLX_Datapath/RegisterFile/N24540 ) );
  AOI22_X1 U84558 ( .A1(n105394), .A2(n94588), .B1(n105392), .B2(n109932), 
        .ZN(n96819) );
  OAI21_X1 U84559 ( .B1(n106109), .B2(n105397), .A(n96820), .ZN(
        \DLX_Datapath/RegisterFile/N24539 ) );
  AOI22_X1 U84560 ( .A1(n105394), .A2(n94590), .B1(n105392), .B2(n109815), 
        .ZN(n96820) );
  OAI21_X1 U84561 ( .B1(n106231), .B2(n105397), .A(n96821), .ZN(
        \DLX_Datapath/RegisterFile/N24538 ) );
  AOI22_X1 U84562 ( .A1(n105394), .A2(n94592), .B1(n105392), .B2(n108189), 
        .ZN(n96821) );
  OAI21_X1 U84563 ( .B1(n106171), .B2(n105397), .A(n96822), .ZN(
        \DLX_Datapath/RegisterFile/N24537 ) );
  AOI22_X1 U84564 ( .A1(n105394), .A2(n94594), .B1(n105392), .B2(n108312), 
        .ZN(n96822) );
  OAI21_X1 U84565 ( .B1(n81281), .B2(n105397), .A(n96823), .ZN(
        \DLX_Datapath/RegisterFile/N24536 ) );
  AOI22_X1 U84566 ( .A1(n105394), .A2(n94596), .B1(n105392), .B2(n108423), 
        .ZN(n96823) );
  OAI21_X1 U84567 ( .B1(n106070), .B2(n105397), .A(n96824), .ZN(
        \DLX_Datapath/RegisterFile/N24535 ) );
  AOI22_X1 U84568 ( .A1(n105394), .A2(n94598), .B1(n105392), .B2(n107661), 
        .ZN(n96824) );
  OAI21_X1 U84569 ( .B1(n81310), .B2(n105397), .A(n96825), .ZN(
        \DLX_Datapath/RegisterFile/N24534 ) );
  AOI22_X1 U84570 ( .A1(n105394), .A2(n94600), .B1(n105393), .B2(n109579), 
        .ZN(n96825) );
  OAI21_X1 U84571 ( .B1(n81278), .B2(n105396), .A(n96826), .ZN(
        \DLX_Datapath/RegisterFile/N24533 ) );
  AOI22_X1 U84572 ( .A1(n105395), .A2(n94602), .B1(n96805), .B2(n108540), .ZN(
        n96826) );
  OAI21_X1 U84573 ( .B1(n106158), .B2(n105396), .A(n96827), .ZN(
        \DLX_Datapath/RegisterFile/N24532 ) );
  AOI22_X1 U84574 ( .A1(n105394), .A2(n94604), .B1(n105393), .B2(n109684), 
        .ZN(n96827) );
  OAI21_X1 U84575 ( .B1(n106114), .B2(n105396), .A(n96828), .ZN(
        \DLX_Datapath/RegisterFile/N24531 ) );
  AOI22_X1 U84576 ( .A1(n105395), .A2(n94606), .B1(n96805), .B2(n109468), .ZN(
        n96828) );
  OAI21_X1 U84577 ( .B1(n81588), .B2(n105396), .A(n96829), .ZN(
        \DLX_Datapath/RegisterFile/N24530 ) );
  AOI22_X1 U84578 ( .A1(n96804), .A2(n94608), .B1(n105393), .B2(n109005), .ZN(
        n96829) );
  OAI21_X1 U84579 ( .B1(n81267), .B2(n105396), .A(n96830), .ZN(
        \DLX_Datapath/RegisterFile/N24529 ) );
  AOI22_X1 U84580 ( .A1(n96804), .A2(n94610), .B1(n105393), .B2(n109353), .ZN(
        n96830) );
  OAI21_X1 U84581 ( .B1(n106045), .B2(n105396), .A(n96831), .ZN(
        \DLX_Datapath/RegisterFile/N24528 ) );
  AOI22_X1 U84582 ( .A1(n105395), .A2(n94612), .B1(n105392), .B2(n109235), 
        .ZN(n96831) );
  OAI21_X1 U84583 ( .B1(n81501), .B2(n105396), .A(n96832), .ZN(
        \DLX_Datapath/RegisterFile/N24527 ) );
  AOI22_X1 U84584 ( .A1(n96804), .A2(n94614), .B1(n105393), .B2(n109127), .ZN(
        n96832) );
  OAI21_X1 U84585 ( .B1(n106093), .B2(n105396), .A(n96833), .ZN(
        \DLX_Datapath/RegisterFile/N24526 ) );
  AOI22_X1 U84586 ( .A1(n105395), .A2(n94616), .B1(n96805), .B2(n108662), .ZN(
        n96833) );
  OAI21_X1 U84587 ( .B1(n106054), .B2(n105396), .A(n96834), .ZN(
        \DLX_Datapath/RegisterFile/N24525 ) );
  AOI22_X1 U84588 ( .A1(n105395), .A2(n94618), .B1(n105393), .B2(n108889), 
        .ZN(n96834) );
  OAI21_X1 U84589 ( .B1(n105218), .B2(n105396), .A(n96835), .ZN(
        \DLX_Datapath/RegisterFile/N24524 ) );
  AOI22_X1 U84590 ( .A1(n105395), .A2(n94620), .B1(n105393), .B2(n108777), 
        .ZN(n96835) );
  OAI21_X1 U84591 ( .B1(n81262), .B2(n105396), .A(n96836), .ZN(
        \DLX_Datapath/RegisterFile/N24523 ) );
  AOI22_X1 U84592 ( .A1(n105395), .A2(n94622), .B1(n96805), .B2(n107317), .ZN(
        n96836) );
  NOR2_X1 U84593 ( .A1(n96837), .A2(n96838), .ZN(n96805) );
  NOR2_X1 U84594 ( .A1(n96801), .A2(n96838), .ZN(n96804) );
  NOR2_X1 U84595 ( .A1(n96802), .A2(n105091), .ZN(n96838) );
  NAND2_X1 U84596 ( .A1(n94625), .A2(n105129), .ZN(n96802) );
  OAI21_X1 U84597 ( .B1(n106147), .B2(n105390), .A(n96840), .ZN(
        \DLX_Datapath/RegisterFile/N24522 ) );
  AOI22_X1 U84598 ( .A1(n105389), .A2(n81521), .B1(n96842), .B2(n107881), .ZN(
        n96840) );
  OAI21_X1 U84599 ( .B1(n105971), .B2(n105390), .A(n96843), .ZN(
        \DLX_Datapath/RegisterFile/N24521 ) );
  AOI22_X1 U84600 ( .A1(n105389), .A2(n81653), .B1(n96842), .B2(n107976), .ZN(
        n96843) );
  OAI21_X1 U84601 ( .B1(n106137), .B2(n105391), .A(n96844), .ZN(
        \DLX_Datapath/RegisterFile/N24520 ) );
  AOI22_X1 U84602 ( .A1(n105389), .A2(n81380), .B1(n96842), .B2(n107243), .ZN(
        n96844) );
  OAI21_X1 U84603 ( .B1(n81299), .B2(n105390), .A(n96845), .ZN(
        \DLX_Datapath/RegisterFile/N24519 ) );
  AOI22_X1 U84604 ( .A1(n96841), .A2(n81377), .B1(n105387), .B2(n107782), .ZN(
        n96845) );
  OAI21_X1 U84605 ( .B1(n81306), .B2(n105390), .A(n96846), .ZN(
        \DLX_Datapath/RegisterFile/N24518 ) );
  AOI22_X1 U84606 ( .A1(n105389), .A2(n81428), .B1(n96842), .B2(n110683), .ZN(
        n96846) );
  OAI21_X1 U84607 ( .B1(n106099), .B2(n105391), .A(n96847), .ZN(
        \DLX_Datapath/RegisterFile/N24517 ) );
  AOI22_X1 U84608 ( .A1(n105388), .A2(n81410), .B1(n105387), .B2(n108083), 
        .ZN(n96847) );
  OAI21_X1 U84609 ( .B1(n81270), .B2(n105391), .A(n96848), .ZN(
        \DLX_Datapath/RegisterFile/N24516 ) );
  AOI22_X1 U84610 ( .A1(n96841), .A2(n81700), .B1(n105387), .B2(n110781), .ZN(
        n96848) );
  OAI21_X1 U84611 ( .B1(n105991), .B2(n105390), .A(n96849), .ZN(
        \DLX_Datapath/RegisterFile/N24515 ) );
  AOI22_X1 U84612 ( .A1(n96841), .A2(n81632), .B1(n105387), .B2(n110882), .ZN(
        n96849) );
  OAI21_X1 U84613 ( .B1(n106332), .B2(n105391), .A(n96850), .ZN(
        \DLX_Datapath/RegisterFile/N24514 ) );
  AOI22_X1 U84614 ( .A1(n96841), .A2(n81414), .B1(n105387), .B2(n110476), .ZN(
        n96850) );
  OAI21_X1 U84615 ( .B1(n81315), .B2(n105391), .A(n96851), .ZN(
        \DLX_Datapath/RegisterFile/N24513 ) );
  AOI22_X1 U84616 ( .A1(n105388), .A2(n81317), .B1(n105386), .B2(n110258), 
        .ZN(n96851) );
  OAI21_X1 U84617 ( .B1(n106129), .B2(n105391), .A(n96852), .ZN(
        \DLX_Datapath/RegisterFile/N24512 ) );
  AOI22_X1 U84618 ( .A1(n105388), .A2(n81386), .B1(n105386), .B2(n110575), 
        .ZN(n96852) );
  OAI21_X1 U84619 ( .B1(n106187), .B2(n105391), .A(n96853), .ZN(
        \DLX_Datapath/RegisterFile/N24511 ) );
  AOI22_X1 U84620 ( .A1(n105388), .A2(n81320), .B1(n105386), .B2(n110366), 
        .ZN(n96853) );
  OAI21_X1 U84621 ( .B1(n106162), .B2(n105391), .A(n96854), .ZN(
        \DLX_Datapath/RegisterFile/N24510 ) );
  AOI22_X1 U84622 ( .A1(n105388), .A2(n81604), .B1(n105387), .B2(n110042), 
        .ZN(n96854) );
  OAI21_X1 U84623 ( .B1(n106104), .B2(n105391), .A(n96855), .ZN(
        \DLX_Datapath/RegisterFile/N24509 ) );
  AOI22_X1 U84624 ( .A1(n105388), .A2(n81405), .B1(n105386), .B2(n110149), 
        .ZN(n96855) );
  OAI21_X1 U84625 ( .B1(n106219), .B2(n105391), .A(n96856), .ZN(
        \DLX_Datapath/RegisterFile/N24508 ) );
  AOI22_X1 U84626 ( .A1(n105388), .A2(n81402), .B1(n105386), .B2(n109933), 
        .ZN(n96856) );
  OAI21_X1 U84627 ( .B1(n106109), .B2(n105391), .A(n96857), .ZN(
        \DLX_Datapath/RegisterFile/N24507 ) );
  AOI22_X1 U84628 ( .A1(n105388), .A2(n81400), .B1(n105386), .B2(n109816), 
        .ZN(n96857) );
  OAI21_X1 U84629 ( .B1(n106231), .B2(n105391), .A(n96858), .ZN(
        \DLX_Datapath/RegisterFile/N24506 ) );
  AOI22_X1 U84630 ( .A1(n105388), .A2(n81332), .B1(n105386), .B2(n108190), 
        .ZN(n96858) );
  OAI21_X1 U84631 ( .B1(n106171), .B2(n105391), .A(n96859), .ZN(
        \DLX_Datapath/RegisterFile/N24505 ) );
  AOI22_X1 U84632 ( .A1(n105388), .A2(n81373), .B1(n105386), .B2(n108313), 
        .ZN(n96859) );
  OAI21_X1 U84633 ( .B1(n81281), .B2(n105391), .A(n96860), .ZN(
        \DLX_Datapath/RegisterFile/N24504 ) );
  AOI22_X1 U84634 ( .A1(n105388), .A2(n81322), .B1(n105386), .B2(n108424), 
        .ZN(n96860) );
  OAI21_X1 U84635 ( .B1(n106070), .B2(n105391), .A(n96861), .ZN(
        \DLX_Datapath/RegisterFile/N24503 ) );
  AOI22_X1 U84636 ( .A1(n105388), .A2(n81506), .B1(n105386), .B2(n107662), 
        .ZN(n96861) );
  OAI21_X1 U84637 ( .B1(n81310), .B2(n105391), .A(n96862), .ZN(
        \DLX_Datapath/RegisterFile/N24502 ) );
  AOI22_X1 U84638 ( .A1(n105388), .A2(n81313), .B1(n105386), .B2(n109580), 
        .ZN(n96862) );
  OAI21_X1 U84639 ( .B1(n81278), .B2(n105390), .A(n96863), .ZN(
        \DLX_Datapath/RegisterFile/N24501 ) );
  AOI22_X1 U84640 ( .A1(n105389), .A2(n81330), .B1(n96842), .B2(n108541), .ZN(
        n96863) );
  OAI21_X1 U84641 ( .B1(n106158), .B2(n105390), .A(n96864), .ZN(
        \DLX_Datapath/RegisterFile/N24500 ) );
  AOI22_X1 U84642 ( .A1(n105389), .A2(n81425), .B1(n105387), .B2(n109685), 
        .ZN(n96864) );
  OAI21_X1 U84643 ( .B1(n106114), .B2(n105390), .A(n96865), .ZN(
        \DLX_Datapath/RegisterFile/N24499 ) );
  AOI22_X1 U84644 ( .A1(n105389), .A2(n81396), .B1(n96842), .B2(n109469), .ZN(
        n96865) );
  OAI21_X1 U84645 ( .B1(n81588), .B2(n105390), .A(n96866), .ZN(
        \DLX_Datapath/RegisterFile/N24498 ) );
  AOI22_X1 U84646 ( .A1(n96841), .A2(n81590), .B1(n105387), .B2(n109006), .ZN(
        n96866) );
  OAI21_X1 U84647 ( .B1(n81267), .B2(n105390), .A(n96867), .ZN(
        \DLX_Datapath/RegisterFile/N24497 ) );
  AOI22_X1 U84648 ( .A1(n96841), .A2(n81423), .B1(n105387), .B2(n109354), .ZN(
        n96867) );
  OAI21_X1 U84649 ( .B1(n106043), .B2(n105390), .A(n96868), .ZN(
        \DLX_Datapath/RegisterFile/N24496 ) );
  AOI22_X1 U84650 ( .A1(n105389), .A2(n81511), .B1(n105387), .B2(n109236), 
        .ZN(n96868) );
  OAI21_X1 U84651 ( .B1(n81501), .B2(n105390), .A(n96869), .ZN(
        \DLX_Datapath/RegisterFile/N24495 ) );
  AOI22_X1 U84652 ( .A1(n96841), .A2(n81503), .B1(n105387), .B2(n109128), .ZN(
        n96869) );
  OAI21_X1 U84653 ( .B1(n106093), .B2(n105390), .A(n96870), .ZN(
        \DLX_Datapath/RegisterFile/N24494 ) );
  AOI22_X1 U84654 ( .A1(n105389), .A2(n81417), .B1(n96842), .B2(n108663), .ZN(
        n96870) );
  OAI21_X1 U84655 ( .B1(n106054), .B2(n105390), .A(n96871), .ZN(
        \DLX_Datapath/RegisterFile/N24493 ) );
  AOI22_X1 U84656 ( .A1(n105388), .A2(n81500), .B1(n105387), .B2(n108890), 
        .ZN(n96871) );
  OAI21_X1 U84657 ( .B1(n105218), .B2(n105390), .A(n96872), .ZN(
        \DLX_Datapath/RegisterFile/N24492 ) );
  AOI22_X1 U84658 ( .A1(n105389), .A2(n81335), .B1(n105386), .B2(n108778), 
        .ZN(n96872) );
  OAI21_X1 U84659 ( .B1(n81262), .B2(n105390), .A(n96873), .ZN(
        \DLX_Datapath/RegisterFile/N24491 ) );
  AOI22_X1 U84660 ( .A1(n105389), .A2(n81327), .B1(n96842), .B2(n107318), .ZN(
        n96873) );
  NOR2_X1 U84661 ( .A1(n96837), .A2(n96874), .ZN(n96842) );
  NOR2_X1 U84662 ( .A1(n96801), .A2(n96874), .ZN(n96841) );
  NOR2_X1 U84663 ( .A1(n96839), .A2(n105091), .ZN(n96874) );
  NAND2_X1 U84664 ( .A1(n105130), .A2(n94664), .ZN(n96839) );
  OAI21_X1 U84665 ( .B1(n81358), .B2(n105385), .A(n96876), .ZN(
        \DLX_Datapath/RegisterFile/N24490 ) );
  AOI22_X1 U84666 ( .A1(n105384), .A2(n94667), .B1(n105381), .B2(n70334), .ZN(
        n96876) );
  OAI21_X1 U84667 ( .B1(n105970), .B2(n96875), .A(n96879), .ZN(
        \DLX_Datapath/RegisterFile/N24489 ) );
  AOI22_X1 U84668 ( .A1(n105383), .A2(n94670), .B1(n105381), .B2(n70476), .ZN(
        n96879) );
  OAI21_X1 U84669 ( .B1(n106135), .B2(n96875), .A(n96880), .ZN(
        \DLX_Datapath/RegisterFile/N24488 ) );
  AOI22_X1 U84670 ( .A1(n105384), .A2(n94672), .B1(n105381), .B2(n69529), .ZN(
        n96880) );
  OAI21_X1 U84671 ( .B1(n106209), .B2(n96875), .A(n96881), .ZN(
        \DLX_Datapath/RegisterFile/N24487 ) );
  AOI22_X1 U84672 ( .A1(n105383), .A2(n94674), .B1(n105381), .B2(n70190), .ZN(
        n96881) );
  OAI21_X1 U84673 ( .B1(n106204), .B2(n96875), .A(n96882), .ZN(
        \DLX_Datapath/RegisterFile/N24486 ) );
  AOI22_X1 U84674 ( .A1(n105384), .A2(n94676), .B1(n105381), .B2(n74036), .ZN(
        n96882) );
  OAI21_X1 U84675 ( .B1(n106099), .B2(n96875), .A(n96883), .ZN(
        \DLX_Datapath/RegisterFile/N24485 ) );
  AOI22_X1 U84676 ( .A1(n105383), .A2(n94678), .B1(n105381), .B2(n70623), .ZN(
        n96883) );
  OAI21_X1 U84677 ( .B1(n106255), .B2(n96875), .A(n96884), .ZN(
        \DLX_Datapath/RegisterFile/N24484 ) );
  AOI22_X1 U84678 ( .A1(n105384), .A2(n94680), .B1(n105381), .B2(n74177), .ZN(
        n96884) );
  OAI21_X1 U84679 ( .B1(n105991), .B2(n105385), .A(n96885), .ZN(
        \DLX_Datapath/RegisterFile/N24483 ) );
  AOI22_X1 U84680 ( .A1(n105383), .A2(n94682), .B1(n105381), .B2(n74317), .ZN(
        n96885) );
  OAI21_X1 U84681 ( .B1(n106332), .B2(n96875), .A(n96886), .ZN(
        \DLX_Datapath/RegisterFile/N24482 ) );
  AOI22_X1 U84682 ( .A1(n105383), .A2(n94684), .B1(n105380), .B2(n73753), .ZN(
        n96886) );
  OAI21_X1 U84683 ( .B1(n81315), .B2(n105385), .A(n96887), .ZN(
        \DLX_Datapath/RegisterFile/N24481 ) );
  AOI22_X1 U84684 ( .A1(n105382), .A2(n94686), .B1(n105380), .B2(n73457), .ZN(
        n96887) );
  OAI21_X1 U84685 ( .B1(n106129), .B2(n105385), .A(n96888), .ZN(
        \DLX_Datapath/RegisterFile/N24480 ) );
  AOI22_X1 U84686 ( .A1(n105382), .A2(n94688), .B1(n105380), .B2(n73894), .ZN(
        n96888) );
  OAI21_X1 U84687 ( .B1(n106185), .B2(n105385), .A(n96889), .ZN(
        \DLX_Datapath/RegisterFile/N24479 ) );
  AOI22_X1 U84688 ( .A1(n105382), .A2(n94690), .B1(n105380), .B2(n73606), .ZN(
        n96889) );
  OAI21_X1 U84689 ( .B1(n106162), .B2(n105385), .A(n96890), .ZN(
        \DLX_Datapath/RegisterFile/N24478 ) );
  AOI22_X1 U84690 ( .A1(n105382), .A2(n94692), .B1(n105380), .B2(n73168), .ZN(
        n96890) );
  OAI21_X1 U84691 ( .B1(n106104), .B2(n105385), .A(n96891), .ZN(
        \DLX_Datapath/RegisterFile/N24477 ) );
  AOI22_X1 U84692 ( .A1(n105382), .A2(n94694), .B1(n105380), .B2(n73310), .ZN(
        n96891) );
  OAI21_X1 U84693 ( .B1(n106220), .B2(n105385), .A(n96892), .ZN(
        \DLX_Datapath/RegisterFile/N24476 ) );
  AOI22_X1 U84694 ( .A1(n105382), .A2(n94696), .B1(n105380), .B2(n73026), .ZN(
        n96892) );
  OAI21_X1 U84695 ( .B1(n106109), .B2(n105385), .A(n96893), .ZN(
        \DLX_Datapath/RegisterFile/N24475 ) );
  AOI22_X1 U84696 ( .A1(n105382), .A2(n94698), .B1(n105380), .B2(n72876), .ZN(
        n96893) );
  OAI21_X1 U84697 ( .B1(n106231), .B2(n105385), .A(n96894), .ZN(
        \DLX_Datapath/RegisterFile/N24474 ) );
  AOI22_X1 U84698 ( .A1(n105382), .A2(n94700), .B1(n105380), .B2(n70772), .ZN(
        n96894) );
  OAI21_X1 U84699 ( .B1(n106171), .B2(n105385), .A(n96895), .ZN(
        \DLX_Datapath/RegisterFile/N24473 ) );
  AOI22_X1 U84700 ( .A1(n105382), .A2(n94702), .B1(n105380), .B2(n70931), .ZN(
        n96895) );
  OAI21_X1 U84701 ( .B1(n106238), .B2(n105385), .A(n96896), .ZN(
        \DLX_Datapath/RegisterFile/N24472 ) );
  AOI22_X1 U84702 ( .A1(n105382), .A2(n94704), .B1(n105380), .B2(n71076), .ZN(
        n96896) );
  OAI21_X1 U84703 ( .B1(n106070), .B2(n105385), .A(n96897), .ZN(
        \DLX_Datapath/RegisterFile/N24471 ) );
  AOI22_X1 U84704 ( .A1(n105382), .A2(n94706), .B1(n105380), .B2(n70037), .ZN(
        n96897) );
  OAI21_X1 U84705 ( .B1(n81310), .B2(n105385), .A(n96898), .ZN(
        \DLX_Datapath/RegisterFile/N24470 ) );
  AOI22_X1 U84706 ( .A1(n105383), .A2(n94708), .B1(n105379), .B2(n72566), .ZN(
        n96898) );
  OAI21_X1 U84707 ( .B1(n106246), .B2(n105385), .A(n96899), .ZN(
        \DLX_Datapath/RegisterFile/N24469 ) );
  AOI22_X1 U84708 ( .A1(n105384), .A2(n94710), .B1(n105379), .B2(n71225), .ZN(
        n96899) );
  OAI21_X1 U84709 ( .B1(n106158), .B2(n105385), .A(n96900), .ZN(
        \DLX_Datapath/RegisterFile/N24468 ) );
  AOI22_X1 U84710 ( .A1(n105383), .A2(n94712), .B1(n105379), .B2(n72708), .ZN(
        n96900) );
  OAI21_X1 U84711 ( .B1(n106114), .B2(n105385), .A(n96901), .ZN(
        \DLX_Datapath/RegisterFile/N24467 ) );
  AOI22_X1 U84712 ( .A1(n105384), .A2(n94714), .B1(n105379), .B2(n72418), .ZN(
        n96901) );
  OAI21_X1 U84713 ( .B1(n81588), .B2(n105385), .A(n96902), .ZN(
        \DLX_Datapath/RegisterFile/N24466 ) );
  AOI22_X1 U84714 ( .A1(n105383), .A2(n81259), .B1(n105379), .B2(n71818), .ZN(
        n96902) );
  OAI21_X1 U84715 ( .B1(n81267), .B2(n105385), .A(n96903), .ZN(
        \DLX_Datapath/RegisterFile/N24465 ) );
  AOI22_X1 U84716 ( .A1(n105384), .A2(n94717), .B1(n105379), .B2(n72267), .ZN(
        n96903) );
  OAI21_X1 U84717 ( .B1(n106046), .B2(n105385), .A(n96904), .ZN(
        \DLX_Datapath/RegisterFile/N24464 ) );
  AOI22_X1 U84718 ( .A1(n105383), .A2(n94719), .B1(n105379), .B2(n72116), .ZN(
        n96904) );
  OAI21_X1 U84719 ( .B1(n106050), .B2(n105385), .A(n96905), .ZN(
        \DLX_Datapath/RegisterFile/N24463 ) );
  AOI22_X1 U84720 ( .A1(n105384), .A2(n94721), .B1(n105379), .B2(n71972), .ZN(
        n96905) );
  OAI21_X1 U84721 ( .B1(n106093), .B2(n105385), .A(n96906), .ZN(
        \DLX_Datapath/RegisterFile/N24462 ) );
  AOI22_X1 U84722 ( .A1(n105383), .A2(n94723), .B1(n105379), .B2(n71374), .ZN(
        n96906) );
  OAI21_X1 U84723 ( .B1(n106054), .B2(n96875), .A(n96907), .ZN(
        \DLX_Datapath/RegisterFile/N24461 ) );
  AOI22_X1 U84724 ( .A1(n105384), .A2(n94725), .B1(n105379), .B2(n71669), .ZN(
        n96907) );
  OAI21_X1 U84725 ( .B1(n105218), .B2(n105385), .A(n96908), .ZN(
        \DLX_Datapath/RegisterFile/N24460 ) );
  AOI22_X1 U84726 ( .A1(n105384), .A2(n94727), .B1(n105379), .B2(n71525), .ZN(
        n96908) );
  OAI21_X1 U84727 ( .B1(n81262), .B2(n105385), .A(n96909), .ZN(
        \DLX_Datapath/RegisterFile/N24459 ) );
  AOI22_X1 U84728 ( .A1(n105383), .A2(n94729), .B1(n105379), .B2(n69634), .ZN(
        n96909) );
  AOI21_X1 U84730 ( .B1(n105205), .B2(n96801), .A(n94663), .ZN(n96837) );
  NOR2_X1 U84731 ( .A1(n96801), .A2(n96910), .ZN(n96877) );
  NOR2_X1 U84732 ( .A1(n96875), .A2(n105095), .ZN(n96910) );
  OR2_X1 U84733 ( .A1(n96558), .A2(n86230), .ZN(n96801) );
  NAND2_X1 U84734 ( .A1(n94734), .A2(n105130), .ZN(n96875) );
  OAI21_X1 U84735 ( .B1(n106032), .B2(n81651), .A(n96911), .ZN(
        \DLX_Datapath/RegisterFile/N24457 ) );
  AOI22_X1 U84736 ( .A1(n94511), .A2(n104877), .B1(n106030), .B2(n107977), 
        .ZN(n96911) );
  OAI21_X1 U84737 ( .B1(n106136), .B2(n106032), .A(n96912), .ZN(
        \DLX_Datapath/RegisterFile/N24456 ) );
  AOI22_X1 U84738 ( .A1(n104875), .A2(n81539), .B1(n106030), .B2(n107244), 
        .ZN(n96912) );
  OAI21_X1 U84739 ( .B1(n106208), .B2(n106032), .A(n96913), .ZN(
        \DLX_Datapath/RegisterFile/N24455 ) );
  AOI22_X1 U84740 ( .A1(n104876), .A2(n81301), .B1(n106030), .B2(n107783), 
        .ZN(n96913) );
  OAI21_X1 U84741 ( .B1(n106099), .B2(n106032), .A(n96914), .ZN(
        \DLX_Datapath/RegisterFile/N24453 ) );
  AOI22_X1 U84742 ( .A1(n94516), .A2(n104876), .B1(n106030), .B2(n108084), 
        .ZN(n96914) );
  OAI21_X1 U84743 ( .B1(n106032), .B2(n105990), .A(n96915), .ZN(
        \DLX_Datapath/RegisterFile/N24451 ) );
  AOI22_X1 U84744 ( .A1(n94519), .A2(n104875), .B1(n106030), .B2(n110883), 
        .ZN(n96915) );
  OAI21_X1 U84745 ( .B1(n106332), .B2(n106032), .A(n96916), .ZN(
        \DLX_Datapath/RegisterFile/N24450 ) );
  AOI22_X1 U84746 ( .A1(n104876), .A2(n80192), .B1(n106030), .B2(n110477), 
        .ZN(n96916) );
  OAI21_X1 U84747 ( .B1(n106129), .B2(n106032), .A(n96917), .ZN(
        \DLX_Datapath/RegisterFile/N24448 ) );
  AOI22_X1 U84748 ( .A1(n94523), .A2(n104877), .B1(n106030), .B2(n110576), 
        .ZN(n96917) );
  OAI21_X1 U84749 ( .B1(n106104), .B2(n106032), .A(n96918), .ZN(
        \DLX_Datapath/RegisterFile/N24445 ) );
  AOI22_X1 U84750 ( .A1(n94527), .A2(n104875), .B1(n106030), .B2(n110150), 
        .ZN(n96918) );
  OAI21_X1 U84751 ( .B1(n106221), .B2(n106032), .A(n96919), .ZN(
        \DLX_Datapath/RegisterFile/N24444 ) );
  AOI22_X1 U84752 ( .A1(n104877), .A2(n81297), .B1(n106030), .B2(n109934), 
        .ZN(n96919) );
  OAI21_X1 U84753 ( .B1(n106109), .B2(n106032), .A(n96920), .ZN(
        \DLX_Datapath/RegisterFile/N24443 ) );
  AOI22_X1 U84754 ( .A1(n94530), .A2(n104876), .B1(n106029), .B2(n109817), 
        .ZN(n96920) );
  OAI21_X1 U84755 ( .B1(n106171), .B2(n106032), .A(n96921), .ZN(
        \DLX_Datapath/RegisterFile/N24441 ) );
  AOI22_X1 U84756 ( .A1(n104875), .A2(n106167), .B1(n106029), .B2(n108314), 
        .ZN(n96921) );
  OAI21_X1 U84757 ( .B1(n106070), .B2(n81540), .A(n96922), .ZN(
        \DLX_Datapath/RegisterFile/N24439 ) );
  AOI22_X1 U84758 ( .A1(n104876), .A2(n81453), .B1(n106029), .B2(n107663), 
        .ZN(n96922) );
  OAI21_X1 U84759 ( .B1(n106200), .B2(n81540), .A(n96923), .ZN(
        \DLX_Datapath/RegisterFile/N24438 ) );
  AOI22_X1 U84760 ( .A1(n105626), .A2(n104875), .B1(n106029), .B2(n109581), 
        .ZN(n96923) );
  OAI21_X1 U84761 ( .B1(n106158), .B2(n81540), .A(n96924), .ZN(
        \DLX_Datapath/RegisterFile/N24436 ) );
  AOI22_X1 U84762 ( .A1(n104875), .A2(n81351), .B1(n106029), .B2(n109686), 
        .ZN(n96924) );
  OAI21_X1 U84763 ( .B1(n106114), .B2(n81540), .A(n96925), .ZN(
        \DLX_Datapath/RegisterFile/N24435 ) );
  AOI22_X1 U84764 ( .A1(n106020), .A2(n104875), .B1(n106029), .B2(n109470), 
        .ZN(n96925) );
  OAI21_X1 U84765 ( .B1(n81588), .B2(n106032), .A(n96926), .ZN(
        \DLX_Datapath/RegisterFile/N24434 ) );
  AOI22_X1 U84766 ( .A1(n94541), .A2(n104877), .B1(n106029), .B2(n109007), 
        .ZN(n96926) );
  OAI21_X1 U84767 ( .B1(n106044), .B2(n81540), .A(n96927), .ZN(
        \DLX_Datapath/RegisterFile/N24432 ) );
  AOI22_X1 U84768 ( .A1(n105623), .A2(n104876), .B1(n106029), .B2(n109237), 
        .ZN(n96927) );
  OAI21_X1 U84769 ( .B1(n106050), .B2(n81540), .A(n96928), .ZN(
        \DLX_Datapath/RegisterFile/N24431 ) );
  AOI22_X1 U84770 ( .A1(n105622), .A2(n104876), .B1(n106029), .B2(n109129), 
        .ZN(n96928) );
  OAI21_X1 U84771 ( .B1(n106093), .B2(n81540), .A(n96929), .ZN(
        \DLX_Datapath/RegisterFile/N24430 ) );
  AOI22_X1 U84772 ( .A1(n105621), .A2(n104875), .B1(n106029), .B2(n108664), 
        .ZN(n96929) );
  OAI21_X1 U84773 ( .B1(n106054), .B2(n81540), .A(n96930), .ZN(
        \DLX_Datapath/RegisterFile/N24429 ) );
  AOI22_X1 U84774 ( .A1(n81783), .A2(n104877), .B1(n106029), .B2(n108891), 
        .ZN(n96930) );
  OAI21_X1 U84775 ( .B1(n106268), .B2(n106032), .A(n96931), .ZN(
        \DLX_Datapath/RegisterFile/N24427 ) );
  AOI22_X1 U84776 ( .A1(n104877), .A2(n81265), .B1(n106029), .B2(n107319), 
        .ZN(n96931) );
  AOI21_X1 U84777 ( .B1(n96560), .B2(n94771), .A(n96932), .ZN(n81543) );
  NAND2_X1 U84778 ( .A1(n96558), .A2(n105205), .ZN(n96560) );
  NOR2_X1 U84780 ( .A1(n81540), .A2(n105091), .ZN(n96932) );
  NAND2_X1 U84781 ( .A1(n105129), .A2(n94772), .ZN(n81540) );
  OAI21_X1 U84782 ( .B1(n81358), .B2(n105378), .A(n96935), .ZN(
        \DLX_Datapath/RegisterFile/N24426 ) );
  AOI22_X1 U84783 ( .A1(n104862), .A2(n94559), .B1(n105377), .B2(n107883), 
        .ZN(n96935) );
  OAI21_X1 U84784 ( .B1(n105970), .B2(n96934), .A(n96938), .ZN(
        \DLX_Datapath/RegisterFile/N24425 ) );
  AOI22_X1 U84785 ( .A1(n104860), .A2(n94562), .B1(n105377), .B2(n107978), 
        .ZN(n96938) );
  OAI21_X1 U84786 ( .B1(n106136), .B2(n96934), .A(n96939), .ZN(
        \DLX_Datapath/RegisterFile/N24424 ) );
  AOI22_X1 U84787 ( .A1(n104860), .A2(n94564), .B1(n105377), .B2(n107245), 
        .ZN(n96939) );
  OAI21_X1 U84788 ( .B1(n106208), .B2(n96934), .A(n96940), .ZN(
        \DLX_Datapath/RegisterFile/N24423 ) );
  AOI22_X1 U84789 ( .A1(n104861), .A2(n94566), .B1(n105377), .B2(n107784), 
        .ZN(n96940) );
  OAI21_X1 U84790 ( .B1(n106205), .B2(n96934), .A(n96941), .ZN(
        \DLX_Datapath/RegisterFile/N24422 ) );
  AOI22_X1 U84791 ( .A1(n104862), .A2(n94568), .B1(n105377), .B2(n110685), 
        .ZN(n96941) );
  OAI21_X1 U84792 ( .B1(n106099), .B2(n96934), .A(n96942), .ZN(
        \DLX_Datapath/RegisterFile/N24421 ) );
  AOI22_X1 U84793 ( .A1(n104861), .A2(n94570), .B1(n105377), .B2(n108085), 
        .ZN(n96942) );
  OAI21_X1 U84794 ( .B1(n106256), .B2(n96934), .A(n96943), .ZN(
        \DLX_Datapath/RegisterFile/N24420 ) );
  AOI22_X1 U84795 ( .A1(n104860), .A2(n94572), .B1(n105377), .B2(n110783), 
        .ZN(n96943) );
  OAI21_X1 U84796 ( .B1(n105991), .B2(n105378), .A(n96944), .ZN(
        \DLX_Datapath/RegisterFile/N24419 ) );
  AOI22_X1 U84797 ( .A1(n104861), .A2(n94574), .B1(n105377), .B2(n74319), .ZN(
        n96944) );
  OAI21_X1 U84798 ( .B1(n106332), .B2(n96934), .A(n96945), .ZN(
        \DLX_Datapath/RegisterFile/N24418 ) );
  AOI22_X1 U84799 ( .A1(n104862), .A2(n94576), .B1(n105376), .B2(n110478), 
        .ZN(n96945) );
  OAI21_X1 U84800 ( .B1(n81315), .B2(n105378), .A(n96946), .ZN(
        \DLX_Datapath/RegisterFile/N24417 ) );
  AOI22_X1 U84801 ( .A1(n104861), .A2(n94578), .B1(n105376), .B2(n110260), 
        .ZN(n96946) );
  OAI21_X1 U84802 ( .B1(n106129), .B2(n105378), .A(n96947), .ZN(
        \DLX_Datapath/RegisterFile/N24416 ) );
  AOI22_X1 U84803 ( .A1(n104862), .A2(n94580), .B1(n105376), .B2(n110577), 
        .ZN(n96947) );
  OAI21_X1 U84804 ( .B1(n106187), .B2(n105378), .A(n96948), .ZN(
        \DLX_Datapath/RegisterFile/N24415 ) );
  AOI22_X1 U84805 ( .A1(n104860), .A2(n94582), .B1(n105376), .B2(n110368), 
        .ZN(n96948) );
  OAI21_X1 U84806 ( .B1(n106162), .B2(n105378), .A(n96949), .ZN(
        \DLX_Datapath/RegisterFile/N24414 ) );
  AOI22_X1 U84807 ( .A1(n104860), .A2(n94584), .B1(n105376), .B2(n110044), 
        .ZN(n96949) );
  OAI21_X1 U84808 ( .B1(n106104), .B2(n105378), .A(n96950), .ZN(
        \DLX_Datapath/RegisterFile/N24413 ) );
  AOI22_X1 U84809 ( .A1(n104861), .A2(n94586), .B1(n105376), .B2(n110151), 
        .ZN(n96950) );
  OAI21_X1 U84810 ( .B1(n106221), .B2(n105378), .A(n96951), .ZN(
        \DLX_Datapath/RegisterFile/N24412 ) );
  AOI22_X1 U84811 ( .A1(n104861), .A2(n94588), .B1(n105376), .B2(n109935), 
        .ZN(n96951) );
  OAI21_X1 U84812 ( .B1(n106109), .B2(n105378), .A(n96952), .ZN(
        \DLX_Datapath/RegisterFile/N24411 ) );
  AOI22_X1 U84813 ( .A1(n104862), .A2(n94590), .B1(n105376), .B2(n109818), 
        .ZN(n96952) );
  OAI21_X1 U84814 ( .B1(n106231), .B2(n105378), .A(n96953), .ZN(
        \DLX_Datapath/RegisterFile/N24410 ) );
  AOI22_X1 U84815 ( .A1(n104860), .A2(n94592), .B1(n105376), .B2(n108192), 
        .ZN(n96953) );
  OAI21_X1 U84816 ( .B1(n106171), .B2(n105378), .A(n96954), .ZN(
        \DLX_Datapath/RegisterFile/N24409 ) );
  AOI22_X1 U84817 ( .A1(n104862), .A2(n94594), .B1(n105376), .B2(n108315), 
        .ZN(n96954) );
  OAI21_X1 U84818 ( .B1(n81281), .B2(n105378), .A(n96955), .ZN(
        \DLX_Datapath/RegisterFile/N24408 ) );
  AOI22_X1 U84819 ( .A1(n104861), .A2(n94596), .B1(n105376), .B2(n108426), 
        .ZN(n96955) );
  OAI21_X1 U84820 ( .B1(n106070), .B2(n105378), .A(n96956), .ZN(
        \DLX_Datapath/RegisterFile/N24407 ) );
  AOI22_X1 U84821 ( .A1(n104862), .A2(n94598), .B1(n105376), .B2(n107664), 
        .ZN(n96956) );
  OAI21_X1 U84822 ( .B1(n81310), .B2(n105378), .A(n96957), .ZN(
        \DLX_Datapath/RegisterFile/N24406 ) );
  AOI22_X1 U84823 ( .A1(n104860), .A2(n94600), .B1(n105375), .B2(n109582), 
        .ZN(n96957) );
  OAI21_X1 U84824 ( .B1(n106244), .B2(n105378), .A(n96958), .ZN(
        \DLX_Datapath/RegisterFile/N24405 ) );
  AOI22_X1 U84825 ( .A1(n104860), .A2(n94602), .B1(n105375), .B2(n108543), 
        .ZN(n96958) );
  OAI21_X1 U84826 ( .B1(n106158), .B2(n105378), .A(n96959), .ZN(
        \DLX_Datapath/RegisterFile/N24404 ) );
  AOI22_X1 U84827 ( .A1(n104860), .A2(n94604), .B1(n105375), .B2(n109687), 
        .ZN(n96959) );
  OAI21_X1 U84828 ( .B1(n106114), .B2(n105378), .A(n96960), .ZN(
        \DLX_Datapath/RegisterFile/N24403 ) );
  AOI22_X1 U84829 ( .A1(n104861), .A2(n94606), .B1(n105375), .B2(n109471), 
        .ZN(n96960) );
  OAI21_X1 U84830 ( .B1(n81588), .B2(n105378), .A(n96961), .ZN(
        \DLX_Datapath/RegisterFile/N24402 ) );
  AOI22_X1 U84831 ( .A1(n104861), .A2(n94608), .B1(n105375), .B2(n109008), 
        .ZN(n96961) );
  OAI21_X1 U84832 ( .B1(n81267), .B2(n105378), .A(n96962), .ZN(
        \DLX_Datapath/RegisterFile/N24401 ) );
  AOI22_X1 U84833 ( .A1(n104862), .A2(n94610), .B1(n105375), .B2(n109356), 
        .ZN(n96962) );
  OAI21_X1 U84834 ( .B1(n106044), .B2(n105378), .A(n96963), .ZN(
        \DLX_Datapath/RegisterFile/N24400 ) );
  AOI22_X1 U84835 ( .A1(n104860), .A2(n94612), .B1(n105375), .B2(n109238), 
        .ZN(n96963) );
  OAI21_X1 U84836 ( .B1(n106049), .B2(n105378), .A(n96964), .ZN(
        \DLX_Datapath/RegisterFile/N24399 ) );
  AOI22_X1 U84837 ( .A1(n104861), .A2(n94614), .B1(n105375), .B2(n109130), 
        .ZN(n96964) );
  OAI21_X1 U84838 ( .B1(n106093), .B2(n105378), .A(n96965), .ZN(
        \DLX_Datapath/RegisterFile/N24398 ) );
  AOI22_X1 U84839 ( .A1(n104861), .A2(n94616), .B1(n105375), .B2(n108665), 
        .ZN(n96965) );
  OAI21_X1 U84840 ( .B1(n106054), .B2(n96934), .A(n96966), .ZN(
        \DLX_Datapath/RegisterFile/N24397 ) );
  AOI22_X1 U84841 ( .A1(n104862), .A2(n94618), .B1(n105375), .B2(n108892), 
        .ZN(n96966) );
  OAI21_X1 U84842 ( .B1(n105218), .B2(n105378), .A(n96967), .ZN(
        \DLX_Datapath/RegisterFile/N24396 ) );
  AOI22_X1 U84843 ( .A1(n104860), .A2(n94620), .B1(n105375), .B2(n108780), 
        .ZN(n96967) );
  OAI21_X1 U84844 ( .B1(n106267), .B2(n105378), .A(n96968), .ZN(
        \DLX_Datapath/RegisterFile/N24395 ) );
  AOI22_X1 U84845 ( .A1(n104862), .A2(n94622), .B1(n105375), .B2(n107320), 
        .ZN(n96968) );
  NOR2_X1 U84847 ( .A1(n96933), .A2(n96970), .ZN(n96936) );
  NOR2_X1 U84848 ( .A1(n96934), .A2(n105094), .ZN(n96970) );
  NAND2_X1 U84849 ( .A1(n105130), .A2(n94810), .ZN(n96934) );
  OAI21_X1 U84850 ( .B1(n106002), .B2(n81651), .A(n96971), .ZN(
        \DLX_Datapath/RegisterFile/N24393 ) );
  AOI22_X1 U84851 ( .A1(n81653), .A2(n104850), .B1(n104866), .B2(n107979), 
        .ZN(n96971) );
  OAI21_X1 U84852 ( .B1(n106138), .B2(n106002), .A(n96972), .ZN(
        \DLX_Datapath/RegisterFile/N24392 ) );
  AOI22_X1 U84853 ( .A1(n104850), .A2(n81380), .B1(n104866), .B2(n107246), 
        .ZN(n96972) );
  OAI21_X1 U84854 ( .B1(n106208), .B2(n106002), .A(n96973), .ZN(
        \DLX_Datapath/RegisterFile/N24391 ) );
  AOI22_X1 U84855 ( .A1(n104851), .A2(n81377), .B1(n104867), .B2(n107785), 
        .ZN(n96973) );
  OAI21_X1 U84856 ( .B1(n106205), .B2(n106002), .A(n96974), .ZN(
        \DLX_Datapath/RegisterFile/N24390 ) );
  AOI22_X1 U84857 ( .A1(n104851), .A2(n81428), .B1(n104867), .B2(n110686), 
        .ZN(n96974) );
  OAI21_X1 U84858 ( .B1(n106099), .B2(n106002), .A(n96975), .ZN(
        \DLX_Datapath/RegisterFile/N24389 ) );
  AOI22_X1 U84859 ( .A1(n104849), .A2(n81410), .B1(n104865), .B2(n108086), 
        .ZN(n96975) );
  OAI21_X1 U84860 ( .B1(n106254), .B2(n106002), .A(n96976), .ZN(
        \DLX_Datapath/RegisterFile/N24388 ) );
  AOI22_X1 U84861 ( .A1(n81700), .A2(n104849), .B1(n104867), .B2(n110784), 
        .ZN(n96976) );
  OAI21_X1 U84862 ( .B1(n106002), .B2(n105991), .A(n96977), .ZN(
        \DLX_Datapath/RegisterFile/N24387 ) );
  AOI22_X1 U84863 ( .A1(n81632), .A2(n104851), .B1(n104865), .B2(n110884), 
        .ZN(n96977) );
  OAI21_X1 U84864 ( .B1(n106332), .B2(n106002), .A(n96978), .ZN(
        \DLX_Datapath/RegisterFile/N24386 ) );
  AOI22_X1 U84865 ( .A1(n104851), .A2(n81414), .B1(n104865), .B2(n110479), 
        .ZN(n96978) );
  OAI21_X1 U84866 ( .B1(n106192), .B2(n106002), .A(n96979), .ZN(
        \DLX_Datapath/RegisterFile/N24385 ) );
  AOI22_X1 U84867 ( .A1(n104850), .A2(n81317), .B1(n104866), .B2(n110261), 
        .ZN(n96979) );
  OAI21_X1 U84868 ( .B1(n106129), .B2(n106002), .A(n96980), .ZN(
        \DLX_Datapath/RegisterFile/N24384 ) );
  AOI22_X1 U84869 ( .A1(n104849), .A2(n81386), .B1(n104867), .B2(n110578), 
        .ZN(n96980) );
  OAI21_X1 U84870 ( .B1(n106186), .B2(n106002), .A(n96981), .ZN(
        \DLX_Datapath/RegisterFile/N24383 ) );
  AOI22_X1 U84871 ( .A1(n104851), .A2(n81320), .B1(n104866), .B2(n110369), 
        .ZN(n96981) );
  OAI21_X1 U84872 ( .B1(n106162), .B2(n106002), .A(n96982), .ZN(
        \DLX_Datapath/RegisterFile/N24382 ) );
  AOI22_X1 U84873 ( .A1(n104849), .A2(n81604), .B1(n104865), .B2(n110045), 
        .ZN(n96982) );
  OAI21_X1 U84874 ( .B1(n106104), .B2(n106002), .A(n96983), .ZN(
        \DLX_Datapath/RegisterFile/N24381 ) );
  AOI22_X1 U84875 ( .A1(n104850), .A2(n81405), .B1(n104865), .B2(n110152), 
        .ZN(n96983) );
  OAI21_X1 U84876 ( .B1(n106218), .B2(n106002), .A(n96984), .ZN(
        \DLX_Datapath/RegisterFile/N24380 ) );
  AOI22_X1 U84877 ( .A1(n104849), .A2(n81402), .B1(n104866), .B2(n109936), 
        .ZN(n96984) );
  OAI21_X1 U84878 ( .B1(n106109), .B2(n81608), .A(n96985), .ZN(
        \DLX_Datapath/RegisterFile/N24379 ) );
  AOI22_X1 U84879 ( .A1(n104851), .A2(n81400), .B1(n104867), .B2(n109819), 
        .ZN(n96985) );
  OAI21_X1 U84880 ( .B1(n106171), .B2(n81608), .A(n96986), .ZN(
        \DLX_Datapath/RegisterFile/N24377 ) );
  AOI22_X1 U84881 ( .A1(n104850), .A2(n81373), .B1(n104867), .B2(n108316), 
        .ZN(n96986) );
  OAI21_X1 U84882 ( .B1(n106070), .B2(n81608), .A(n96987), .ZN(
        \DLX_Datapath/RegisterFile/N24375 ) );
  AOI22_X1 U84883 ( .A1(n104849), .A2(n81506), .B1(n104865), .B2(n107665), 
        .ZN(n96987) );
  OAI21_X1 U84884 ( .B1(n106198), .B2(n81608), .A(n96988), .ZN(
        \DLX_Datapath/RegisterFile/N24374 ) );
  AOI22_X1 U84885 ( .A1(n104850), .A2(n81313), .B1(n104865), .B2(n109583), 
        .ZN(n96988) );
  OAI21_X1 U84886 ( .B1(n106158), .B2(n81608), .A(n96989), .ZN(
        \DLX_Datapath/RegisterFile/N24372 ) );
  AOI22_X1 U84887 ( .A1(n104851), .A2(n81425), .B1(n104866), .B2(n109688), 
        .ZN(n96989) );
  OAI21_X1 U84888 ( .B1(n106114), .B2(n81608), .A(n96990), .ZN(
        \DLX_Datapath/RegisterFile/N24371 ) );
  AOI22_X1 U84889 ( .A1(n104850), .A2(n81396), .B1(n104867), .B2(n109472), 
        .ZN(n96990) );
  OAI21_X1 U84890 ( .B1(n81588), .B2(n106002), .A(n96991), .ZN(
        \DLX_Datapath/RegisterFile/N24370 ) );
  AOI22_X1 U84891 ( .A1(n104849), .A2(n81590), .B1(n104866), .B2(n109009), 
        .ZN(n96991) );
  OAI21_X1 U84892 ( .B1(n106045), .B2(n81608), .A(n96992), .ZN(
        \DLX_Datapath/RegisterFile/N24368 ) );
  AOI22_X1 U84893 ( .A1(n104849), .A2(n81511), .B1(n104865), .B2(n109239), 
        .ZN(n96992) );
  OAI21_X1 U84894 ( .B1(n106054), .B2(n106002), .A(n96993), .ZN(
        \DLX_Datapath/RegisterFile/N24365 ) );
  AOI22_X1 U84895 ( .A1(n104851), .A2(n81500), .B1(n104866), .B2(n108893), 
        .ZN(n96993) );
  OAI21_X1 U84896 ( .B1(n106269), .B2(n106002), .A(n96994), .ZN(
        \DLX_Datapath/RegisterFile/N24363 ) );
  AOI22_X1 U84897 ( .A1(n104850), .A2(n81327), .B1(n104867), .B2(n107321), 
        .ZN(n96994) );
  NOR2_X1 U84898 ( .A1(n96969), .A2(n96995), .ZN(n81611) );
  NOR2_X1 U84899 ( .A1(n96933), .A2(n96995), .ZN(n81610) );
  NOR2_X1 U84900 ( .A1(n81608), .A2(n105091), .ZN(n96995) );
  NAND2_X1 U84901 ( .A1(n105129), .A2(n94853), .ZN(n81608) );
  OAI21_X1 U84902 ( .B1(n81358), .B2(n105374), .A(n96997), .ZN(
        \DLX_Datapath/RegisterFile/N24362 ) );
  AOI22_X1 U84903 ( .A1(n104858), .A2(n94667), .B1(n105372), .B2(n107885), 
        .ZN(n96997) );
  OAI21_X1 U84904 ( .B1(n105970), .B2(n105374), .A(n97000), .ZN(
        \DLX_Datapath/RegisterFile/N24361 ) );
  AOI22_X1 U84905 ( .A1(n104858), .A2(n94670), .B1(n105372), .B2(n107980), 
        .ZN(n97000) );
  OAI21_X1 U84906 ( .B1(n106138), .B2(n105374), .A(n97001), .ZN(
        \DLX_Datapath/RegisterFile/N24360 ) );
  AOI22_X1 U84907 ( .A1(n96998), .A2(n94672), .B1(n105372), .B2(n107247), .ZN(
        n97001) );
  OAI21_X1 U84908 ( .B1(n106208), .B2(n105374), .A(n97002), .ZN(
        \DLX_Datapath/RegisterFile/N24359 ) );
  AOI22_X1 U84909 ( .A1(n104859), .A2(n94674), .B1(n105372), .B2(n107786), 
        .ZN(n97002) );
  OAI21_X1 U84910 ( .B1(n81306), .B2(n105374), .A(n97003), .ZN(
        \DLX_Datapath/RegisterFile/N24358 ) );
  AOI22_X1 U84911 ( .A1(n104858), .A2(n94676), .B1(n105372), .B2(n110687), 
        .ZN(n97003) );
  OAI21_X1 U84912 ( .B1(n106099), .B2(n105374), .A(n97004), .ZN(
        \DLX_Datapath/RegisterFile/N24357 ) );
  AOI22_X1 U84913 ( .A1(n104858), .A2(n94678), .B1(n105372), .B2(n108087), 
        .ZN(n97004) );
  OAI21_X1 U84914 ( .B1(n81270), .B2(n105374), .A(n97005), .ZN(
        \DLX_Datapath/RegisterFile/N24356 ) );
  AOI22_X1 U84915 ( .A1(n104858), .A2(n94680), .B1(n105372), .B2(n110785), 
        .ZN(n97005) );
  OAI21_X1 U84916 ( .B1(n105991), .B2(n105374), .A(n97006), .ZN(
        \DLX_Datapath/RegisterFile/N24355 ) );
  AOI22_X1 U84917 ( .A1(n104859), .A2(n94682), .B1(n105372), .B2(n110885), 
        .ZN(n97006) );
  OAI21_X1 U84918 ( .B1(n106332), .B2(n105374), .A(n97007), .ZN(
        \DLX_Datapath/RegisterFile/N24354 ) );
  AOI22_X1 U84919 ( .A1(n104858), .A2(n94684), .B1(n105371), .B2(n73757), .ZN(
        n97007) );
  OAI21_X1 U84920 ( .B1(n106193), .B2(n105373), .A(n97008), .ZN(
        \DLX_Datapath/RegisterFile/N24353 ) );
  AOI22_X1 U84921 ( .A1(n96998), .A2(n94686), .B1(n105371), .B2(n73461), .ZN(
        n97008) );
  OAI21_X1 U84922 ( .B1(n106130), .B2(n105373), .A(n97009), .ZN(
        \DLX_Datapath/RegisterFile/N24352 ) );
  AOI22_X1 U84923 ( .A1(n104858), .A2(n94688), .B1(n105371), .B2(n110579), 
        .ZN(n97009) );
  OAI21_X1 U84924 ( .B1(n106186), .B2(n105373), .A(n97010), .ZN(
        \DLX_Datapath/RegisterFile/N24351 ) );
  AOI22_X1 U84925 ( .A1(n104859), .A2(n94690), .B1(n105371), .B2(n110370), 
        .ZN(n97010) );
  OAI21_X1 U84926 ( .B1(n106163), .B2(n105373), .A(n97011), .ZN(
        \DLX_Datapath/RegisterFile/N24350 ) );
  AOI22_X1 U84927 ( .A1(n104859), .A2(n94692), .B1(n105371), .B2(n110046), 
        .ZN(n97011) );
  OAI21_X1 U84928 ( .B1(n106104), .B2(n105373), .A(n97012), .ZN(
        \DLX_Datapath/RegisterFile/N24349 ) );
  AOI22_X1 U84929 ( .A1(n96998), .A2(n94694), .B1(n105371), .B2(n110153), .ZN(
        n97012) );
  OAI21_X1 U84930 ( .B1(n106218), .B2(n105373), .A(n97013), .ZN(
        \DLX_Datapath/RegisterFile/N24348 ) );
  AOI22_X1 U84931 ( .A1(n96998), .A2(n94696), .B1(n105371), .B2(n109937), .ZN(
        n97013) );
  OAI21_X1 U84932 ( .B1(n106109), .B2(n105373), .A(n97014), .ZN(
        \DLX_Datapath/RegisterFile/N24347 ) );
  AOI22_X1 U84933 ( .A1(n104858), .A2(n94698), .B1(n105371), .B2(n109820), 
        .ZN(n97014) );
  OAI21_X1 U84934 ( .B1(n106232), .B2(n105373), .A(n97015), .ZN(
        \DLX_Datapath/RegisterFile/N24346 ) );
  AOI22_X1 U84935 ( .A1(n104859), .A2(n94700), .B1(n105371), .B2(n108194), 
        .ZN(n97015) );
  OAI21_X1 U84936 ( .B1(n106171), .B2(n105373), .A(n97016), .ZN(
        \DLX_Datapath/RegisterFile/N24345 ) );
  AOI22_X1 U84937 ( .A1(n104858), .A2(n94702), .B1(n105371), .B2(n108317), 
        .ZN(n97016) );
  OAI21_X1 U84938 ( .B1(n81281), .B2(n105373), .A(n97017), .ZN(
        \DLX_Datapath/RegisterFile/N24344 ) );
  AOI22_X1 U84939 ( .A1(n104859), .A2(n94704), .B1(n105371), .B2(n108428), 
        .ZN(n97017) );
  OAI21_X1 U84940 ( .B1(n106070), .B2(n105373), .A(n97018), .ZN(
        \DLX_Datapath/RegisterFile/N24343 ) );
  AOI22_X1 U84941 ( .A1(n104858), .A2(n94706), .B1(n105371), .B2(n107666), 
        .ZN(n97018) );
  OAI21_X1 U84942 ( .B1(n106198), .B2(n105373), .A(n97019), .ZN(
        \DLX_Datapath/RegisterFile/N24342 ) );
  AOI22_X1 U84943 ( .A1(n104859), .A2(n94708), .B1(n96999), .B2(n109584), .ZN(
        n97019) );
  OAI21_X1 U84944 ( .B1(n106243), .B2(n105374), .A(n97020), .ZN(
        \DLX_Datapath/RegisterFile/N24341 ) );
  AOI22_X1 U84945 ( .A1(n104859), .A2(n94710), .B1(n105372), .B2(n108545), 
        .ZN(n97020) );
  OAI21_X1 U84946 ( .B1(n106158), .B2(n105374), .A(n97021), .ZN(
        \DLX_Datapath/RegisterFile/N24340 ) );
  AOI22_X1 U84947 ( .A1(n104859), .A2(n94712), .B1(n96999), .B2(n109689), .ZN(
        n97021) );
  OAI21_X1 U84948 ( .B1(n106114), .B2(n105373), .A(n97022), .ZN(
        \DLX_Datapath/RegisterFile/N24339 ) );
  AOI22_X1 U84949 ( .A1(n96998), .A2(n94714), .B1(n96999), .B2(n109473), .ZN(
        n97022) );
  OAI21_X1 U84950 ( .B1(n81588), .B2(n105374), .A(n97023), .ZN(
        \DLX_Datapath/RegisterFile/N24338 ) );
  AOI22_X1 U84951 ( .A1(n104858), .A2(n81259), .B1(n105372), .B2(n109010), 
        .ZN(n97023) );
  OAI21_X1 U84952 ( .B1(n81267), .B2(n105374), .A(n97024), .ZN(
        \DLX_Datapath/RegisterFile/N24337 ) );
  AOI22_X1 U84953 ( .A1(n104858), .A2(n94717), .B1(n105372), .B2(n109358), 
        .ZN(n97024) );
  OAI21_X1 U84954 ( .B1(n106045), .B2(n105373), .A(n97025), .ZN(
        \DLX_Datapath/RegisterFile/N24336 ) );
  AOI22_X1 U84955 ( .A1(n104859), .A2(n94719), .B1(n105371), .B2(n109240), 
        .ZN(n97025) );
  OAI21_X1 U84956 ( .B1(n106049), .B2(n105374), .A(n97026), .ZN(
        \DLX_Datapath/RegisterFile/N24335 ) );
  AOI22_X1 U84957 ( .A1(n104858), .A2(n94721), .B1(n96999), .B2(n109132), .ZN(
        n97026) );
  OAI21_X1 U84958 ( .B1(n106093), .B2(n105373), .A(n97027), .ZN(
        \DLX_Datapath/RegisterFile/N24334 ) );
  AOI22_X1 U84959 ( .A1(n96998), .A2(n94723), .B1(n96999), .B2(n108667), .ZN(
        n97027) );
  OAI21_X1 U84960 ( .B1(n106054), .B2(n105374), .A(n97028), .ZN(
        \DLX_Datapath/RegisterFile/N24333 ) );
  AOI22_X1 U84961 ( .A1(n104858), .A2(n94725), .B1(n96999), .B2(n108894), .ZN(
        n97028) );
  OAI21_X1 U84962 ( .B1(n105218), .B2(n105374), .A(n97029), .ZN(
        \DLX_Datapath/RegisterFile/N24332 ) );
  AOI22_X1 U84963 ( .A1(n96998), .A2(n94727), .B1(n96999), .B2(n108782), .ZN(
        n97029) );
  OAI21_X1 U84964 ( .B1(n106266), .B2(n105373), .A(n97030), .ZN(
        \DLX_Datapath/RegisterFile/N24331 ) );
  AOI22_X1 U84965 ( .A1(n104859), .A2(n94729), .B1(n96999), .B2(n107322), .ZN(
        n97030) );
  NOR2_X1 U84966 ( .A1(n97031), .A2(n96969), .ZN(n96999) );
  AOI21_X1 U84967 ( .B1(n105199), .B2(n96933), .A(n105601), .ZN(n96969) );
  NOR2_X1 U84968 ( .A1(n96933), .A2(n97031), .ZN(n96998) );
  NOR2_X1 U84969 ( .A1(n96996), .A2(n105094), .ZN(n97031) );
  OR2_X1 U84970 ( .A1(n96558), .A2(n94848), .ZN(n96933) );
  NAND2_X1 U84971 ( .A1(n97032), .A2(n107028), .ZN(n96558) );
  NOR2_X1 U84972 ( .A1(n94851), .A2(n96488), .ZN(n97032) );
  NAND2_X1 U84973 ( .A1(n94892), .A2(n105129), .ZN(n96996) );
  NOR2_X1 U84974 ( .A1(n97033), .A2(n107126), .ZN(n96561) );
  OAI21_X1 U84975 ( .B1(n81358), .B2(n106086), .A(n97034), .ZN(
        \DLX_Datapath/RegisterFile/N24330 ) );
  AOI22_X1 U84976 ( .A1(n106084), .A2(n81360), .B1(n106081), .B2(n107886), 
        .ZN(n97034) );
  OAI21_X1 U84977 ( .B1(n81439), .B2(n81651), .A(n97035), .ZN(
        \DLX_Datapath/RegisterFile/N24329 ) );
  AOI22_X1 U84978 ( .A1(n94511), .A2(n106085), .B1(n106082), .B2(n107981), 
        .ZN(n97035) );
  OAI21_X1 U84979 ( .B1(n106136), .B2(n106086), .A(n97036), .ZN(
        \DLX_Datapath/RegisterFile/N24328 ) );
  AOI22_X1 U84980 ( .A1(n81539), .A2(n106085), .B1(n106081), .B2(n107248), 
        .ZN(n97036) );
  OAI21_X1 U84981 ( .B1(n106208), .B2(n106086), .A(n97037), .ZN(
        \DLX_Datapath/RegisterFile/N24327 ) );
  AOI22_X1 U84982 ( .A1(n106083), .A2(n81301), .B1(n106081), .B2(n107787), 
        .ZN(n97037) );
  OAI21_X1 U84983 ( .B1(n81306), .B2(n106086), .A(n97038), .ZN(
        \DLX_Datapath/RegisterFile/N24326 ) );
  AOI22_X1 U84984 ( .A1(n106084), .A2(n81308), .B1(n106081), .B2(n110688), 
        .ZN(n97038) );
  OAI21_X1 U84985 ( .B1(n106099), .B2(n106086), .A(n97039), .ZN(
        \DLX_Datapath/RegisterFile/N24325 ) );
  AOI22_X1 U84986 ( .A1(n94516), .A2(n106085), .B1(n106082), .B2(n108088), 
        .ZN(n97039) );
  OAI21_X1 U84987 ( .B1(n81270), .B2(n106086), .A(n97040), .ZN(
        \DLX_Datapath/RegisterFile/N24324 ) );
  AOI22_X1 U84988 ( .A1(n106083), .A2(n81272), .B1(n106081), .B2(n110786), 
        .ZN(n97040) );
  OAI21_X1 U84989 ( .B1(n81439), .B2(n105991), .A(n97041), .ZN(
        \DLX_Datapath/RegisterFile/N24323 ) );
  AOI22_X1 U84990 ( .A1(n94519), .A2(n106085), .B1(n106080), .B2(n110886), 
        .ZN(n97041) );
  OAI21_X1 U84991 ( .B1(n106332), .B2(n106086), .A(n97042), .ZN(
        \DLX_Datapath/RegisterFile/N24322 ) );
  AOI22_X1 U84992 ( .A1(n106084), .A2(n80192), .B1(n106081), .B2(n110480), 
        .ZN(n97042) );
  OAI21_X1 U84993 ( .B1(n106130), .B2(n106086), .A(n97043), .ZN(
        \DLX_Datapath/RegisterFile/N24320 ) );
  AOI22_X1 U84994 ( .A1(n94523), .A2(n106085), .B1(n106080), .B2(n110580), 
        .ZN(n97043) );
  OAI21_X1 U84995 ( .B1(n106163), .B2(n106086), .A(n97044), .ZN(
        \DLX_Datapath/RegisterFile/N24318 ) );
  AOI22_X1 U84996 ( .A1(n106083), .A2(n81347), .B1(n106081), .B2(n110047), 
        .ZN(n97044) );
  OAI21_X1 U84997 ( .B1(n106103), .B2(n106086), .A(n97045), .ZN(
        \DLX_Datapath/RegisterFile/N24317 ) );
  AOI22_X1 U84998 ( .A1(n94527), .A2(n106085), .B1(n106082), .B2(n110154), 
        .ZN(n97045) );
  OAI21_X1 U84999 ( .B1(n106218), .B2(n106086), .A(n97046), .ZN(
        \DLX_Datapath/RegisterFile/N24316 ) );
  AOI22_X1 U85000 ( .A1(n106083), .A2(n81297), .B1(n106081), .B2(n109938), 
        .ZN(n97046) );
  OAI21_X1 U85001 ( .B1(n106109), .B2(n106086), .A(n97047), .ZN(
        \DLX_Datapath/RegisterFile/N24315 ) );
  AOI22_X1 U85002 ( .A1(n94530), .A2(n106084), .B1(n106080), .B2(n109821), 
        .ZN(n97047) );
  OAI21_X1 U85003 ( .B1(n81439), .B2(n81451), .A(n97048), .ZN(
        \DLX_Datapath/RegisterFile/N24311 ) );
  AOI22_X1 U85004 ( .A1(n81453), .A2(n106085), .B1(n106082), .B2(n107667), 
        .ZN(n97048) );
  OAI21_X1 U85005 ( .B1(n106198), .B2(n106086), .A(n97049), .ZN(
        \DLX_Datapath/RegisterFile/N24310 ) );
  AOI22_X1 U85006 ( .A1(n105626), .A2(n106083), .B1(n106082), .B2(n109585), 
        .ZN(n97049) );
  OAI21_X1 U85007 ( .B1(n106157), .B2(n106086), .A(n97050), .ZN(
        \DLX_Datapath/RegisterFile/N24308 ) );
  AOI22_X1 U85008 ( .A1(n106084), .A2(n81351), .B1(n106081), .B2(n109690), 
        .ZN(n97050) );
  OAI21_X1 U85009 ( .B1(n106114), .B2(n106086), .A(n97051), .ZN(
        \DLX_Datapath/RegisterFile/N24307 ) );
  AOI22_X1 U85010 ( .A1(n106019), .A2(n106084), .B1(n106080), .B2(n109474), 
        .ZN(n97051) );
  OAI21_X1 U85011 ( .B1(n81588), .B2(n106086), .A(n97052), .ZN(
        \DLX_Datapath/RegisterFile/N24306 ) );
  AOI22_X1 U85012 ( .A1(n94541), .A2(n106083), .B1(n106080), .B2(n109011), 
        .ZN(n97052) );
  OAI21_X1 U85013 ( .B1(n81439), .B2(n106043), .A(n97053), .ZN(
        \DLX_Datapath/RegisterFile/N24304 ) );
  AOI22_X1 U85014 ( .A1(n105623), .A2(n106084), .B1(n106080), .B2(n109241), 
        .ZN(n97053) );
  OAI21_X1 U85015 ( .B1(n106086), .B2(n81501), .A(n97054), .ZN(
        \DLX_Datapath/RegisterFile/N24303 ) );
  AOI22_X1 U85016 ( .A1(n105622), .A2(n106085), .B1(n106082), .B2(n109133), 
        .ZN(n97054) );
  OAI21_X1 U85017 ( .B1(n106094), .B2(n106086), .A(n97055), .ZN(
        \DLX_Datapath/RegisterFile/N24302 ) );
  AOI22_X1 U85018 ( .A1(n105621), .A2(n106084), .B1(n106082), .B2(n108668), 
        .ZN(n97055) );
  OAI21_X1 U85019 ( .B1(n106086), .B2(n81498), .A(n97056), .ZN(
        \DLX_Datapath/RegisterFile/N24301 ) );
  AOI22_X1 U85020 ( .A1(n105911), .A2(n106085), .B1(n106080), .B2(n108895), 
        .ZN(n97056) );
  OAI21_X1 U85021 ( .B1(n106267), .B2(n81439), .A(n97057), .ZN(
        \DLX_Datapath/RegisterFile/N24299 ) );
  AOI22_X1 U85022 ( .A1(n106084), .A2(n81265), .B1(n106081), .B2(n107323), 
        .ZN(n97057) );
  AOI21_X1 U85023 ( .B1(n97058), .B2(n94258), .A(n104724), .ZN(n81442) );
  NOR2_X1 U85024 ( .A1(n97060), .A2(n97061), .ZN(n81441) );
  OR2_X1 U85025 ( .A1(n97059), .A2(n94999), .ZN(n97060) );
  NOR2_X1 U85026 ( .A1(n81439), .A2(n105091), .ZN(n97059) );
  NAND2_X1 U85027 ( .A1(n105127), .A2(n94934), .ZN(n81439) );
  OAI21_X1 U85028 ( .B1(n81358), .B2(n105370), .A(n97064), .ZN(
        \DLX_Datapath/RegisterFile/N24298 ) );
  AOI22_X1 U85029 ( .A1(n97065), .A2(n107887), .B1(n97066), .B2(n94559), .ZN(
        n97064) );
  OAI21_X1 U85030 ( .B1(n105970), .B2(n97063), .A(n97067), .ZN(
        \DLX_Datapath/RegisterFile/N24297 ) );
  AOI22_X1 U85031 ( .A1(n97065), .A2(n107982), .B1(n97066), .B2(n94562), .ZN(
        n97067) );
  OAI21_X1 U85032 ( .B1(n81378), .B2(n105370), .A(n97068), .ZN(
        \DLX_Datapath/RegisterFile/N24296 ) );
  AOI22_X1 U85033 ( .A1(n97065), .A2(n107249), .B1(n97066), .B2(n94564), .ZN(
        n97068) );
  OAI21_X1 U85034 ( .B1(n106208), .B2(n97063), .A(n97069), .ZN(
        \DLX_Datapath/RegisterFile/N24295 ) );
  AOI22_X1 U85035 ( .A1(n97065), .A2(n107788), .B1(n97066), .B2(n94566), .ZN(
        n97069) );
  OAI21_X1 U85036 ( .B1(n81306), .B2(n105370), .A(n97070), .ZN(
        \DLX_Datapath/RegisterFile/N24294 ) );
  AOI22_X1 U85037 ( .A1(n97065), .A2(n110689), .B1(n97066), .B2(n94568), .ZN(
        n97070) );
  OAI21_X1 U85038 ( .B1(n106101), .B2(n97063), .A(n97071), .ZN(
        \DLX_Datapath/RegisterFile/N24293 ) );
  AOI22_X1 U85039 ( .A1(n97065), .A2(n108089), .B1(n97066), .B2(n94570), .ZN(
        n97071) );
  OAI21_X1 U85040 ( .B1(n81270), .B2(n105370), .A(n97072), .ZN(
        \DLX_Datapath/RegisterFile/N24292 ) );
  AOI22_X1 U85041 ( .A1(n97065), .A2(n110787), .B1(n97066), .B2(n94572), .ZN(
        n97072) );
  OAI21_X1 U85042 ( .B1(n105991), .B2(n105370), .A(n97073), .ZN(
        \DLX_Datapath/RegisterFile/N24291 ) );
  AOI22_X1 U85043 ( .A1(n97065), .A2(n110887), .B1(n97066), .B2(n94574), .ZN(
        n97073) );
  OAI21_X1 U85044 ( .B1(n106332), .B2(n97063), .A(n97074), .ZN(
        \DLX_Datapath/RegisterFile/N24290 ) );
  AOI22_X1 U85045 ( .A1(n97065), .A2(n110481), .B1(n97066), .B2(n94576), .ZN(
        n97074) );
  OAI21_X1 U85046 ( .B1(n106190), .B2(n97063), .A(n97075), .ZN(
        \DLX_Datapath/RegisterFile/N24289 ) );
  AOI22_X1 U85047 ( .A1(n97065), .A2(n110263), .B1(n97066), .B2(n94578), .ZN(
        n97075) );
  OAI21_X1 U85048 ( .B1(n106130), .B2(n97063), .A(n97076), .ZN(
        \DLX_Datapath/RegisterFile/N24288 ) );
  AOI22_X1 U85049 ( .A1(n97065), .A2(n110581), .B1(n97066), .B2(n94580), .ZN(
        n97076) );
  OAI21_X1 U85050 ( .B1(n106188), .B2(n105370), .A(n97077), .ZN(
        \DLX_Datapath/RegisterFile/N24287 ) );
  AOI22_X1 U85051 ( .A1(n97065), .A2(n110372), .B1(n97066), .B2(n94582), .ZN(
        n97077) );
  OAI21_X1 U85052 ( .B1(n106163), .B2(n105370), .A(n97078), .ZN(
        \DLX_Datapath/RegisterFile/N24286 ) );
  AOI22_X1 U85053 ( .A1(n97065), .A2(n110048), .B1(n97066), .B2(n94584), .ZN(
        n97078) );
  OAI21_X1 U85054 ( .B1(n106103), .B2(n105370), .A(n97079), .ZN(
        \DLX_Datapath/RegisterFile/N24285 ) );
  AOI22_X1 U85055 ( .A1(n97065), .A2(n110155), .B1(n97066), .B2(n94586), .ZN(
        n97079) );
  OAI21_X1 U85056 ( .B1(n106218), .B2(n105370), .A(n97080), .ZN(
        \DLX_Datapath/RegisterFile/N24284 ) );
  AOI22_X1 U85057 ( .A1(n97065), .A2(n109939), .B1(n97066), .B2(n94588), .ZN(
        n97080) );
  OAI21_X1 U85058 ( .B1(n81398), .B2(n105370), .A(n97081), .ZN(
        \DLX_Datapath/RegisterFile/N24283 ) );
  AOI22_X1 U85059 ( .A1(n97065), .A2(n109822), .B1(n97066), .B2(n94590), .ZN(
        n97081) );
  OAI21_X1 U85060 ( .B1(n106231), .B2(n105370), .A(n97082), .ZN(
        \DLX_Datapath/RegisterFile/N24282 ) );
  AOI22_X1 U85061 ( .A1(n97065), .A2(n108196), .B1(n97066), .B2(n94592), .ZN(
        n97082) );
  OAI21_X1 U85062 ( .B1(n106171), .B2(n105370), .A(n97083), .ZN(
        \DLX_Datapath/RegisterFile/N24281 ) );
  AOI22_X1 U85063 ( .A1(n97065), .A2(n108319), .B1(n97066), .B2(n94594), .ZN(
        n97083) );
  OAI21_X1 U85064 ( .B1(n81281), .B2(n105370), .A(n97084), .ZN(
        \DLX_Datapath/RegisterFile/N24280 ) );
  AOI22_X1 U85065 ( .A1(n97065), .A2(n108430), .B1(n97066), .B2(n94596), .ZN(
        n97084) );
  OAI21_X1 U85066 ( .B1(n106070), .B2(n105370), .A(n97085), .ZN(
        \DLX_Datapath/RegisterFile/N24279 ) );
  AOI22_X1 U85067 ( .A1(n97065), .A2(n107668), .B1(n97066), .B2(n94598), .ZN(
        n97085) );
  OAI21_X1 U85068 ( .B1(n106198), .B2(n105370), .A(n97086), .ZN(
        \DLX_Datapath/RegisterFile/N24278 ) );
  AOI22_X1 U85069 ( .A1(n97065), .A2(n109586), .B1(n97066), .B2(n94600), .ZN(
        n97086) );
  OAI21_X1 U85070 ( .B1(n106245), .B2(n105370), .A(n97087), .ZN(
        \DLX_Datapath/RegisterFile/N24277 ) );
  AOI22_X1 U85071 ( .A1(n97065), .A2(n108547), .B1(n97066), .B2(n94602), .ZN(
        n97087) );
  OAI21_X1 U85072 ( .B1(n106160), .B2(n105370), .A(n97088), .ZN(
        \DLX_Datapath/RegisterFile/N24276 ) );
  AOI22_X1 U85073 ( .A1(n97065), .A2(n109691), .B1(n97066), .B2(n94604), .ZN(
        n97088) );
  OAI21_X1 U85074 ( .B1(n81394), .B2(n105370), .A(n97089), .ZN(
        \DLX_Datapath/RegisterFile/N24275 ) );
  AOI22_X1 U85075 ( .A1(n97065), .A2(n109475), .B1(n97066), .B2(n94606), .ZN(
        n97089) );
  OAI21_X1 U85076 ( .B1(n106009), .B2(n105370), .A(n97090), .ZN(
        \DLX_Datapath/RegisterFile/N24274 ) );
  AOI22_X1 U85077 ( .A1(n97065), .A2(n109012), .B1(n97066), .B2(n94608), .ZN(
        n97090) );
  OAI21_X1 U85078 ( .B1(n106260), .B2(n105370), .A(n97091), .ZN(
        \DLX_Datapath/RegisterFile/N24273 ) );
  AOI22_X1 U85079 ( .A1(n97065), .A2(n109360), .B1(n97066), .B2(n94610), .ZN(
        n97091) );
  OAI21_X1 U85080 ( .B1(n106044), .B2(n105370), .A(n97092), .ZN(
        \DLX_Datapath/RegisterFile/N24272 ) );
  AOI22_X1 U85081 ( .A1(n97065), .A2(n109242), .B1(n97066), .B2(n94612), .ZN(
        n97092) );
  OAI21_X1 U85082 ( .B1(n106051), .B2(n105370), .A(n97093), .ZN(
        \DLX_Datapath/RegisterFile/N24271 ) );
  AOI22_X1 U85083 ( .A1(n97065), .A2(n109134), .B1(n97066), .B2(n94614), .ZN(
        n97093) );
  OAI21_X1 U85084 ( .B1(n106094), .B2(n105370), .A(n97094), .ZN(
        \DLX_Datapath/RegisterFile/N24270 ) );
  AOI22_X1 U85085 ( .A1(n97065), .A2(n108669), .B1(n97066), .B2(n94616), .ZN(
        n97094) );
  OAI21_X1 U85086 ( .B1(n106053), .B2(n105370), .A(n97095), .ZN(
        \DLX_Datapath/RegisterFile/N24269 ) );
  AOI22_X1 U85087 ( .A1(n97065), .A2(n108896), .B1(n97066), .B2(n94618), .ZN(
        n97095) );
  OAI21_X1 U85088 ( .B1(n105218), .B2(n105370), .A(n97096), .ZN(
        \DLX_Datapath/RegisterFile/N24268 ) );
  AOI22_X1 U85089 ( .A1(n97065), .A2(n108784), .B1(n97066), .B2(n94620), .ZN(
        n97096) );
  OAI21_X1 U85090 ( .B1(n106269), .B2(n105370), .A(n97097), .ZN(
        \DLX_Datapath/RegisterFile/N24267 ) );
  AOI22_X1 U85091 ( .A1(n97065), .A2(n107324), .B1(n97066), .B2(n94622), .ZN(
        n97097) );
  AND2_X2 U85092 ( .A1(n97098), .A2(n97099), .ZN(n97066) );
  AND2_X2 U85093 ( .A1(n97100), .A2(n97099), .ZN(n97065) );
  OR2_X1 U85094 ( .A1(n97063), .A2(n105091), .ZN(n97099) );
  NAND2_X1 U85095 ( .A1(n94296), .A2(n105127), .ZN(n97063) );
  OAI21_X1 U85096 ( .B1(n81358), .B2(n105369), .A(n97102), .ZN(
        \DLX_Datapath/RegisterFile/N24266 ) );
  AOI22_X1 U85097 ( .A1(n97103), .A2(n81521), .B1(n97104), .B2(n107888), .ZN(
        n97102) );
  OAI21_X1 U85098 ( .B1(n105970), .B2(n97101), .A(n97105), .ZN(
        \DLX_Datapath/RegisterFile/N24265 ) );
  AOI22_X1 U85099 ( .A1(n97103), .A2(n81653), .B1(n97104), .B2(n107983), .ZN(
        n97105) );
  OAI21_X1 U85100 ( .B1(n81378), .B2(n105369), .A(n97106), .ZN(
        \DLX_Datapath/RegisterFile/N24264 ) );
  AOI22_X1 U85101 ( .A1(n97103), .A2(n81380), .B1(n97104), .B2(n107250), .ZN(
        n97106) );
  OAI21_X1 U85102 ( .B1(n106208), .B2(n97101), .A(n97107), .ZN(
        \DLX_Datapath/RegisterFile/N24263 ) );
  AOI22_X1 U85103 ( .A1(n97103), .A2(n81377), .B1(n97104), .B2(n107789), .ZN(
        n97107) );
  OAI21_X1 U85104 ( .B1(n81306), .B2(n105369), .A(n97108), .ZN(
        \DLX_Datapath/RegisterFile/N24262 ) );
  AOI22_X1 U85105 ( .A1(n97103), .A2(n81428), .B1(n97104), .B2(n110690), .ZN(
        n97108) );
  OAI21_X1 U85106 ( .B1(n106099), .B2(n97101), .A(n97109), .ZN(
        \DLX_Datapath/RegisterFile/N24261 ) );
  AOI22_X1 U85107 ( .A1(n97103), .A2(n81410), .B1(n97104), .B2(n108090), .ZN(
        n97109) );
  OAI21_X1 U85108 ( .B1(n81270), .B2(n105369), .A(n97110), .ZN(
        \DLX_Datapath/RegisterFile/N24260 ) );
  AOI22_X1 U85109 ( .A1(n97103), .A2(n81700), .B1(n97104), .B2(n110788), .ZN(
        n97110) );
  OAI21_X1 U85110 ( .B1(n105991), .B2(n105369), .A(n97111), .ZN(
        \DLX_Datapath/RegisterFile/N24259 ) );
  AOI22_X1 U85111 ( .A1(n97103), .A2(n81632), .B1(n97104), .B2(n110888), .ZN(
        n97111) );
  OAI21_X1 U85112 ( .B1(n106332), .B2(n97101), .A(n97112), .ZN(
        \DLX_Datapath/RegisterFile/N24258 ) );
  AOI22_X1 U85113 ( .A1(n97103), .A2(n81414), .B1(n97104), .B2(n110482), .ZN(
        n97112) );
  OAI21_X1 U85114 ( .B1(n106192), .B2(n97101), .A(n97113), .ZN(
        \DLX_Datapath/RegisterFile/N24257 ) );
  AOI22_X1 U85115 ( .A1(n97103), .A2(n81317), .B1(n97104), .B2(n110264), .ZN(
        n97113) );
  OAI21_X1 U85116 ( .B1(n106130), .B2(n97101), .A(n97114), .ZN(
        \DLX_Datapath/RegisterFile/N24256 ) );
  AOI22_X1 U85117 ( .A1(n97103), .A2(n81386), .B1(n97104), .B2(n110582), .ZN(
        n97114) );
  OAI21_X1 U85118 ( .B1(n106185), .B2(n105369), .A(n97115), .ZN(
        \DLX_Datapath/RegisterFile/N24255 ) );
  AOI22_X1 U85119 ( .A1(n97103), .A2(n81320), .B1(n97104), .B2(n110373), .ZN(
        n97115) );
  OAI21_X1 U85120 ( .B1(n106163), .B2(n105369), .A(n97116), .ZN(
        \DLX_Datapath/RegisterFile/N24254 ) );
  AOI22_X1 U85121 ( .A1(n97103), .A2(n81604), .B1(n97104), .B2(n110049), .ZN(
        n97116) );
  OAI21_X1 U85122 ( .B1(n106106), .B2(n105369), .A(n97117), .ZN(
        \DLX_Datapath/RegisterFile/N24253 ) );
  AOI22_X1 U85123 ( .A1(n97103), .A2(n81405), .B1(n97104), .B2(n110156), .ZN(
        n97117) );
  OAI21_X1 U85124 ( .B1(n106218), .B2(n105369), .A(n97118), .ZN(
        \DLX_Datapath/RegisterFile/N24252 ) );
  AOI22_X1 U85125 ( .A1(n97103), .A2(n81402), .B1(n97104), .B2(n109940), .ZN(
        n97118) );
  OAI21_X1 U85126 ( .B1(n81398), .B2(n105369), .A(n97119), .ZN(
        \DLX_Datapath/RegisterFile/N24251 ) );
  AOI22_X1 U85127 ( .A1(n97103), .A2(n81400), .B1(n97104), .B2(n109823), .ZN(
        n97119) );
  OAI21_X1 U85128 ( .B1(n106230), .B2(n105369), .A(n97120), .ZN(
        \DLX_Datapath/RegisterFile/N24250 ) );
  AOI22_X1 U85129 ( .A1(n97103), .A2(n81332), .B1(n97104), .B2(n108197), .ZN(
        n97120) );
  OAI21_X1 U85130 ( .B1(n106171), .B2(n105369), .A(n97121), .ZN(
        \DLX_Datapath/RegisterFile/N24249 ) );
  AOI22_X1 U85131 ( .A1(n97103), .A2(n81373), .B1(n97104), .B2(n108320), .ZN(
        n97121) );
  OAI21_X1 U85132 ( .B1(n81281), .B2(n105369), .A(n97122), .ZN(
        \DLX_Datapath/RegisterFile/N24248 ) );
  AOI22_X1 U85133 ( .A1(n97103), .A2(n81322), .B1(n97104), .B2(n108431), .ZN(
        n97122) );
  OAI21_X1 U85134 ( .B1(n106070), .B2(n105369), .A(n97123), .ZN(
        \DLX_Datapath/RegisterFile/N24247 ) );
  AOI22_X1 U85135 ( .A1(n97103), .A2(n81506), .B1(n97104), .B2(n107669), .ZN(
        n97123) );
  OAI21_X1 U85136 ( .B1(n106198), .B2(n105369), .A(n97124), .ZN(
        \DLX_Datapath/RegisterFile/N24246 ) );
  AOI22_X1 U85137 ( .A1(n97103), .A2(n81313), .B1(n97104), .B2(n109587), .ZN(
        n97124) );
  OAI21_X1 U85138 ( .B1(n106245), .B2(n105369), .A(n97125), .ZN(
        \DLX_Datapath/RegisterFile/N24245 ) );
  AOI22_X1 U85139 ( .A1(n97103), .A2(n81330), .B1(n97104), .B2(n108548), .ZN(
        n97125) );
  OAI21_X1 U85140 ( .B1(n106157), .B2(n105369), .A(n97126), .ZN(
        \DLX_Datapath/RegisterFile/N24244 ) );
  AOI22_X1 U85141 ( .A1(n97103), .A2(n81425), .B1(n97104), .B2(n109692), .ZN(
        n97126) );
  OAI21_X1 U85142 ( .B1(n81394), .B2(n105369), .A(n97127), .ZN(
        \DLX_Datapath/RegisterFile/N24243 ) );
  AOI22_X1 U85143 ( .A1(n97103), .A2(n81396), .B1(n97104), .B2(n109476), .ZN(
        n97127) );
  OAI21_X1 U85144 ( .B1(n106009), .B2(n105369), .A(n97128), .ZN(
        \DLX_Datapath/RegisterFile/N24242 ) );
  AOI22_X1 U85145 ( .A1(n97103), .A2(n81590), .B1(n97104), .B2(n109013), .ZN(
        n97128) );
  OAI21_X1 U85146 ( .B1(n106261), .B2(n105369), .A(n97129), .ZN(
        \DLX_Datapath/RegisterFile/N24241 ) );
  AOI22_X1 U85147 ( .A1(n97103), .A2(n81423), .B1(n97104), .B2(n109361), .ZN(
        n97129) );
  OAI21_X1 U85148 ( .B1(n106044), .B2(n105369), .A(n97130), .ZN(
        \DLX_Datapath/RegisterFile/N24240 ) );
  AOI22_X1 U85149 ( .A1(n97103), .A2(n81511), .B1(n97104), .B2(n109243), .ZN(
        n97130) );
  OAI21_X1 U85150 ( .B1(n106050), .B2(n105369), .A(n97131), .ZN(
        \DLX_Datapath/RegisterFile/N24239 ) );
  AOI22_X1 U85151 ( .A1(n97103), .A2(n81503), .B1(n97104), .B2(n109135), .ZN(
        n97131) );
  OAI21_X1 U85152 ( .B1(n106094), .B2(n105369), .A(n97132), .ZN(
        \DLX_Datapath/RegisterFile/N24238 ) );
  AOI22_X1 U85153 ( .A1(n97103), .A2(n81417), .B1(n97104), .B2(n108670), .ZN(
        n97132) );
  OAI21_X1 U85154 ( .B1(n106055), .B2(n105369), .A(n97133), .ZN(
        \DLX_Datapath/RegisterFile/N24237 ) );
  AOI22_X1 U85155 ( .A1(n97103), .A2(n81500), .B1(n97104), .B2(n108897), .ZN(
        n97133) );
  OAI21_X1 U85156 ( .B1(n105218), .B2(n105369), .A(n97134), .ZN(
        \DLX_Datapath/RegisterFile/N24236 ) );
  AOI22_X1 U85157 ( .A1(n97103), .A2(n81335), .B1(n97104), .B2(n108785), .ZN(
        n97134) );
  OAI21_X1 U85158 ( .B1(n106268), .B2(n105369), .A(n97135), .ZN(
        \DLX_Datapath/RegisterFile/N24235 ) );
  AOI22_X1 U85159 ( .A1(n97103), .A2(n81327), .B1(n97104), .B2(n107325), .ZN(
        n97135) );
  AND2_X2 U85160 ( .A1(n97100), .A2(n97136), .ZN(n97104) );
  AND2_X2 U85161 ( .A1(n97098), .A2(n97136), .ZN(n97103) );
  OR2_X1 U85162 ( .A1(n97101), .A2(n105091), .ZN(n97136) );
  NAND2_X1 U85163 ( .A1(n105127), .A2(n94331), .ZN(n97101) );
  OAI21_X1 U85164 ( .B1(n81358), .B2(n105368), .A(n97138), .ZN(
        \DLX_Datapath/RegisterFile/N24234 ) );
  AOI22_X1 U85165 ( .A1(n97139), .A2(n94667), .B1(n97140), .B2(n70342), .ZN(
        n97138) );
  OAI21_X1 U85166 ( .B1(n105970), .B2(n105368), .A(n97141), .ZN(
        \DLX_Datapath/RegisterFile/N24233 ) );
  AOI22_X1 U85167 ( .A1(n97139), .A2(n94670), .B1(n97140), .B2(n70484), .ZN(
        n97141) );
  OAI21_X1 U85168 ( .B1(n81378), .B2(n105368), .A(n97142), .ZN(
        \DLX_Datapath/RegisterFile/N24232 ) );
  AOI22_X1 U85169 ( .A1(n97139), .A2(n94672), .B1(n97140), .B2(n107251), .ZN(
        n97142) );
  OAI21_X1 U85170 ( .B1(n106208), .B2(n105368), .A(n97143), .ZN(
        \DLX_Datapath/RegisterFile/N24231 ) );
  AOI22_X1 U85171 ( .A1(n97139), .A2(n94674), .B1(n97140), .B2(n107790), .ZN(
        n97143) );
  OAI21_X1 U85172 ( .B1(n106205), .B2(n105368), .A(n97144), .ZN(
        \DLX_Datapath/RegisterFile/N24230 ) );
  AOI22_X1 U85173 ( .A1(n97139), .A2(n94676), .B1(n97140), .B2(n74044), .ZN(
        n97144) );
  OAI21_X1 U85174 ( .B1(n106098), .B2(n105368), .A(n97145), .ZN(
        \DLX_Datapath/RegisterFile/N24229 ) );
  AOI22_X1 U85175 ( .A1(n97139), .A2(n94678), .B1(n97140), .B2(n70631), .ZN(
        n97145) );
  OAI21_X1 U85176 ( .B1(n81270), .B2(n105368), .A(n97146), .ZN(
        \DLX_Datapath/RegisterFile/N24228 ) );
  AOI22_X1 U85177 ( .A1(n97139), .A2(n94680), .B1(n97140), .B2(n110789), .ZN(
        n97146) );
  OAI21_X1 U85178 ( .B1(n105991), .B2(n105368), .A(n97147), .ZN(
        \DLX_Datapath/RegisterFile/N24227 ) );
  AOI22_X1 U85179 ( .A1(n97139), .A2(n94682), .B1(n97140), .B2(n110889), .ZN(
        n97147) );
  OAI21_X1 U85180 ( .B1(n106332), .B2(n105368), .A(n97148), .ZN(
        \DLX_Datapath/RegisterFile/N24226 ) );
  AOI22_X1 U85181 ( .A1(n97139), .A2(n94684), .B1(n97140), .B2(n110483), .ZN(
        n97148) );
  OAI21_X1 U85182 ( .B1(n106191), .B2(n105368), .A(n97149), .ZN(
        \DLX_Datapath/RegisterFile/N24225 ) );
  AOI22_X1 U85183 ( .A1(n97139), .A2(n94686), .B1(n97140), .B2(n110265), .ZN(
        n97149) );
  OAI21_X1 U85184 ( .B1(n106130), .B2(n105368), .A(n97150), .ZN(
        \DLX_Datapath/RegisterFile/N24224 ) );
  AOI22_X1 U85185 ( .A1(n97139), .A2(n94688), .B1(n97140), .B2(n110583), .ZN(
        n97150) );
  OAI21_X1 U85186 ( .B1(n106186), .B2(n105368), .A(n97151), .ZN(
        \DLX_Datapath/RegisterFile/N24223 ) );
  AOI22_X1 U85187 ( .A1(n97139), .A2(n94690), .B1(n97140), .B2(n110374), .ZN(
        n97151) );
  OAI21_X1 U85188 ( .B1(n106163), .B2(n105368), .A(n97152), .ZN(
        \DLX_Datapath/RegisterFile/N24222 ) );
  AOI22_X1 U85189 ( .A1(n97139), .A2(n94692), .B1(n97140), .B2(n110050), .ZN(
        n97152) );
  OAI21_X1 U85190 ( .B1(n106106), .B2(n105368), .A(n97153), .ZN(
        \DLX_Datapath/RegisterFile/N24221 ) );
  AOI22_X1 U85191 ( .A1(n97139), .A2(n94694), .B1(n97140), .B2(n110157), .ZN(
        n97153) );
  OAI21_X1 U85192 ( .B1(n106218), .B2(n105368), .A(n97154), .ZN(
        \DLX_Datapath/RegisterFile/N24220 ) );
  AOI22_X1 U85193 ( .A1(n97139), .A2(n94696), .B1(n97140), .B2(n109941), .ZN(
        n97154) );
  OAI21_X1 U85194 ( .B1(n81398), .B2(n105368), .A(n97155), .ZN(
        \DLX_Datapath/RegisterFile/N24219 ) );
  AOI22_X1 U85195 ( .A1(n97139), .A2(n94698), .B1(n97140), .B2(n109824), .ZN(
        n97155) );
  OAI21_X1 U85196 ( .B1(n106231), .B2(n105368), .A(n97156), .ZN(
        \DLX_Datapath/RegisterFile/N24218 ) );
  AOI22_X1 U85197 ( .A1(n97139), .A2(n94700), .B1(n97140), .B2(n108198), .ZN(
        n97156) );
  OAI21_X1 U85198 ( .B1(n106171), .B2(n105368), .A(n97157), .ZN(
        \DLX_Datapath/RegisterFile/N24217 ) );
  AOI22_X1 U85199 ( .A1(n97139), .A2(n94702), .B1(n97140), .B2(n108321), .ZN(
        n97157) );
  OAI21_X1 U85200 ( .B1(n81281), .B2(n105368), .A(n97158), .ZN(
        \DLX_Datapath/RegisterFile/N24216 ) );
  AOI22_X1 U85201 ( .A1(n97139), .A2(n94704), .B1(n97140), .B2(n108432), .ZN(
        n97158) );
  OAI21_X1 U85202 ( .B1(n106070), .B2(n105368), .A(n97159), .ZN(
        \DLX_Datapath/RegisterFile/N24215 ) );
  AOI22_X1 U85203 ( .A1(n97139), .A2(n94706), .B1(n97140), .B2(n107670), .ZN(
        n97159) );
  OAI21_X1 U85204 ( .B1(n106198), .B2(n105368), .A(n97160), .ZN(
        \DLX_Datapath/RegisterFile/N24214 ) );
  AOI22_X1 U85205 ( .A1(n97139), .A2(n94708), .B1(n97140), .B2(n109588), .ZN(
        n97160) );
  OAI21_X1 U85206 ( .B1(n106245), .B2(n105368), .A(n97161), .ZN(
        \DLX_Datapath/RegisterFile/N24213 ) );
  AOI22_X1 U85207 ( .A1(n97139), .A2(n94710), .B1(n97140), .B2(n108549), .ZN(
        n97161) );
  OAI21_X1 U85208 ( .B1(n106159), .B2(n105368), .A(n97162), .ZN(
        \DLX_Datapath/RegisterFile/N24212 ) );
  AOI22_X1 U85209 ( .A1(n97139), .A2(n94712), .B1(n97140), .B2(n109693), .ZN(
        n97162) );
  OAI21_X1 U85210 ( .B1(n81394), .B2(n105368), .A(n97163), .ZN(
        \DLX_Datapath/RegisterFile/N24211 ) );
  AOI22_X1 U85211 ( .A1(n97139), .A2(n94714), .B1(n97140), .B2(n109477), .ZN(
        n97163) );
  OAI21_X1 U85212 ( .B1(n106009), .B2(n105368), .A(n97164), .ZN(
        \DLX_Datapath/RegisterFile/N24210 ) );
  AOI22_X1 U85213 ( .A1(n97139), .A2(n81259), .B1(n97140), .B2(n109014), .ZN(
        n97164) );
  OAI21_X1 U85214 ( .B1(n106260), .B2(n105368), .A(n97165), .ZN(
        \DLX_Datapath/RegisterFile/N24209 ) );
  AOI22_X1 U85215 ( .A1(n97139), .A2(n94717), .B1(n97140), .B2(n109362), .ZN(
        n97165) );
  OAI21_X1 U85216 ( .B1(n106044), .B2(n105368), .A(n97166), .ZN(
        \DLX_Datapath/RegisterFile/N24208 ) );
  AOI22_X1 U85217 ( .A1(n97139), .A2(n94719), .B1(n97140), .B2(n109244), .ZN(
        n97166) );
  OAI21_X1 U85218 ( .B1(n106051), .B2(n105368), .A(n97167), .ZN(
        \DLX_Datapath/RegisterFile/N24207 ) );
  AOI22_X1 U85219 ( .A1(n97139), .A2(n94721), .B1(n97140), .B2(n109136), .ZN(
        n97167) );
  OAI21_X1 U85220 ( .B1(n106094), .B2(n105368), .A(n97168), .ZN(
        \DLX_Datapath/RegisterFile/N24206 ) );
  AOI22_X1 U85221 ( .A1(n97139), .A2(n94723), .B1(n97140), .B2(n108671), .ZN(
        n97168) );
  OAI21_X1 U85222 ( .B1(n106054), .B2(n105368), .A(n97169), .ZN(
        \DLX_Datapath/RegisterFile/N24205 ) );
  AOI22_X1 U85223 ( .A1(n97139), .A2(n94725), .B1(n97140), .B2(n108898), .ZN(
        n97169) );
  OAI21_X1 U85224 ( .B1(n105218), .B2(n105368), .A(n97170), .ZN(
        \DLX_Datapath/RegisterFile/N24204 ) );
  AOI22_X1 U85225 ( .A1(n97139), .A2(n94727), .B1(n97140), .B2(n108786), .ZN(
        n97170) );
  OAI21_X1 U85226 ( .B1(n106268), .B2(n105368), .A(n97171), .ZN(
        \DLX_Datapath/RegisterFile/N24203 ) );
  AOI22_X1 U85227 ( .A1(n97139), .A2(n94729), .B1(n97140), .B2(n107326), .ZN(
        n97171) );
  AND2_X2 U85228 ( .A1(n97100), .A2(n97172), .ZN(n97140) );
  OAI21_X1 U85229 ( .B1(n94366), .B2(n97098), .A(n105602), .ZN(n97100) );
  AND2_X2 U85230 ( .A1(n97098), .A2(n97172), .ZN(n97139) );
  OR2_X1 U85231 ( .A1(n97137), .A2(n105089), .ZN(n97172) );
  NOR2_X1 U85232 ( .A1(n97061), .A2(n94999), .ZN(n97098) );
  NAND2_X1 U85233 ( .A1(n94367), .A2(n105127), .ZN(n97137) );
  OAI21_X1 U85234 ( .B1(n106059), .B2(n81651), .A(n97173), .ZN(
        \DLX_Datapath/RegisterFile/N24201 ) );
  AOI22_X1 U85235 ( .A1(n94511), .A2(n104765), .B1(n70485), .B2(n104827), .ZN(
        n97173) );
  AOI22_X1 U85237 ( .A1(n81539), .A2(n104766), .B1(n69538), .B2(n104827), .ZN(
        n97174) );
  OAI21_X1 U85238 ( .B1(n106208), .B2(n106059), .A(n97175), .ZN(
        \DLX_Datapath/RegisterFile/N24199 ) );
  AOI22_X1 U85239 ( .A1(n104765), .A2(n81301), .B1(n70199), .B2(n81479), .ZN(
        n97175) );
  OAI21_X1 U85240 ( .B1(n106206), .B2(n106059), .A(n97176), .ZN(
        \DLX_Datapath/RegisterFile/N24198 ) );
  AOI22_X1 U85241 ( .A1(n104765), .A2(n81308), .B1(n74045), .B2(n104828), .ZN(
        n97176) );
  OAI21_X1 U85242 ( .B1(n106101), .B2(n106059), .A(n97177), .ZN(
        \DLX_Datapath/RegisterFile/N24197 ) );
  AOI22_X1 U85243 ( .A1(n94516), .A2(n104764), .B1(n70632), .B2(n81479), .ZN(
        n97177) );
  OAI21_X1 U85244 ( .B1(n106256), .B2(n106059), .A(n97178), .ZN(
        \DLX_Datapath/RegisterFile/N24196 ) );
  AOI22_X1 U85245 ( .A1(n104765), .A2(n81272), .B1(n74186), .B2(n81479), .ZN(
        n97178) );
  OAI21_X1 U85246 ( .B1(n106059), .B2(n105992), .A(n97179), .ZN(
        \DLX_Datapath/RegisterFile/N24195 ) );
  AOI22_X1 U85247 ( .A1(n94519), .A2(n104764), .B1(n74326), .B2(n104827), .ZN(
        n97179) );
  OAI21_X1 U85248 ( .B1(n106330), .B2(n106059), .A(n97180), .ZN(
        \DLX_Datapath/RegisterFile/N24194 ) );
  AOI22_X1 U85249 ( .A1(n104765), .A2(n80192), .B1(n73762), .B2(n104827), .ZN(
        n97180) );
  OAI21_X1 U85250 ( .B1(n106193), .B2(n106059), .A(n97181), .ZN(
        \DLX_Datapath/RegisterFile/N24193 ) );
  AOI22_X1 U85251 ( .A1(n104766), .A2(n81474), .B1(n73466), .B2(n104827), .ZN(
        n97181) );
  OAI21_X1 U85252 ( .B1(n106130), .B2(n106059), .A(n97182), .ZN(
        \DLX_Datapath/RegisterFile/N24192 ) );
  AOI22_X1 U85253 ( .A1(n94523), .A2(n104764), .B1(n73903), .B2(n104828), .ZN(
        n97182) );
  OAI21_X1 U85254 ( .B1(n106188), .B2(n106059), .A(n97183), .ZN(
        \DLX_Datapath/RegisterFile/N24191 ) );
  AOI22_X1 U85255 ( .A1(n104764), .A2(n106060), .B1(n73615), .B2(n104828), 
        .ZN(n97183) );
  OAI21_X1 U85256 ( .B1(n106163), .B2(n106059), .A(n97184), .ZN(
        \DLX_Datapath/RegisterFile/N24190 ) );
  AOI22_X1 U85257 ( .A1(n104765), .A2(n81347), .B1(n73177), .B2(n104828), .ZN(
        n97184) );
  OAI21_X1 U85258 ( .B1(n81403), .B2(n106059), .A(n97185), .ZN(
        \DLX_Datapath/RegisterFile/N24189 ) );
  AOI22_X1 U85259 ( .A1(n94527), .A2(n104764), .B1(n73319), .B2(n104827), .ZN(
        n97185) );
  OAI21_X1 U85260 ( .B1(n106218), .B2(n106059), .A(n97186), .ZN(
        \DLX_Datapath/RegisterFile/N24188 ) );
  AOI22_X1 U85261 ( .A1(n104766), .A2(n81297), .B1(n73035), .B2(n81479), .ZN(
        n97186) );
  OAI21_X1 U85262 ( .B1(n81398), .B2(n106059), .A(n97187), .ZN(
        \DLX_Datapath/RegisterFile/N24187 ) );
  AOI22_X1 U85263 ( .A1(n94530), .A2(n104764), .B1(n72885), .B2(n104828), .ZN(
        n97187) );
  OAI21_X1 U85264 ( .B1(n106072), .B2(n106059), .A(n97188), .ZN(
        \DLX_Datapath/RegisterFile/N24183 ) );
  AOI22_X1 U85265 ( .A1(n104765), .A2(n81453), .B1(n70046), .B2(n104827), .ZN(
        n97188) );
  OAI21_X1 U85266 ( .B1(n106198), .B2(n106059), .A(n97189), .ZN(
        \DLX_Datapath/RegisterFile/N24182 ) );
  AOI22_X1 U85267 ( .A1(n105626), .A2(n104764), .B1(n72575), .B2(n104828), 
        .ZN(n97189) );
  OAI21_X1 U85268 ( .B1(n106159), .B2(n106059), .A(n97190), .ZN(
        \DLX_Datapath/RegisterFile/N24180 ) );
  AOI22_X1 U85269 ( .A1(n104766), .A2(n81351), .B1(n72717), .B2(n81479), .ZN(
        n97190) );
  OAI21_X1 U85270 ( .B1(n106114), .B2(n106059), .A(n97191), .ZN(
        \DLX_Datapath/RegisterFile/N24179 ) );
  AOI22_X1 U85271 ( .A1(n106019), .A2(n104764), .B1(n72427), .B2(n104827), 
        .ZN(n97191) );
  OAI21_X1 U85272 ( .B1(n106009), .B2(n106059), .A(n97192), .ZN(
        \DLX_Datapath/RegisterFile/N24178 ) );
  AOI22_X1 U85273 ( .A1(n94541), .A2(n104765), .B1(n71827), .B2(n104827), .ZN(
        n97192) );
  OAI21_X1 U85274 ( .B1(n106059), .B2(n81509), .A(n97193), .ZN(
        \DLX_Datapath/RegisterFile/N24176 ) );
  AOI22_X1 U85275 ( .A1(n105623), .A2(n104766), .B1(n72125), .B2(n104827), 
        .ZN(n97193) );
  OAI21_X1 U85276 ( .B1(n106059), .B2(n81501), .A(n97194), .ZN(
        \DLX_Datapath/RegisterFile/N24175 ) );
  AOI22_X1 U85277 ( .A1(n105622), .A2(n104765), .B1(n71981), .B2(n104828), 
        .ZN(n97194) );
  OAI21_X1 U85278 ( .B1(n106094), .B2(n106059), .A(n97195), .ZN(
        \DLX_Datapath/RegisterFile/N24174 ) );
  AOI22_X1 U85279 ( .A1(n105621), .A2(n104766), .B1(n71383), .B2(n104828), 
        .ZN(n97195) );
  OAI21_X1 U85280 ( .B1(n106059), .B2(n81498), .A(n97196), .ZN(
        \DLX_Datapath/RegisterFile/N24173 ) );
  AOI22_X1 U85281 ( .A1(n105911), .A2(n104766), .B1(n71678), .B2(n104828), 
        .ZN(n97196) );
  OAI21_X1 U85282 ( .B1(n106267), .B2(n106059), .A(n97197), .ZN(
        \DLX_Datapath/RegisterFile/N24171 ) );
  AOI22_X1 U85283 ( .A1(n104765), .A2(n81265), .B1(n69643), .B2(n104828), .ZN(
        n97197) );
  AOI21_X1 U85284 ( .B1(n97058), .B2(n94398), .A(n104725), .ZN(n81479) );
  NOR2_X1 U85285 ( .A1(n97199), .A2(n97061), .ZN(n81478) );
  OR2_X1 U85286 ( .A1(n97198), .A2(n95131), .ZN(n97199) );
  NOR2_X1 U85287 ( .A1(n81476), .A2(n105094), .ZN(n97198) );
  NAND2_X1 U85288 ( .A1(n105127), .A2(n94399), .ZN(n81476) );
  OAI21_X1 U85289 ( .B1(n81358), .B2(n105367), .A(n97201), .ZN(
        \DLX_Datapath/RegisterFile/N24170 ) );
  AOI22_X1 U85290 ( .A1(n97202), .A2(n94559), .B1(n97203), .B2(n107889), .ZN(
        n97201) );
  OAI21_X1 U85291 ( .B1(n105970), .B2(n105367), .A(n97204), .ZN(
        \DLX_Datapath/RegisterFile/N24169 ) );
  AOI22_X1 U85292 ( .A1(n97202), .A2(n94562), .B1(n97203), .B2(n107984), .ZN(
        n97204) );
  OAI21_X1 U85293 ( .B1(n81378), .B2(n105367), .A(n97205), .ZN(
        \DLX_Datapath/RegisterFile/N24168 ) );
  AOI22_X1 U85294 ( .A1(n97202), .A2(n94564), .B1(n97203), .B2(n107252), .ZN(
        n97205) );
  OAI21_X1 U85295 ( .B1(n106208), .B2(n105367), .A(n97206), .ZN(
        \DLX_Datapath/RegisterFile/N24167 ) );
  AOI22_X1 U85296 ( .A1(n97202), .A2(n94566), .B1(n97203), .B2(n107791), .ZN(
        n97206) );
  OAI21_X1 U85297 ( .B1(n106206), .B2(n105367), .A(n97207), .ZN(
        \DLX_Datapath/RegisterFile/N24166 ) );
  AOI22_X1 U85298 ( .A1(n97202), .A2(n94568), .B1(n97203), .B2(n110691), .ZN(
        n97207) );
  OAI21_X1 U85299 ( .B1(n106101), .B2(n105367), .A(n97208), .ZN(
        \DLX_Datapath/RegisterFile/N24165 ) );
  AOI22_X1 U85300 ( .A1(n97202), .A2(n94570), .B1(n97203), .B2(n108091), .ZN(
        n97208) );
  OAI21_X1 U85301 ( .B1(n81270), .B2(n105367), .A(n97209), .ZN(
        \DLX_Datapath/RegisterFile/N24164 ) );
  AOI22_X1 U85302 ( .A1(n97202), .A2(n94572), .B1(n97203), .B2(n110790), .ZN(
        n97209) );
  OAI21_X1 U85303 ( .B1(n105991), .B2(n105367), .A(n97210), .ZN(
        \DLX_Datapath/RegisterFile/N24163 ) );
  AOI22_X1 U85304 ( .A1(n97202), .A2(n94574), .B1(n97203), .B2(n110890), .ZN(
        n97210) );
  OAI21_X1 U85305 ( .B1(n106333), .B2(n105367), .A(n97211), .ZN(
        \DLX_Datapath/RegisterFile/N24162 ) );
  AOI22_X1 U85306 ( .A1(n97202), .A2(n94576), .B1(n97203), .B2(n110484), .ZN(
        n97211) );
  OAI21_X1 U85307 ( .B1(n106193), .B2(n105367), .A(n97212), .ZN(
        \DLX_Datapath/RegisterFile/N24161 ) );
  AOI22_X1 U85308 ( .A1(n97202), .A2(n94578), .B1(n97203), .B2(n110266), .ZN(
        n97212) );
  OAI21_X1 U85309 ( .B1(n106130), .B2(n105367), .A(n97213), .ZN(
        \DLX_Datapath/RegisterFile/N24160 ) );
  AOI22_X1 U85310 ( .A1(n97202), .A2(n94580), .B1(n97203), .B2(n110584), .ZN(
        n97213) );
  OAI21_X1 U85311 ( .B1(n106188), .B2(n105367), .A(n97214), .ZN(
        \DLX_Datapath/RegisterFile/N24159 ) );
  AOI22_X1 U85312 ( .A1(n97202), .A2(n94582), .B1(n97203), .B2(n110375), .ZN(
        n97214) );
  OAI21_X1 U85313 ( .B1(n106163), .B2(n105367), .A(n97215), .ZN(
        \DLX_Datapath/RegisterFile/N24158 ) );
  AOI22_X1 U85314 ( .A1(n97202), .A2(n94584), .B1(n97203), .B2(n110051), .ZN(
        n97215) );
  OAI21_X1 U85315 ( .B1(n106104), .B2(n105367), .A(n97216), .ZN(
        \DLX_Datapath/RegisterFile/N24157 ) );
  AOI22_X1 U85316 ( .A1(n97202), .A2(n94586), .B1(n97203), .B2(n110158), .ZN(
        n97216) );
  OAI21_X1 U85317 ( .B1(n106218), .B2(n105367), .A(n97217), .ZN(
        \DLX_Datapath/RegisterFile/N24156 ) );
  AOI22_X1 U85318 ( .A1(n97202), .A2(n94588), .B1(n97203), .B2(n109942), .ZN(
        n97217) );
  OAI21_X1 U85319 ( .B1(n81398), .B2(n105367), .A(n97218), .ZN(
        \DLX_Datapath/RegisterFile/N24155 ) );
  AOI22_X1 U85320 ( .A1(n97202), .A2(n94590), .B1(n97203), .B2(n109825), .ZN(
        n97218) );
  OAI21_X1 U85321 ( .B1(n106230), .B2(n105367), .A(n97219), .ZN(
        \DLX_Datapath/RegisterFile/N24154 ) );
  AOI22_X1 U85322 ( .A1(n97202), .A2(n94592), .B1(n97203), .B2(n108199), .ZN(
        n97219) );
  OAI21_X1 U85323 ( .B1(n106171), .B2(n105367), .A(n97220), .ZN(
        \DLX_Datapath/RegisterFile/N24153 ) );
  AOI22_X1 U85324 ( .A1(n97202), .A2(n94594), .B1(n97203), .B2(n108322), .ZN(
        n97220) );
  OAI21_X1 U85325 ( .B1(n81281), .B2(n105367), .A(n97221), .ZN(
        \DLX_Datapath/RegisterFile/N24152 ) );
  AOI22_X1 U85326 ( .A1(n97202), .A2(n94596), .B1(n97203), .B2(n108433), .ZN(
        n97221) );
  OAI21_X1 U85327 ( .B1(n106072), .B2(n105367), .A(n97222), .ZN(
        \DLX_Datapath/RegisterFile/N24151 ) );
  AOI22_X1 U85328 ( .A1(n97202), .A2(n94598), .B1(n97203), .B2(n107671), .ZN(
        n97222) );
  OAI21_X1 U85329 ( .B1(n106198), .B2(n105367), .A(n97223), .ZN(
        \DLX_Datapath/RegisterFile/N24150 ) );
  AOI22_X1 U85330 ( .A1(n97202), .A2(n94600), .B1(n97203), .B2(n109589), .ZN(
        n97223) );
  OAI21_X1 U85331 ( .B1(n106245), .B2(n105367), .A(n97224), .ZN(
        \DLX_Datapath/RegisterFile/N24149 ) );
  AOI22_X1 U85332 ( .A1(n97202), .A2(n94602), .B1(n97203), .B2(n108550), .ZN(
        n97224) );
  OAI21_X1 U85333 ( .B1(n106158), .B2(n105367), .A(n97225), .ZN(
        \DLX_Datapath/RegisterFile/N24148 ) );
  AOI22_X1 U85334 ( .A1(n97202), .A2(n94604), .B1(n97203), .B2(n109694), .ZN(
        n97225) );
  OAI21_X1 U85335 ( .B1(n81394), .B2(n105367), .A(n97226), .ZN(
        \DLX_Datapath/RegisterFile/N24147 ) );
  AOI22_X1 U85336 ( .A1(n97202), .A2(n94606), .B1(n97203), .B2(n109478), .ZN(
        n97226) );
  OAI21_X1 U85337 ( .B1(n106009), .B2(n105367), .A(n97227), .ZN(
        \DLX_Datapath/RegisterFile/N24146 ) );
  AOI22_X1 U85338 ( .A1(n97202), .A2(n94608), .B1(n97203), .B2(n109015), .ZN(
        n97227) );
  OAI21_X1 U85339 ( .B1(n106260), .B2(n105367), .A(n97228), .ZN(
        \DLX_Datapath/RegisterFile/N24145 ) );
  AOI22_X1 U85340 ( .A1(n97202), .A2(n94610), .B1(n97203), .B2(n109363), .ZN(
        n97228) );
  OAI21_X1 U85341 ( .B1(n106044), .B2(n105367), .A(n97229), .ZN(
        \DLX_Datapath/RegisterFile/N24144 ) );
  AOI22_X1 U85342 ( .A1(n97202), .A2(n94612), .B1(n97203), .B2(n109245), .ZN(
        n97229) );
  OAI21_X1 U85343 ( .B1(n106050), .B2(n105367), .A(n97230), .ZN(
        \DLX_Datapath/RegisterFile/N24143 ) );
  AOI22_X1 U85344 ( .A1(n97202), .A2(n94614), .B1(n97203), .B2(n109137), .ZN(
        n97230) );
  OAI21_X1 U85345 ( .B1(n106094), .B2(n105367), .A(n97231), .ZN(
        \DLX_Datapath/RegisterFile/N24142 ) );
  AOI22_X1 U85346 ( .A1(n97202), .A2(n94616), .B1(n97203), .B2(n108672), .ZN(
        n97231) );
  OAI21_X1 U85347 ( .B1(n106053), .B2(n105367), .A(n97232), .ZN(
        \DLX_Datapath/RegisterFile/N24141 ) );
  AOI22_X1 U85348 ( .A1(n97202), .A2(n94618), .B1(n97203), .B2(n108899), .ZN(
        n97232) );
  OAI21_X1 U85349 ( .B1(n105218), .B2(n105367), .A(n97233), .ZN(
        \DLX_Datapath/RegisterFile/N24140 ) );
  AOI22_X1 U85350 ( .A1(n97202), .A2(n94620), .B1(n97203), .B2(n108787), .ZN(
        n97233) );
  OAI21_X1 U85351 ( .B1(n106267), .B2(n105367), .A(n97234), .ZN(
        \DLX_Datapath/RegisterFile/N24139 ) );
  AOI22_X1 U85352 ( .A1(n97202), .A2(n94622), .B1(n97203), .B2(n107327), .ZN(
        n97234) );
  AND2_X2 U85353 ( .A1(n97235), .A2(n97236), .ZN(n97203) );
  AND2_X2 U85354 ( .A1(n97237), .A2(n97236), .ZN(n97202) );
  OR2_X1 U85355 ( .A1(n97200), .A2(n105091), .ZN(n97236) );
  NAND2_X1 U85356 ( .A1(n94434), .A2(n105127), .ZN(n97200) );
  OAI21_X1 U85357 ( .B1(n81358), .B2(n106058), .A(n97238), .ZN(
        \DLX_Datapath/RegisterFile/N24138 ) );
  AOI22_X1 U85358 ( .A1(n81495), .A2(n107890), .B1(n81521), .B2(n104777), .ZN(
        n97238) );
  OAI21_X1 U85359 ( .B1(n106058), .B2(n81651), .A(n97239), .ZN(
        \DLX_Datapath/RegisterFile/N24137 ) );
  AOI22_X1 U85360 ( .A1(n81495), .A2(n107985), .B1(n81653), .B2(n104777), .ZN(
        n97239) );
  OAI21_X1 U85361 ( .B1(n81378), .B2(n106058), .A(n97240), .ZN(
        \DLX_Datapath/RegisterFile/N24136 ) );
  AOI22_X1 U85362 ( .A1(n81495), .A2(n107253), .B1(n104777), .B2(n81380), .ZN(
        n97240) );
  OAI21_X1 U85363 ( .B1(n106208), .B2(n106058), .A(n97241), .ZN(
        \DLX_Datapath/RegisterFile/N24135 ) );
  AOI22_X1 U85364 ( .A1(n81495), .A2(n107792), .B1(n104777), .B2(n81377), .ZN(
        n97241) );
  OAI21_X1 U85365 ( .B1(n106203), .B2(n106058), .A(n97242), .ZN(
        \DLX_Datapath/RegisterFile/N24134 ) );
  AOI22_X1 U85366 ( .A1(n81495), .A2(n110692), .B1(n81496), .B2(n81428), .ZN(
        n97242) );
  OAI21_X1 U85367 ( .B1(n106098), .B2(n106058), .A(n97243), .ZN(
        \DLX_Datapath/RegisterFile/N24133 ) );
  AOI22_X1 U85368 ( .A1(n81495), .A2(n108092), .B1(n104777), .B2(n81410), .ZN(
        n97243) );
  OAI21_X1 U85369 ( .B1(n81270), .B2(n106058), .A(n97244), .ZN(
        \DLX_Datapath/RegisterFile/N24132 ) );
  AOI22_X1 U85370 ( .A1(n81495), .A2(n110791), .B1(n81700), .B2(n81496), .ZN(
        n97244) );
  OAI21_X1 U85371 ( .B1(n81493), .B2(n105990), .A(n97245), .ZN(
        \DLX_Datapath/RegisterFile/N24131 ) );
  AOI22_X1 U85372 ( .A1(n81495), .A2(n110891), .B1(n81632), .B2(n81496), .ZN(
        n97245) );
  OAI21_X1 U85373 ( .B1(n106332), .B2(n106058), .A(n97246), .ZN(
        \DLX_Datapath/RegisterFile/N24130 ) );
  AOI22_X1 U85374 ( .A1(n81495), .A2(n110485), .B1(n81496), .B2(n81414), .ZN(
        n97246) );
  OAI21_X1 U85375 ( .B1(n106190), .B2(n106058), .A(n97247), .ZN(
        \DLX_Datapath/RegisterFile/N24129 ) );
  AOI22_X1 U85376 ( .A1(n81495), .A2(n110267), .B1(n81496), .B2(n81317), .ZN(
        n97247) );
  OAI21_X1 U85377 ( .B1(n106130), .B2(n106058), .A(n97248), .ZN(
        \DLX_Datapath/RegisterFile/N24128 ) );
  AOI22_X1 U85378 ( .A1(n81495), .A2(n110585), .B1(n81496), .B2(n81386), .ZN(
        n97248) );
  OAI21_X1 U85379 ( .B1(n106185), .B2(n81493), .A(n97249), .ZN(
        \DLX_Datapath/RegisterFile/N24127 ) );
  AOI22_X1 U85380 ( .A1(n81495), .A2(n110376), .B1(n104777), .B2(n81320), .ZN(
        n97249) );
  OAI21_X1 U85381 ( .B1(n106163), .B2(n81493), .A(n97250), .ZN(
        \DLX_Datapath/RegisterFile/N24126 ) );
  AOI22_X1 U85382 ( .A1(n81495), .A2(n110052), .B1(n81604), .B2(n104777), .ZN(
        n97250) );
  OAI21_X1 U85383 ( .B1(n106105), .B2(n106058), .A(n97251), .ZN(
        \DLX_Datapath/RegisterFile/N24125 ) );
  AOI22_X1 U85384 ( .A1(n81495), .A2(n110159), .B1(n104777), .B2(n81405), .ZN(
        n97251) );
  OAI21_X1 U85385 ( .B1(n106218), .B2(n106058), .A(n97252), .ZN(
        \DLX_Datapath/RegisterFile/N24124 ) );
  AOI22_X1 U85386 ( .A1(n81495), .A2(n109943), .B1(n81496), .B2(n81402), .ZN(
        n97252) );
  OAI21_X1 U85387 ( .B1(n81398), .B2(n106058), .A(n97253), .ZN(
        \DLX_Datapath/RegisterFile/N24123 ) );
  AOI22_X1 U85388 ( .A1(n81495), .A2(n109826), .B1(n104777), .B2(n81400), .ZN(
        n97253) );
  OAI21_X1 U85389 ( .B1(n106198), .B2(n106058), .A(n97254), .ZN(
        \DLX_Datapath/RegisterFile/N24118 ) );
  AOI22_X1 U85390 ( .A1(n81495), .A2(n109590), .B1(n104777), .B2(n81313), .ZN(
        n97254) );
  OAI21_X1 U85391 ( .B1(n106160), .B2(n106058), .A(n97255), .ZN(
        \DLX_Datapath/RegisterFile/N24116 ) );
  AOI22_X1 U85392 ( .A1(n81495), .A2(n109695), .B1(n104777), .B2(n81425), .ZN(
        n97255) );
  OAI21_X1 U85393 ( .B1(n81394), .B2(n106058), .A(n97256), .ZN(
        \DLX_Datapath/RegisterFile/N24115 ) );
  AOI22_X1 U85394 ( .A1(n81495), .A2(n109479), .B1(n104777), .B2(n81396), .ZN(
        n97256) );
  OAI21_X1 U85395 ( .B1(n106009), .B2(n106058), .A(n97257), .ZN(
        \DLX_Datapath/RegisterFile/N24114 ) );
  AOI22_X1 U85396 ( .A1(n81495), .A2(n109016), .B1(n81590), .B2(n104777), .ZN(
        n97257) );
  OAI21_X1 U85397 ( .B1(n106094), .B2(n106058), .A(n97258), .ZN(
        \DLX_Datapath/RegisterFile/N24110 ) );
  AOI22_X1 U85398 ( .A1(n81495), .A2(n108673), .B1(n81496), .B2(n81417), .ZN(
        n97258) );
  OAI21_X1 U85399 ( .B1(n106266), .B2(n106058), .A(n97259), .ZN(
        \DLX_Datapath/RegisterFile/N24107 ) );
  AOI22_X1 U85400 ( .A1(n81495), .A2(n107328), .B1(n81496), .B2(n81327), .ZN(
        n97259) );
  AND2_X2 U85401 ( .A1(n97237), .A2(n97260), .ZN(n81496) );
  AND2_X2 U85402 ( .A1(n97235), .A2(n97260), .ZN(n81495) );
  OR2_X1 U85403 ( .A1(n81493), .A2(n105095), .ZN(n97260) );
  NAND2_X1 U85404 ( .A1(n105127), .A2(n95132), .ZN(n81493) );
  OAI21_X1 U85405 ( .B1(n81358), .B2(n105366), .A(n97262), .ZN(
        \DLX_Datapath/RegisterFile/N24106 ) );
  AOI22_X1 U85406 ( .A1(n97263), .A2(n94667), .B1(n104731), .B2(n70346), .ZN(
        n97262) );
  OAI21_X1 U85407 ( .B1(n105971), .B2(n97261), .A(n97265), .ZN(
        \DLX_Datapath/RegisterFile/N24105 ) );
  AOI22_X1 U85408 ( .A1(n97263), .A2(n94670), .B1(n97264), .B2(n70488), .ZN(
        n97265) );
  OAI21_X1 U85409 ( .B1(n81378), .B2(n105366), .A(n97266), .ZN(
        \DLX_Datapath/RegisterFile/N24104 ) );
  AOI22_X1 U85410 ( .A1(n97263), .A2(n94672), .B1(n104731), .B2(n69541), .ZN(
        n97266) );
  OAI21_X1 U85411 ( .B1(n106208), .B2(n97261), .A(n97267), .ZN(
        \DLX_Datapath/RegisterFile/N24103 ) );
  AOI22_X1 U85412 ( .A1(n97263), .A2(n94674), .B1(n97264), .B2(n70202), .ZN(
        n97267) );
  OAI21_X1 U85413 ( .B1(n81306), .B2(n105366), .A(n97268), .ZN(
        \DLX_Datapath/RegisterFile/N24102 ) );
  AOI22_X1 U85414 ( .A1(n97263), .A2(n94676), .B1(n104731), .B2(n74048), .ZN(
        n97268) );
  OAI21_X1 U85415 ( .B1(n106100), .B2(n97261), .A(n97269), .ZN(
        \DLX_Datapath/RegisterFile/N24101 ) );
  AOI22_X1 U85416 ( .A1(n97263), .A2(n94678), .B1(n97264), .B2(n70635), .ZN(
        n97269) );
  OAI21_X1 U85417 ( .B1(n81270), .B2(n105366), .A(n97270), .ZN(
        \DLX_Datapath/RegisterFile/N24100 ) );
  AOI22_X1 U85418 ( .A1(n97263), .A2(n94680), .B1(n104731), .B2(n74189), .ZN(
        n97270) );
  OAI21_X1 U85419 ( .B1(n105991), .B2(n105366), .A(n97271), .ZN(
        \DLX_Datapath/RegisterFile/N24099 ) );
  AOI22_X1 U85420 ( .A1(n97263), .A2(n94682), .B1(n97264), .B2(n74329), .ZN(
        n97271) );
  OAI21_X1 U85421 ( .B1(n106332), .B2(n97261), .A(n97272), .ZN(
        \DLX_Datapath/RegisterFile/N24098 ) );
  AOI22_X1 U85422 ( .A1(n97263), .A2(n94684), .B1(n97264), .B2(n73765), .ZN(
        n97272) );
  OAI21_X1 U85423 ( .B1(n106191), .B2(n97261), .A(n97273), .ZN(
        \DLX_Datapath/RegisterFile/N24097 ) );
  AOI22_X1 U85424 ( .A1(n97263), .A2(n94686), .B1(n104731), .B2(n73469), .ZN(
        n97273) );
  OAI21_X1 U85425 ( .B1(n106130), .B2(n97261), .A(n97274), .ZN(
        \DLX_Datapath/RegisterFile/N24096 ) );
  AOI22_X1 U85426 ( .A1(n97263), .A2(n94688), .B1(n97264), .B2(n73906), .ZN(
        n97274) );
  OAI21_X1 U85427 ( .B1(n106187), .B2(n105366), .A(n97275), .ZN(
        \DLX_Datapath/RegisterFile/N24095 ) );
  AOI22_X1 U85428 ( .A1(n97263), .A2(n94690), .B1(n104731), .B2(n73618), .ZN(
        n97275) );
  OAI21_X1 U85429 ( .B1(n106163), .B2(n105366), .A(n97276), .ZN(
        \DLX_Datapath/RegisterFile/N24094 ) );
  AOI22_X1 U85430 ( .A1(n97263), .A2(n94692), .B1(n97264), .B2(n73180), .ZN(
        n97276) );
  OAI21_X1 U85431 ( .B1(n106104), .B2(n105366), .A(n97277), .ZN(
        \DLX_Datapath/RegisterFile/N24093 ) );
  AOI22_X1 U85432 ( .A1(n97263), .A2(n94694), .B1(n104731), .B2(n73322), .ZN(
        n97277) );
  OAI21_X1 U85433 ( .B1(n106218), .B2(n105366), .A(n97278), .ZN(
        \DLX_Datapath/RegisterFile/N24092 ) );
  AOI22_X1 U85434 ( .A1(n97263), .A2(n94696), .B1(n104731), .B2(n73038), .ZN(
        n97278) );
  OAI21_X1 U85435 ( .B1(n81398), .B2(n105366), .A(n97279), .ZN(
        \DLX_Datapath/RegisterFile/N24091 ) );
  AOI22_X1 U85436 ( .A1(n97263), .A2(n94698), .B1(n97264), .B2(n72888), .ZN(
        n97279) );
  OAI21_X1 U85437 ( .B1(n106233), .B2(n105366), .A(n97280), .ZN(
        \DLX_Datapath/RegisterFile/N24090 ) );
  AOI22_X1 U85438 ( .A1(n97263), .A2(n94700), .B1(n104731), .B2(n70784), .ZN(
        n97280) );
  OAI21_X1 U85439 ( .B1(n106172), .B2(n105366), .A(n97281), .ZN(
        \DLX_Datapath/RegisterFile/N24089 ) );
  AOI22_X1 U85440 ( .A1(n97263), .A2(n94702), .B1(n97264), .B2(n70943), .ZN(
        n97281) );
  OAI21_X1 U85441 ( .B1(n81281), .B2(n105366), .A(n97282), .ZN(
        \DLX_Datapath/RegisterFile/N24088 ) );
  AOI22_X1 U85442 ( .A1(n97263), .A2(n94704), .B1(n97264), .B2(n71088), .ZN(
        n97282) );
  OAI21_X1 U85443 ( .B1(n106071), .B2(n105366), .A(n97283), .ZN(
        \DLX_Datapath/RegisterFile/N24087 ) );
  AOI22_X1 U85444 ( .A1(n97263), .A2(n94706), .B1(n104731), .B2(n70049), .ZN(
        n97283) );
  OAI21_X1 U85445 ( .B1(n106198), .B2(n105366), .A(n97284), .ZN(
        \DLX_Datapath/RegisterFile/N24086 ) );
  AOI22_X1 U85446 ( .A1(n97263), .A2(n94708), .B1(n97264), .B2(n72578), .ZN(
        n97284) );
  OAI21_X1 U85447 ( .B1(n106245), .B2(n105366), .A(n97285), .ZN(
        \DLX_Datapath/RegisterFile/N24085 ) );
  AOI22_X1 U85448 ( .A1(n97263), .A2(n94710), .B1(n104731), .B2(n71237), .ZN(
        n97285) );
  OAI21_X1 U85449 ( .B1(n106159), .B2(n105366), .A(n97286), .ZN(
        \DLX_Datapath/RegisterFile/N24084 ) );
  AOI22_X1 U85450 ( .A1(n97263), .A2(n94712), .B1(n104731), .B2(n72720), .ZN(
        n97286) );
  OAI21_X1 U85451 ( .B1(n81394), .B2(n105366), .A(n97287), .ZN(
        \DLX_Datapath/RegisterFile/N24083 ) );
  AOI22_X1 U85452 ( .A1(n97263), .A2(n94714), .B1(n97264), .B2(n72430), .ZN(
        n97287) );
  OAI21_X1 U85453 ( .B1(n106009), .B2(n105366), .A(n97288), .ZN(
        \DLX_Datapath/RegisterFile/N24082 ) );
  AOI22_X1 U85454 ( .A1(n97263), .A2(n81259), .B1(n104731), .B2(n71830), .ZN(
        n97288) );
  OAI21_X1 U85455 ( .B1(n106260), .B2(n105366), .A(n97289), .ZN(
        \DLX_Datapath/RegisterFile/N24081 ) );
  AOI22_X1 U85456 ( .A1(n97263), .A2(n94717), .B1(n104731), .B2(n72279), .ZN(
        n97289) );
  OAI21_X1 U85457 ( .B1(n106044), .B2(n105366), .A(n97290), .ZN(
        \DLX_Datapath/RegisterFile/N24080 ) );
  AOI22_X1 U85458 ( .A1(n97263), .A2(n94719), .B1(n97264), .B2(n72128), .ZN(
        n97290) );
  OAI21_X1 U85459 ( .B1(n106049), .B2(n105366), .A(n97291), .ZN(
        \DLX_Datapath/RegisterFile/N24079 ) );
  AOI22_X1 U85460 ( .A1(n97263), .A2(n94721), .B1(n104731), .B2(n71984), .ZN(
        n97291) );
  OAI21_X1 U85461 ( .B1(n106094), .B2(n105366), .A(n97292), .ZN(
        \DLX_Datapath/RegisterFile/N24078 ) );
  AOI22_X1 U85462 ( .A1(n97263), .A2(n94723), .B1(n97264), .B2(n71386), .ZN(
        n97292) );
  OAI21_X1 U85463 ( .B1(n106054), .B2(n105366), .A(n97293), .ZN(
        \DLX_Datapath/RegisterFile/N24077 ) );
  AOI22_X1 U85464 ( .A1(n97263), .A2(n94725), .B1(n97264), .B2(n71681), .ZN(
        n97293) );
  OAI21_X1 U85465 ( .B1(n105217), .B2(n105366), .A(n97294), .ZN(
        \DLX_Datapath/RegisterFile/N24076 ) );
  AOI22_X1 U85466 ( .A1(n97263), .A2(n94727), .B1(n97264), .B2(n71537), .ZN(
        n97294) );
  OAI21_X1 U85467 ( .B1(n106267), .B2(n105366), .A(n97295), .ZN(
        \DLX_Datapath/RegisterFile/N24075 ) );
  AOI22_X1 U85468 ( .A1(n97263), .A2(n94729), .B1(n104731), .B2(n69646), .ZN(
        n97295) );
  AND2_X2 U85469 ( .A1(n97235), .A2(n97296), .ZN(n97264) );
  OAI21_X1 U85470 ( .B1(n94366), .B2(n97237), .A(n105602), .ZN(n97235) );
  AND2_X2 U85471 ( .A1(n97237), .A2(n97296), .ZN(n97263) );
  OR2_X1 U85472 ( .A1(n97261), .A2(n105089), .ZN(n97296) );
  NOR2_X1 U85473 ( .A1(n97061), .A2(n95131), .ZN(n97237) );
  NAND2_X1 U85474 ( .A1(n105127), .A2(n94505), .ZN(n97261) );
  OAI21_X1 U85475 ( .B1(n106078), .B2(n105970), .A(n97297), .ZN(
        \DLX_Datapath/RegisterFile/N24073 ) );
  AOI22_X1 U85476 ( .A1(n81445), .A2(n107986), .B1(n94511), .B2(n106074), .ZN(
        n97297) );
  OAI21_X1 U85477 ( .B1(n106135), .B2(n106078), .A(n97298), .ZN(
        \DLX_Datapath/RegisterFile/N24072 ) );
  AOI22_X1 U85478 ( .A1(n81445), .A2(n107254), .B1(n81539), .B2(n81446), .ZN(
        n97298) );
  OAI21_X1 U85479 ( .B1(n106209), .B2(n106078), .A(n97299), .ZN(
        \DLX_Datapath/RegisterFile/N24071 ) );
  AOI22_X1 U85480 ( .A1(n81445), .A2(n107793), .B1(n106074), .B2(n81301), .ZN(
        n97299) );
  OAI21_X1 U85481 ( .B1(n106098), .B2(n106078), .A(n97300), .ZN(
        \DLX_Datapath/RegisterFile/N24069 ) );
  AOI22_X1 U85482 ( .A1(n81445), .A2(n108093), .B1(n94516), .B2(n81446), .ZN(
        n97300) );
  OAI21_X1 U85483 ( .B1(n106079), .B2(n81629), .A(n97301), .ZN(
        \DLX_Datapath/RegisterFile/N24067 ) );
  AOI22_X1 U85484 ( .A1(n106077), .A2(n111016), .B1(n94519), .B2(n106075), 
        .ZN(n97301) );
  OAI21_X1 U85485 ( .B1(n106331), .B2(n106078), .A(n97302), .ZN(
        \DLX_Datapath/RegisterFile/N24066 ) );
  AOI22_X1 U85486 ( .A1(n81445), .A2(n111017), .B1(n106074), .B2(n80192), .ZN(
        n97302) );
  OAI21_X1 U85487 ( .B1(n106191), .B2(n106078), .A(n97303), .ZN(
        \DLX_Datapath/RegisterFile/N24065 ) );
  AOI22_X1 U85488 ( .A1(n81445), .A2(n110268), .B1(n81474), .B2(n81446), .ZN(
        n97303) );
  OAI21_X1 U85489 ( .B1(n106130), .B2(n106078), .A(n97304), .ZN(
        \DLX_Datapath/RegisterFile/N24064 ) );
  AOI22_X1 U85490 ( .A1(n81445), .A2(n110586), .B1(n94523), .B2(n81446), .ZN(
        n97304) );
  OAI21_X1 U85491 ( .B1(n106186), .B2(n106079), .A(n97305), .ZN(
        \DLX_Datapath/RegisterFile/N24063 ) );
  AOI22_X1 U85492 ( .A1(n106076), .A2(n110377), .B1(n106062), .B2(n81446), 
        .ZN(n97305) );
  OAI21_X1 U85493 ( .B1(n81403), .B2(n106079), .A(n97306), .ZN(
        \DLX_Datapath/RegisterFile/N24061 ) );
  AOI22_X1 U85494 ( .A1(n106077), .A2(n110160), .B1(n94527), .B2(n106075), 
        .ZN(n97306) );
  OAI21_X1 U85495 ( .B1(n106218), .B2(n106079), .A(n97307), .ZN(
        \DLX_Datapath/RegisterFile/N24060 ) );
  AOI22_X1 U85496 ( .A1(n106076), .A2(n109944), .B1(n106074), .B2(n81297), 
        .ZN(n97307) );
  OAI21_X1 U85497 ( .B1(n81398), .B2(n106079), .A(n97308), .ZN(
        \DLX_Datapath/RegisterFile/N24059 ) );
  AOI22_X1 U85498 ( .A1(n106077), .A2(n109827), .B1(n94530), .B2(n106075), 
        .ZN(n97308) );
  OAI21_X1 U85499 ( .B1(n106198), .B2(n106079), .A(n97309), .ZN(
        \DLX_Datapath/RegisterFile/N24054 ) );
  AOI22_X1 U85500 ( .A1(n106076), .A2(n109591), .B1(n94536), .B2(n81446), .ZN(
        n97309) );
  OAI21_X1 U85501 ( .B1(n106157), .B2(n106079), .A(n97310), .ZN(
        \DLX_Datapath/RegisterFile/N24052 ) );
  AOI22_X1 U85502 ( .A1(n106077), .A2(n109696), .B1(n106074), .B2(n81351), 
        .ZN(n97310) );
  OAI21_X1 U85503 ( .B1(n106114), .B2(n106079), .A(n97311), .ZN(
        \DLX_Datapath/RegisterFile/N24051 ) );
  AOI22_X1 U85504 ( .A1(n106076), .A2(n109480), .B1(n106021), .B2(n81446), 
        .ZN(n97311) );
  OAI21_X1 U85505 ( .B1(n106009), .B2(n106079), .A(n97312), .ZN(
        \DLX_Datapath/RegisterFile/N24050 ) );
  AOI22_X1 U85506 ( .A1(n106077), .A2(n109017), .B1(n94541), .B2(n106074), 
        .ZN(n97312) );
  OAI21_X1 U85507 ( .B1(n106079), .B2(n81509), .A(n97313), .ZN(
        \DLX_Datapath/RegisterFile/N24048 ) );
  AOI22_X1 U85508 ( .A1(n106076), .A2(n109247), .B1(n105624), .B2(n106074), 
        .ZN(n97313) );
  OAI21_X1 U85509 ( .B1(n106078), .B2(n106051), .A(n97314), .ZN(
        \DLX_Datapath/RegisterFile/N24047 ) );
  AOI22_X1 U85510 ( .A1(n106076), .A2(n109139), .B1(n94546), .B2(n106074), 
        .ZN(n97314) );
  OAI21_X1 U85511 ( .B1(n106094), .B2(n106079), .A(n97315), .ZN(
        \DLX_Datapath/RegisterFile/N24046 ) );
  AOI22_X1 U85512 ( .A1(n106076), .A2(n108674), .B1(n94548), .B2(n106074), 
        .ZN(n97315) );
  OAI21_X1 U85513 ( .B1(n106078), .B2(n81498), .A(n97316), .ZN(
        \DLX_Datapath/RegisterFile/N24045 ) );
  AOI22_X1 U85514 ( .A1(n106077), .A2(n108901), .B1(n81783), .B2(n106074), 
        .ZN(n97316) );
  OAI21_X1 U85515 ( .B1(n106266), .B2(n106079), .A(n97317), .ZN(
        \DLX_Datapath/RegisterFile/N24043 ) );
  AOI22_X1 U85516 ( .A1(n106077), .A2(n107329), .B1(n106075), .B2(n81265), 
        .ZN(n97317) );
  NOR2_X1 U85517 ( .A1(n97318), .A2(n104692), .ZN(n81446) );
  AOI21_X1 U85518 ( .B1(n97058), .B2(n94554), .A(n104692), .ZN(n81445) );
  NAND2_X1 U85520 ( .A1(n105128), .A2(n94555), .ZN(n81443) );
  OAI21_X1 U85521 ( .B1(n81358), .B2(n105365), .A(n97321), .ZN(
        \DLX_Datapath/RegisterFile/N24042 ) );
  AOI22_X1 U85522 ( .A1(n105363), .A2(n70348), .B1(n105361), .B2(n94559), .ZN(
        n97321) );
  OAI21_X1 U85523 ( .B1(n105969), .B2(n105365), .A(n97324), .ZN(
        \DLX_Datapath/RegisterFile/N24041 ) );
  AOI22_X1 U85524 ( .A1(n105362), .A2(n70490), .B1(n105360), .B2(n94562), .ZN(
        n97324) );
  OAI21_X1 U85525 ( .B1(n81378), .B2(n105365), .A(n97325), .ZN(
        \DLX_Datapath/RegisterFile/N24040 ) );
  AOI22_X1 U85526 ( .A1(n105363), .A2(n69543), .B1(n105361), .B2(n94564), .ZN(
        n97325) );
  OAI21_X1 U85527 ( .B1(n106209), .B2(n105365), .A(n97326), .ZN(
        \DLX_Datapath/RegisterFile/N24039 ) );
  AOI22_X1 U85528 ( .A1(n105362), .A2(n70204), .B1(n105360), .B2(n94566), .ZN(
        n97326) );
  OAI21_X1 U85529 ( .B1(n106204), .B2(n105365), .A(n97327), .ZN(
        \DLX_Datapath/RegisterFile/N24038 ) );
  AOI22_X1 U85530 ( .A1(n105363), .A2(n74050), .B1(n105361), .B2(n94568), .ZN(
        n97327) );
  OAI21_X1 U85531 ( .B1(n106098), .B2(n105365), .A(n97328), .ZN(
        \DLX_Datapath/RegisterFile/N24037 ) );
  AOI22_X1 U85532 ( .A1(n105362), .A2(n70637), .B1(n105360), .B2(n94570), .ZN(
        n97328) );
  OAI21_X1 U85533 ( .B1(n106257), .B2(n105365), .A(n97329), .ZN(
        \DLX_Datapath/RegisterFile/N24036 ) );
  AOI22_X1 U85534 ( .A1(n105363), .A2(n74191), .B1(n105361), .B2(n94572), .ZN(
        n97329) );
  OAI21_X1 U85535 ( .B1(n105990), .B2(n105365), .A(n97330), .ZN(
        \DLX_Datapath/RegisterFile/N24035 ) );
  AOI22_X1 U85536 ( .A1(n105362), .A2(n74331), .B1(n105360), .B2(n94574), .ZN(
        n97330) );
  OAI21_X1 U85537 ( .B1(n106330), .B2(n105365), .A(n97331), .ZN(
        \DLX_Datapath/RegisterFile/N24034 ) );
  AOI22_X1 U85538 ( .A1(n105362), .A2(n73767), .B1(n105360), .B2(n94576), .ZN(
        n97331) );
  OAI21_X1 U85539 ( .B1(n106193), .B2(n105364), .A(n97332), .ZN(
        \DLX_Datapath/RegisterFile/N24033 ) );
  AOI22_X1 U85540 ( .A1(n105362), .A2(n73471), .B1(n97323), .B2(n94578), .ZN(
        n97332) );
  OAI21_X1 U85541 ( .B1(n106130), .B2(n105364), .A(n97333), .ZN(
        \DLX_Datapath/RegisterFile/N24032 ) );
  AOI22_X1 U85542 ( .A1(n97322), .A2(n73908), .B1(n97323), .B2(n94580), .ZN(
        n97333) );
  OAI21_X1 U85543 ( .B1(n106186), .B2(n105364), .A(n97334), .ZN(
        \DLX_Datapath/RegisterFile/N24031 ) );
  AOI22_X1 U85544 ( .A1(n97322), .A2(n73620), .B1(n97323), .B2(n94582), .ZN(
        n97334) );
  OAI21_X1 U85545 ( .B1(n106163), .B2(n105364), .A(n97335), .ZN(
        \DLX_Datapath/RegisterFile/N24030 ) );
  AOI22_X1 U85546 ( .A1(n97322), .A2(n73182), .B1(n97323), .B2(n94584), .ZN(
        n97335) );
  OAI21_X1 U85547 ( .B1(n81403), .B2(n105364), .A(n97336), .ZN(
        \DLX_Datapath/RegisterFile/N24029 ) );
  AOI22_X1 U85548 ( .A1(n105362), .A2(n73324), .B1(n105361), .B2(n94586), .ZN(
        n97336) );
  OAI21_X1 U85549 ( .B1(n106218), .B2(n105364), .A(n97337), .ZN(
        \DLX_Datapath/RegisterFile/N24028 ) );
  AOI22_X1 U85550 ( .A1(n97322), .A2(n73040), .B1(n97323), .B2(n94588), .ZN(
        n97337) );
  OAI21_X1 U85551 ( .B1(n81398), .B2(n105364), .A(n97338), .ZN(
        \DLX_Datapath/RegisterFile/N24027 ) );
  AOI22_X1 U85552 ( .A1(n105362), .A2(n72890), .B1(n105361), .B2(n94590), .ZN(
        n97338) );
  OAI21_X1 U85553 ( .B1(n106232), .B2(n105364), .A(n97339), .ZN(
        \DLX_Datapath/RegisterFile/N24026 ) );
  AOI22_X1 U85554 ( .A1(n97322), .A2(n70786), .B1(n97323), .B2(n94592), .ZN(
        n97339) );
  OAI21_X1 U85555 ( .B1(n106172), .B2(n105364), .A(n97340), .ZN(
        \DLX_Datapath/RegisterFile/N24025 ) );
  AOI22_X1 U85556 ( .A1(n97322), .A2(n70945), .B1(n97323), .B2(n94594), .ZN(
        n97340) );
  OAI21_X1 U85557 ( .B1(n81281), .B2(n105364), .A(n97341), .ZN(
        \DLX_Datapath/RegisterFile/N24024 ) );
  AOI22_X1 U85558 ( .A1(n105363), .A2(n71090), .B1(n105360), .B2(n94596), .ZN(
        n97341) );
  OAI21_X1 U85559 ( .B1(n106069), .B2(n105364), .A(n97342), .ZN(
        \DLX_Datapath/RegisterFile/N24023 ) );
  AOI22_X1 U85560 ( .A1(n97322), .A2(n70051), .B1(n97323), .B2(n94598), .ZN(
        n97342) );
  OAI21_X1 U85561 ( .B1(n106199), .B2(n105364), .A(n97343), .ZN(
        \DLX_Datapath/RegisterFile/N24022 ) );
  AOI22_X1 U85562 ( .A1(n105362), .A2(n72580), .B1(n105360), .B2(n94600), .ZN(
        n97343) );
  OAI21_X1 U85563 ( .B1(n106245), .B2(n105365), .A(n97344), .ZN(
        \DLX_Datapath/RegisterFile/N24021 ) );
  AOI22_X1 U85564 ( .A1(n105363), .A2(n71239), .B1(n105361), .B2(n94602), .ZN(
        n97344) );
  OAI21_X1 U85565 ( .B1(n106158), .B2(n105365), .A(n97345), .ZN(
        \DLX_Datapath/RegisterFile/N24020 ) );
  AOI22_X1 U85566 ( .A1(n105362), .A2(n72722), .B1(n105360), .B2(n94604), .ZN(
        n97345) );
  OAI21_X1 U85567 ( .B1(n81394), .B2(n105364), .A(n97346), .ZN(
        \DLX_Datapath/RegisterFile/N24019 ) );
  AOI22_X1 U85568 ( .A1(n105363), .A2(n72432), .B1(n105361), .B2(n94606), .ZN(
        n97346) );
  OAI21_X1 U85569 ( .B1(n106009), .B2(n105365), .A(n97347), .ZN(
        \DLX_Datapath/RegisterFile/N24018 ) );
  AOI22_X1 U85570 ( .A1(n105362), .A2(n71832), .B1(n105360), .B2(n94608), .ZN(
        n97347) );
  OAI21_X1 U85571 ( .B1(n106260), .B2(n105365), .A(n97348), .ZN(
        \DLX_Datapath/RegisterFile/N24017 ) );
  AOI22_X1 U85572 ( .A1(n105363), .A2(n72281), .B1(n105361), .B2(n94610), .ZN(
        n97348) );
  OAI21_X1 U85573 ( .B1(n106044), .B2(n105364), .A(n97349), .ZN(
        \DLX_Datapath/RegisterFile/N24016 ) );
  AOI22_X1 U85574 ( .A1(n105362), .A2(n72130), .B1(n105360), .B2(n94612), .ZN(
        n97349) );
  OAI21_X1 U85575 ( .B1(n106050), .B2(n105365), .A(n97350), .ZN(
        \DLX_Datapath/RegisterFile/N24015 ) );
  AOI22_X1 U85576 ( .A1(n105363), .A2(n71986), .B1(n105361), .B2(n94614), .ZN(
        n97350) );
  OAI21_X1 U85577 ( .B1(n106094), .B2(n105364), .A(n97351), .ZN(
        \DLX_Datapath/RegisterFile/N24014 ) );
  AOI22_X1 U85578 ( .A1(n105362), .A2(n71388), .B1(n105360), .B2(n94616), .ZN(
        n97351) );
  OAI21_X1 U85579 ( .B1(n106056), .B2(n105365), .A(n97352), .ZN(
        \DLX_Datapath/RegisterFile/N24013 ) );
  AOI22_X1 U85580 ( .A1(n105363), .A2(n71683), .B1(n105361), .B2(n94618), .ZN(
        n97352) );
  OAI21_X1 U85581 ( .B1(n105217), .B2(n105365), .A(n97353), .ZN(
        \DLX_Datapath/RegisterFile/N24012 ) );
  AOI22_X1 U85582 ( .A1(n105363), .A2(n71539), .B1(n105361), .B2(n94620), .ZN(
        n97353) );
  OAI21_X1 U85583 ( .B1(n106268), .B2(n105364), .A(n97354), .ZN(
        \DLX_Datapath/RegisterFile/N24011 ) );
  AOI22_X1 U85584 ( .A1(n105362), .A2(n69648), .B1(n105360), .B2(n94622), .ZN(
        n97354) );
  NOR2_X1 U85585 ( .A1(n97318), .A2(n97355), .ZN(n97323) );
  NOR2_X1 U85586 ( .A1(n97356), .A2(n97355), .ZN(n97322) );
  NOR2_X1 U85587 ( .A1(n97320), .A2(n105094), .ZN(n97355) );
  NAND2_X1 U85588 ( .A1(n94625), .A2(n105128), .ZN(n97320) );
  OAI21_X1 U85589 ( .B1(n106148), .B2(n105359), .A(n97358), .ZN(
        \DLX_Datapath/RegisterFile/N24010 ) );
  AOI22_X1 U85590 ( .A1(n104864), .A2(n81521), .B1(n105357), .B2(n107892), 
        .ZN(n97358) );
  OAI21_X1 U85591 ( .B1(n105971), .B2(n105359), .A(n97361), .ZN(
        \DLX_Datapath/RegisterFile/N24009 ) );
  AOI22_X1 U85592 ( .A1(n104864), .A2(n81653), .B1(n105357), .B2(n107987), 
        .ZN(n97361) );
  OAI21_X1 U85593 ( .B1(n81378), .B2(n105359), .A(n97362), .ZN(
        \DLX_Datapath/RegisterFile/N24008 ) );
  AOI22_X1 U85594 ( .A1(n104863), .A2(n81380), .B1(n105357), .B2(n107255), 
        .ZN(n97362) );
  OAI21_X1 U85595 ( .B1(n106209), .B2(n105359), .A(n97363), .ZN(
        \DLX_Datapath/RegisterFile/N24007 ) );
  AOI22_X1 U85596 ( .A1(n104863), .A2(n81377), .B1(n105357), .B2(n107794), 
        .ZN(n97363) );
  OAI21_X1 U85597 ( .B1(n106205), .B2(n105359), .A(n97364), .ZN(
        \DLX_Datapath/RegisterFile/N24006 ) );
  AOI22_X1 U85598 ( .A1(n97359), .A2(n81428), .B1(n105357), .B2(n110694), .ZN(
        n97364) );
  OAI21_X1 U85599 ( .B1(n106101), .B2(n105359), .A(n97365), .ZN(
        \DLX_Datapath/RegisterFile/N24005 ) );
  AOI22_X1 U85600 ( .A1(n97359), .A2(n81410), .B1(n105357), .B2(n108094), .ZN(
        n97365) );
  OAI21_X1 U85601 ( .B1(n106255), .B2(n105359), .A(n97366), .ZN(
        \DLX_Datapath/RegisterFile/N24004 ) );
  AOI22_X1 U85602 ( .A1(n104863), .A2(n81700), .B1(n105357), .B2(n110793), 
        .ZN(n97366) );
  OAI21_X1 U85603 ( .B1(n105992), .B2(n105359), .A(n97367), .ZN(
        \DLX_Datapath/RegisterFile/N24003 ) );
  AOI22_X1 U85604 ( .A1(n104863), .A2(n81632), .B1(n105357), .B2(n110892), 
        .ZN(n97367) );
  OAI21_X1 U85605 ( .B1(n106333), .B2(n105359), .A(n97368), .ZN(
        \DLX_Datapath/RegisterFile/N24002 ) );
  AOI22_X1 U85606 ( .A1(n104864), .A2(n81414), .B1(n97360), .B2(n110486), .ZN(
        n97368) );
  OAI21_X1 U85607 ( .B1(n106190), .B2(n105358), .A(n97369), .ZN(
        \DLX_Datapath/RegisterFile/N24001 ) );
  AOI22_X1 U85608 ( .A1(n97359), .A2(n81317), .B1(n97360), .B2(n110269), .ZN(
        n97369) );
  OAI21_X1 U85609 ( .B1(n106128), .B2(n105358), .A(n97370), .ZN(
        \DLX_Datapath/RegisterFile/N24000 ) );
  AOI22_X1 U85610 ( .A1(n104864), .A2(n81386), .B1(n97360), .B2(n110587), .ZN(
        n97370) );
  OAI21_X1 U85611 ( .B1(n106186), .B2(n105358), .A(n97371), .ZN(
        \DLX_Datapath/RegisterFile/N23999 ) );
  AOI22_X1 U85612 ( .A1(n104863), .A2(n81320), .B1(n105357), .B2(n110378), 
        .ZN(n97371) );
  OAI21_X1 U85613 ( .B1(n106163), .B2(n105358), .A(n97372), .ZN(
        \DLX_Datapath/RegisterFile/N23998 ) );
  AOI22_X1 U85614 ( .A1(n104863), .A2(n81604), .B1(n97360), .B2(n110054), .ZN(
        n97372) );
  OAI21_X1 U85615 ( .B1(n81403), .B2(n105358), .A(n97373), .ZN(
        \DLX_Datapath/RegisterFile/N23997 ) );
  AOI22_X1 U85616 ( .A1(n104863), .A2(n81405), .B1(n105357), .B2(n110161), 
        .ZN(n97373) );
  OAI21_X1 U85617 ( .B1(n106219), .B2(n105358), .A(n97374), .ZN(
        \DLX_Datapath/RegisterFile/N23996 ) );
  AOI22_X1 U85618 ( .A1(n97359), .A2(n81402), .B1(n97360), .B2(n109945), .ZN(
        n97374) );
  OAI21_X1 U85619 ( .B1(n81398), .B2(n105358), .A(n97375), .ZN(
        \DLX_Datapath/RegisterFile/N23995 ) );
  AOI22_X1 U85620 ( .A1(n104864), .A2(n81400), .B1(n105357), .B2(n109828), 
        .ZN(n97375) );
  OAI21_X1 U85621 ( .B1(n106231), .B2(n105358), .A(n97376), .ZN(
        \DLX_Datapath/RegisterFile/N23994 ) );
  AOI22_X1 U85622 ( .A1(n104863), .A2(n81332), .B1(n105357), .B2(n108202), 
        .ZN(n97376) );
  OAI21_X1 U85623 ( .B1(n106172), .B2(n105358), .A(n97377), .ZN(
        \DLX_Datapath/RegisterFile/N23993 ) );
  AOI22_X1 U85624 ( .A1(n104864), .A2(n81373), .B1(n105356), .B2(n108325), 
        .ZN(n97377) );
  OAI21_X1 U85625 ( .B1(n81281), .B2(n105358), .A(n97378), .ZN(
        \DLX_Datapath/RegisterFile/N23992 ) );
  AOI22_X1 U85626 ( .A1(n104864), .A2(n81322), .B1(n105357), .B2(n108436), 
        .ZN(n97378) );
  OAI21_X1 U85627 ( .B1(n106070), .B2(n105358), .A(n97379), .ZN(
        \DLX_Datapath/RegisterFile/N23991 ) );
  AOI22_X1 U85628 ( .A1(n104864), .A2(n81506), .B1(n97360), .B2(n107674), .ZN(
        n97379) );
  OAI21_X1 U85629 ( .B1(n106198), .B2(n105358), .A(n97380), .ZN(
        \DLX_Datapath/RegisterFile/N23990 ) );
  AOI22_X1 U85630 ( .A1(n104863), .A2(n81313), .B1(n105356), .B2(n109592), 
        .ZN(n97380) );
  OAI21_X1 U85631 ( .B1(n106245), .B2(n105359), .A(n97381), .ZN(
        \DLX_Datapath/RegisterFile/N23989 ) );
  AOI22_X1 U85632 ( .A1(n104863), .A2(n81330), .B1(n105356), .B2(n108553), 
        .ZN(n97381) );
  OAI21_X1 U85633 ( .B1(n106159), .B2(n105359), .A(n97382), .ZN(
        \DLX_Datapath/RegisterFile/N23988 ) );
  AOI22_X1 U85634 ( .A1(n104863), .A2(n81425), .B1(n105356), .B2(n109697), 
        .ZN(n97382) );
  OAI21_X1 U85635 ( .B1(n81394), .B2(n105358), .A(n97383), .ZN(
        \DLX_Datapath/RegisterFile/N23987 ) );
  AOI22_X1 U85636 ( .A1(n104863), .A2(n81396), .B1(n105356), .B2(n109481), 
        .ZN(n97383) );
  OAI21_X1 U85637 ( .B1(n106009), .B2(n105359), .A(n97384), .ZN(
        \DLX_Datapath/RegisterFile/N23986 ) );
  AOI22_X1 U85638 ( .A1(n97359), .A2(n81590), .B1(n105356), .B2(n109018), .ZN(
        n97384) );
  OAI21_X1 U85639 ( .B1(n106260), .B2(n105359), .A(n97385), .ZN(
        \DLX_Datapath/RegisterFile/N23985 ) );
  AOI22_X1 U85640 ( .A1(n104864), .A2(n81423), .B1(n105356), .B2(n109366), 
        .ZN(n97385) );
  OAI21_X1 U85641 ( .B1(n106044), .B2(n105358), .A(n97386), .ZN(
        \DLX_Datapath/RegisterFile/N23984 ) );
  AOI22_X1 U85642 ( .A1(n104863), .A2(n81511), .B1(n105356), .B2(n109248), 
        .ZN(n97386) );
  OAI21_X1 U85643 ( .B1(n106048), .B2(n105359), .A(n97387), .ZN(
        \DLX_Datapath/RegisterFile/N23983 ) );
  AOI22_X1 U85644 ( .A1(n104864), .A2(n81503), .B1(n105356), .B2(n109140), 
        .ZN(n97387) );
  OAI21_X1 U85645 ( .B1(n106094), .B2(n105358), .A(n97388), .ZN(
        \DLX_Datapath/RegisterFile/N23982 ) );
  AOI22_X1 U85646 ( .A1(n97359), .A2(n81417), .B1(n105356), .B2(n108675), .ZN(
        n97388) );
  OAI21_X1 U85647 ( .B1(n106055), .B2(n105359), .A(n97389), .ZN(
        \DLX_Datapath/RegisterFile/N23981 ) );
  AOI22_X1 U85648 ( .A1(n104864), .A2(n81500), .B1(n105356), .B2(n108902), 
        .ZN(n97389) );
  OAI21_X1 U85649 ( .B1(n105217), .B2(n105359), .A(n97390), .ZN(
        \DLX_Datapath/RegisterFile/N23980 ) );
  AOI22_X1 U85650 ( .A1(n97359), .A2(n81335), .B1(n105356), .B2(n108790), .ZN(
        n97390) );
  OAI21_X1 U85651 ( .B1(n106268), .B2(n105358), .A(n97391), .ZN(
        \DLX_Datapath/RegisterFile/N23979 ) );
  AOI22_X1 U85652 ( .A1(n104863), .A2(n81327), .B1(n105356), .B2(n107330), 
        .ZN(n97391) );
  NOR2_X1 U85653 ( .A1(n97356), .A2(n97392), .ZN(n97360) );
  NOR2_X1 U85654 ( .A1(n97318), .A2(n97392), .ZN(n97359) );
  NOR2_X1 U85655 ( .A1(n97357), .A2(n105089), .ZN(n97392) );
  NAND2_X1 U85656 ( .A1(n105127), .A2(n94664), .ZN(n97357) );
  OAI21_X1 U85657 ( .B1(n106148), .B2(n105355), .A(n97394), .ZN(
        \DLX_Datapath/RegisterFile/N23978 ) );
  AOI22_X1 U85658 ( .A1(n105353), .A2(n94667), .B1(n97396), .B2(n70350), .ZN(
        n97394) );
  OAI21_X1 U85659 ( .B1(n105968), .B2(n105355), .A(n97397), .ZN(
        \DLX_Datapath/RegisterFile/N23977 ) );
  AOI22_X1 U85660 ( .A1(n105353), .A2(n94670), .B1(n105351), .B2(n70492), .ZN(
        n97397) );
  OAI21_X1 U85661 ( .B1(n81378), .B2(n105355), .A(n97398), .ZN(
        \DLX_Datapath/RegisterFile/N23976 ) );
  AOI22_X1 U85662 ( .A1(n105353), .A2(n94672), .B1(n105350), .B2(n69545), .ZN(
        n97398) );
  OAI21_X1 U85663 ( .B1(n106209), .B2(n105355), .A(n97399), .ZN(
        \DLX_Datapath/RegisterFile/N23975 ) );
  AOI22_X1 U85664 ( .A1(n105353), .A2(n94674), .B1(n105351), .B2(n70206), .ZN(
        n97399) );
  OAI21_X1 U85665 ( .B1(n106204), .B2(n105355), .A(n97400), .ZN(
        \DLX_Datapath/RegisterFile/N23974 ) );
  AOI22_X1 U85666 ( .A1(n105353), .A2(n94676), .B1(n97396), .B2(n74052), .ZN(
        n97400) );
  OAI21_X1 U85667 ( .B1(n106099), .B2(n105355), .A(n97401), .ZN(
        \DLX_Datapath/RegisterFile/N23973 ) );
  AOI22_X1 U85668 ( .A1(n105353), .A2(n94678), .B1(n105351), .B2(n70639), .ZN(
        n97401) );
  OAI21_X1 U85669 ( .B1(n106255), .B2(n105355), .A(n97402), .ZN(
        \DLX_Datapath/RegisterFile/N23972 ) );
  AOI22_X1 U85670 ( .A1(n105353), .A2(n94680), .B1(n97396), .B2(n110794), .ZN(
        n97402) );
  OAI21_X1 U85671 ( .B1(n105992), .B2(n105355), .A(n97403), .ZN(
        \DLX_Datapath/RegisterFile/N23971 ) );
  AOI22_X1 U85672 ( .A1(n105353), .A2(n94682), .B1(n105351), .B2(n110893), 
        .ZN(n97403) );
  OAI21_X1 U85673 ( .B1(n80190), .B2(n105355), .A(n97404), .ZN(
        \DLX_Datapath/RegisterFile/N23970 ) );
  AOI22_X1 U85674 ( .A1(n105353), .A2(n94684), .B1(n105351), .B2(n110487), 
        .ZN(n97404) );
  OAI21_X1 U85675 ( .B1(n106191), .B2(n105354), .A(n97405), .ZN(
        \DLX_Datapath/RegisterFile/N23969 ) );
  AOI22_X1 U85676 ( .A1(n105352), .A2(n94686), .B1(n105350), .B2(n110270), 
        .ZN(n97405) );
  OAI21_X1 U85677 ( .B1(n106129), .B2(n105354), .A(n97406), .ZN(
        \DLX_Datapath/RegisterFile/N23968 ) );
  AOI22_X1 U85678 ( .A1(n105353), .A2(n94688), .B1(n105350), .B2(n110588), 
        .ZN(n97406) );
  OAI21_X1 U85679 ( .B1(n106186), .B2(n105354), .A(n97407), .ZN(
        \DLX_Datapath/RegisterFile/N23967 ) );
  AOI22_X1 U85680 ( .A1(n97395), .A2(n94690), .B1(n105350), .B2(n110379), .ZN(
        n97407) );
  OAI21_X1 U85681 ( .B1(n106164), .B2(n105354), .A(n97408), .ZN(
        \DLX_Datapath/RegisterFile/N23966 ) );
  AOI22_X1 U85682 ( .A1(n97395), .A2(n94692), .B1(n105350), .B2(n110055), .ZN(
        n97408) );
  OAI21_X1 U85683 ( .B1(n106105), .B2(n105354), .A(n97409), .ZN(
        \DLX_Datapath/RegisterFile/N23965 ) );
  AOI22_X1 U85684 ( .A1(n97395), .A2(n94694), .B1(n105350), .B2(n110162), .ZN(
        n97409) );
  OAI21_X1 U85685 ( .B1(n106219), .B2(n105354), .A(n97410), .ZN(
        \DLX_Datapath/RegisterFile/N23964 ) );
  AOI22_X1 U85686 ( .A1(n97395), .A2(n94696), .B1(n105350), .B2(n109946), .ZN(
        n97410) );
  OAI21_X1 U85687 ( .B1(n81398), .B2(n105354), .A(n97411), .ZN(
        \DLX_Datapath/RegisterFile/N23963 ) );
  AOI22_X1 U85688 ( .A1(n105353), .A2(n94698), .B1(n105350), .B2(n109829), 
        .ZN(n97411) );
  OAI21_X1 U85689 ( .B1(n106230), .B2(n105354), .A(n97412), .ZN(
        \DLX_Datapath/RegisterFile/N23962 ) );
  AOI22_X1 U85690 ( .A1(n105353), .A2(n94700), .B1(n105350), .B2(n108203), 
        .ZN(n97412) );
  OAI21_X1 U85691 ( .B1(n106172), .B2(n105354), .A(n97413), .ZN(
        \DLX_Datapath/RegisterFile/N23961 ) );
  AOI22_X1 U85692 ( .A1(n105353), .A2(n94702), .B1(n105350), .B2(n108326), 
        .ZN(n97413) );
  OAI21_X1 U85693 ( .B1(n106238), .B2(n105354), .A(n97414), .ZN(
        \DLX_Datapath/RegisterFile/N23960 ) );
  AOI22_X1 U85694 ( .A1(n97395), .A2(n94704), .B1(n105350), .B2(n108437), .ZN(
        n97414) );
  OAI21_X1 U85695 ( .B1(n106072), .B2(n105354), .A(n97415), .ZN(
        \DLX_Datapath/RegisterFile/N23959 ) );
  AOI22_X1 U85696 ( .A1(n97395), .A2(n94706), .B1(n105350), .B2(n107675), .ZN(
        n97415) );
  OAI21_X1 U85697 ( .B1(n106200), .B2(n105354), .A(n97416), .ZN(
        \DLX_Datapath/RegisterFile/N23958 ) );
  AOI22_X1 U85698 ( .A1(n105352), .A2(n94708), .B1(n105351), .B2(n109593), 
        .ZN(n97416) );
  OAI21_X1 U85699 ( .B1(n106245), .B2(n105355), .A(n97417), .ZN(
        \DLX_Datapath/RegisterFile/N23957 ) );
  AOI22_X1 U85700 ( .A1(n105352), .A2(n94710), .B1(n97396), .B2(n108554), .ZN(
        n97417) );
  OAI21_X1 U85701 ( .B1(n106159), .B2(n105355), .A(n97418), .ZN(
        \DLX_Datapath/RegisterFile/N23956 ) );
  AOI22_X1 U85702 ( .A1(n105352), .A2(n94712), .B1(n105351), .B2(n109698), 
        .ZN(n97418) );
  OAI21_X1 U85703 ( .B1(n81394), .B2(n105354), .A(n97419), .ZN(
        \DLX_Datapath/RegisterFile/N23955 ) );
  AOI22_X1 U85704 ( .A1(n105352), .A2(n94714), .B1(n105351), .B2(n109482), 
        .ZN(n97419) );
  OAI21_X1 U85705 ( .B1(n106009), .B2(n105355), .A(n97420), .ZN(
        \DLX_Datapath/RegisterFile/N23954 ) );
  AOI22_X1 U85706 ( .A1(n105352), .A2(n81259), .B1(n105351), .B2(n109019), 
        .ZN(n97420) );
  OAI21_X1 U85707 ( .B1(n106260), .B2(n105355), .A(n97421), .ZN(
        \DLX_Datapath/RegisterFile/N23953 ) );
  AOI22_X1 U85708 ( .A1(n105352), .A2(n94717), .B1(n97396), .B2(n109367), .ZN(
        n97421) );
  OAI21_X1 U85709 ( .B1(n106044), .B2(n105354), .A(n97422), .ZN(
        \DLX_Datapath/RegisterFile/N23952 ) );
  AOI22_X1 U85710 ( .A1(n105352), .A2(n94719), .B1(n105351), .B2(n109249), 
        .ZN(n97422) );
  OAI21_X1 U85711 ( .B1(n106049), .B2(n105355), .A(n97423), .ZN(
        \DLX_Datapath/RegisterFile/N23951 ) );
  AOI22_X1 U85712 ( .A1(n105352), .A2(n94721), .B1(n97396), .B2(n109141), .ZN(
        n97423) );
  OAI21_X1 U85713 ( .B1(n106095), .B2(n105354), .A(n97424), .ZN(
        \DLX_Datapath/RegisterFile/N23950 ) );
  AOI22_X1 U85714 ( .A1(n105352), .A2(n94723), .B1(n105351), .B2(n108676), 
        .ZN(n97424) );
  OAI21_X1 U85715 ( .B1(n106054), .B2(n105355), .A(n97425), .ZN(
        \DLX_Datapath/RegisterFile/N23949 ) );
  AOI22_X1 U85716 ( .A1(n105352), .A2(n94725), .B1(n97396), .B2(n108903), .ZN(
        n97425) );
  OAI21_X1 U85717 ( .B1(n105217), .B2(n105355), .A(n97426), .ZN(
        \DLX_Datapath/RegisterFile/N23948 ) );
  AOI22_X1 U85718 ( .A1(n105352), .A2(n94727), .B1(n97396), .B2(n108791), .ZN(
        n97426) );
  OAI21_X1 U85719 ( .B1(n106268), .B2(n105354), .A(n97427), .ZN(
        \DLX_Datapath/RegisterFile/N23947 ) );
  AOI22_X1 U85720 ( .A1(n105352), .A2(n94729), .B1(n105351), .B2(n107331), 
        .ZN(n97427) );
  NOR2_X1 U85721 ( .A1(n97356), .A2(n97428), .ZN(n97396) );
  AOI21_X1 U85722 ( .B1(n105205), .B2(n97318), .A(n94663), .ZN(n97356) );
  NOR2_X1 U85723 ( .A1(n97318), .A2(n97428), .ZN(n97395) );
  NOR2_X1 U85724 ( .A1(n97393), .A2(n105089), .ZN(n97428) );
  OR2_X1 U85725 ( .A1(n97061), .A2(n86230), .ZN(n97318) );
  NAND2_X1 U85726 ( .A1(n94734), .A2(n105127), .ZN(n97393) );
  OAI21_X1 U85727 ( .B1(n106067), .B2(n105970), .A(n97429), .ZN(
        \DLX_Datapath/RegisterFile/N23945 ) );
  AOI22_X1 U85728 ( .A1(n106066), .A2(n107988), .B1(n94511), .B2(n106063), 
        .ZN(n97429) );
  OAI21_X1 U85729 ( .B1(n106137), .B2(n106067), .A(n97430), .ZN(
        \DLX_Datapath/RegisterFile/N23944 ) );
  AOI22_X1 U85730 ( .A1(n106066), .A2(n107256), .B1(n81539), .B2(n81462), .ZN(
        n97430) );
  OAI21_X1 U85731 ( .B1(n106209), .B2(n106067), .A(n97431), .ZN(
        \DLX_Datapath/RegisterFile/N23943 ) );
  AOI22_X1 U85732 ( .A1(n106066), .A2(n107795), .B1(n106063), .B2(n81301), 
        .ZN(n97431) );
  OAI21_X1 U85733 ( .B1(n106100), .B2(n106067), .A(n97432), .ZN(
        \DLX_Datapath/RegisterFile/N23941 ) );
  AOI22_X1 U85734 ( .A1(n106066), .A2(n108095), .B1(n94516), .B2(n81462), .ZN(
        n97432) );
  OAI21_X1 U85735 ( .B1(n106068), .B2(n81629), .A(n97433), .ZN(
        \DLX_Datapath/RegisterFile/N23939 ) );
  AOI22_X1 U85736 ( .A1(n106066), .A2(n110894), .B1(n94519), .B2(n106064), 
        .ZN(n97433) );
  OAI21_X1 U85737 ( .B1(n80190), .B2(n106067), .A(n97434), .ZN(
        \DLX_Datapath/RegisterFile/N23938 ) );
  AOI22_X1 U85738 ( .A1(n106066), .A2(n110488), .B1(n106063), .B2(n80192), 
        .ZN(n97434) );
  OAI21_X1 U85739 ( .B1(n106129), .B2(n106067), .A(n97435), .ZN(
        \DLX_Datapath/RegisterFile/N23936 ) );
  AOI22_X1 U85740 ( .A1(n106066), .A2(n110589), .B1(n94523), .B2(n81462), .ZN(
        n97435) );
  OAI21_X1 U85741 ( .B1(n106105), .B2(n106067), .A(n97436), .ZN(
        \DLX_Datapath/RegisterFile/N23933 ) );
  AOI22_X1 U85742 ( .A1(n106066), .A2(n110163), .B1(n94527), .B2(n81462), .ZN(
        n97436) );
  OAI21_X1 U85743 ( .B1(n106219), .B2(n106067), .A(n97437), .ZN(
        \DLX_Datapath/RegisterFile/N23932 ) );
  AOI22_X1 U85744 ( .A1(n106065), .A2(n109947), .B1(n106063), .B2(n81297), 
        .ZN(n97437) );
  OAI21_X1 U85745 ( .B1(n106110), .B2(n106068), .A(n97438), .ZN(
        \DLX_Datapath/RegisterFile/N23931 ) );
  AOI22_X1 U85746 ( .A1(n106065), .A2(n109830), .B1(n94530), .B2(n81462), .ZN(
        n97438) );
  OAI21_X1 U85747 ( .B1(n106172), .B2(n106068), .A(n97439), .ZN(
        \DLX_Datapath/RegisterFile/N23929 ) );
  AOI22_X1 U85748 ( .A1(n106065), .A2(n108327), .B1(n106063), .B2(n106168), 
        .ZN(n97439) );
  OAI21_X1 U85749 ( .B1(n106198), .B2(n106068), .A(n97440), .ZN(
        \DLX_Datapath/RegisterFile/N23926 ) );
  AOI22_X1 U85750 ( .A1(n106065), .A2(n109594), .B1(n94536), .B2(n81462), .ZN(
        n97440) );
  OAI21_X1 U85751 ( .B1(n106159), .B2(n106067), .A(n97441), .ZN(
        \DLX_Datapath/RegisterFile/N23924 ) );
  AOI22_X1 U85752 ( .A1(n106065), .A2(n109699), .B1(n106063), .B2(n81351), 
        .ZN(n97441) );
  OAI21_X1 U85753 ( .B1(n106115), .B2(n106067), .A(n97442), .ZN(
        \DLX_Datapath/RegisterFile/N23923 ) );
  AOI22_X1 U85754 ( .A1(n106065), .A2(n109483), .B1(n106021), .B2(n81462), 
        .ZN(n97442) );
  OAI21_X1 U85755 ( .B1(n106009), .B2(n106068), .A(n97443), .ZN(
        \DLX_Datapath/RegisterFile/N23922 ) );
  AOI22_X1 U85756 ( .A1(n106065), .A2(n109020), .B1(n94541), .B2(n106063), 
        .ZN(n97443) );
  OAI21_X1 U85757 ( .B1(n106067), .B2(n81509), .A(n97444), .ZN(
        \DLX_Datapath/RegisterFile/N23920 ) );
  AOI22_X1 U85758 ( .A1(n106065), .A2(n109250), .B1(n105625), .B2(n106063), 
        .ZN(n97444) );
  OAI21_X1 U85759 ( .B1(n106068), .B2(n106049), .A(n97445), .ZN(
        \DLX_Datapath/RegisterFile/N23919 ) );
  AOI22_X1 U85760 ( .A1(n106065), .A2(n109142), .B1(n94546), .B2(n106063), 
        .ZN(n97445) );
  OAI21_X1 U85761 ( .B1(n106095), .B2(n106067), .A(n97446), .ZN(
        \DLX_Datapath/RegisterFile/N23918 ) );
  AOI22_X1 U85762 ( .A1(n106065), .A2(n108677), .B1(n94548), .B2(n81462), .ZN(
        n97446) );
  OAI21_X1 U85763 ( .B1(n106067), .B2(n81498), .A(n97447), .ZN(
        \DLX_Datapath/RegisterFile/N23917 ) );
  AOI22_X1 U85764 ( .A1(n106065), .A2(n108904), .B1(n81783), .B2(n106063), 
        .ZN(n97447) );
  OAI21_X1 U85765 ( .B1(n106268), .B2(n106068), .A(n97448), .ZN(
        \DLX_Datapath/RegisterFile/N23915 ) );
  AOI22_X1 U85766 ( .A1(n106065), .A2(n107332), .B1(n106064), .B2(n81265), 
        .ZN(n97448) );
  NOR2_X1 U85767 ( .A1(n97449), .A2(n104691), .ZN(n81462) );
  AOI21_X1 U85768 ( .B1(n97058), .B2(n94771), .A(n97450), .ZN(n81461) );
  NOR2_X1 U85769 ( .A1(n81459), .A2(n105092), .ZN(n97450) );
  NAND2_X1 U85770 ( .A1(n97061), .A2(n105199), .ZN(n97058) );
  NAND2_X1 U85771 ( .A1(n105128), .A2(n94772), .ZN(n81459) );
  OAI21_X1 U85772 ( .B1(n106148), .B2(n105349), .A(n97452), .ZN(
        \DLX_Datapath/RegisterFile/N23914 ) );
  AOI22_X1 U85773 ( .A1(n104870), .A2(n94559), .B1(n105347), .B2(n107894), 
        .ZN(n97452) );
  OAI21_X1 U85774 ( .B1(n105970), .B2(n105349), .A(n97455), .ZN(
        \DLX_Datapath/RegisterFile/N23913 ) );
  AOI22_X1 U85775 ( .A1(n104869), .A2(n94562), .B1(n105346), .B2(n70494), .ZN(
        n97455) );
  OAI21_X1 U85776 ( .B1(n106137), .B2(n105349), .A(n97456), .ZN(
        \DLX_Datapath/RegisterFile/N23912 ) );
  AOI22_X1 U85777 ( .A1(n104869), .A2(n94564), .B1(n105347), .B2(n107257), 
        .ZN(n97456) );
  OAI21_X1 U85778 ( .B1(n106209), .B2(n105349), .A(n97457), .ZN(
        \DLX_Datapath/RegisterFile/N23911 ) );
  AOI22_X1 U85779 ( .A1(n97453), .A2(n94566), .B1(n105346), .B2(n70208), .ZN(
        n97457) );
  OAI21_X1 U85780 ( .B1(n106206), .B2(n105349), .A(n97458), .ZN(
        \DLX_Datapath/RegisterFile/N23910 ) );
  AOI22_X1 U85781 ( .A1(n104870), .A2(n94568), .B1(n105347), .B2(n110696), 
        .ZN(n97458) );
  OAI21_X1 U85782 ( .B1(n106100), .B2(n105349), .A(n97459), .ZN(
        \DLX_Datapath/RegisterFile/N23909 ) );
  AOI22_X1 U85783 ( .A1(n97453), .A2(n94570), .B1(n105346), .B2(n108096), .ZN(
        n97459) );
  OAI21_X1 U85784 ( .B1(n106255), .B2(n105349), .A(n97460), .ZN(
        \DLX_Datapath/RegisterFile/N23908 ) );
  AOI22_X1 U85785 ( .A1(n104869), .A2(n94572), .B1(n105347), .B2(n110796), 
        .ZN(n97460) );
  OAI21_X1 U85786 ( .B1(n105991), .B2(n105349), .A(n97461), .ZN(
        \DLX_Datapath/RegisterFile/N23907 ) );
  AOI22_X1 U85787 ( .A1(n104869), .A2(n94574), .B1(n105346), .B2(n110895), 
        .ZN(n97461) );
  OAI21_X1 U85788 ( .B1(n106331), .B2(n105349), .A(n97462), .ZN(
        \DLX_Datapath/RegisterFile/N23906 ) );
  AOI22_X1 U85789 ( .A1(n104870), .A2(n94576), .B1(n105346), .B2(n110489), 
        .ZN(n97462) );
  OAI21_X1 U85790 ( .B1(n106191), .B2(n105348), .A(n97463), .ZN(
        \DLX_Datapath/RegisterFile/N23905 ) );
  AOI22_X1 U85791 ( .A1(n104870), .A2(n94578), .B1(n97454), .B2(n110272), .ZN(
        n97463) );
  OAI21_X1 U85792 ( .B1(n106130), .B2(n105348), .A(n97464), .ZN(
        \DLX_Datapath/RegisterFile/N23904 ) );
  AOI22_X1 U85793 ( .A1(n104869), .A2(n94580), .B1(n97454), .B2(n110590), .ZN(
        n97464) );
  OAI21_X1 U85794 ( .B1(n106186), .B2(n105348), .A(n97465), .ZN(
        \DLX_Datapath/RegisterFile/N23903 ) );
  AOI22_X1 U85795 ( .A1(n104869), .A2(n94582), .B1(n97454), .B2(n110381), .ZN(
        n97465) );
  OAI21_X1 U85796 ( .B1(n106164), .B2(n105348), .A(n97466), .ZN(
        \DLX_Datapath/RegisterFile/N23902 ) );
  AOI22_X1 U85797 ( .A1(n104869), .A2(n94584), .B1(n97454), .B2(n110057), .ZN(
        n97466) );
  OAI21_X1 U85798 ( .B1(n106105), .B2(n105348), .A(n97467), .ZN(
        \DLX_Datapath/RegisterFile/N23901 ) );
  AOI22_X1 U85799 ( .A1(n104870), .A2(n94586), .B1(n105346), .B2(n110164), 
        .ZN(n97467) );
  OAI21_X1 U85800 ( .B1(n106219), .B2(n105348), .A(n97468), .ZN(
        \DLX_Datapath/RegisterFile/N23900 ) );
  AOI22_X1 U85801 ( .A1(n104869), .A2(n94588), .B1(n97454), .B2(n109948), .ZN(
        n97468) );
  OAI21_X1 U85802 ( .B1(n106110), .B2(n105348), .A(n97469), .ZN(
        \DLX_Datapath/RegisterFile/N23899 ) );
  AOI22_X1 U85803 ( .A1(n97453), .A2(n94590), .B1(n97454), .B2(n109831), .ZN(
        n97469) );
  OAI21_X1 U85804 ( .B1(n106232), .B2(n105348), .A(n97470), .ZN(
        \DLX_Datapath/RegisterFile/N23898 ) );
  AOI22_X1 U85805 ( .A1(n97453), .A2(n94592), .B1(n97454), .B2(n108205), .ZN(
        n97470) );
  OAI21_X1 U85806 ( .B1(n106172), .B2(n105348), .A(n97471), .ZN(
        \DLX_Datapath/RegisterFile/N23897 ) );
  AOI22_X1 U85807 ( .A1(n104870), .A2(n94594), .B1(n105347), .B2(n108328), 
        .ZN(n97471) );
  OAI21_X1 U85808 ( .B1(n106235), .B2(n105348), .A(n97472), .ZN(
        \DLX_Datapath/RegisterFile/N23896 ) );
  AOI22_X1 U85809 ( .A1(n104870), .A2(n94596), .B1(n105346), .B2(n108439), 
        .ZN(n97472) );
  OAI21_X1 U85810 ( .B1(n106071), .B2(n105348), .A(n97473), .ZN(
        \DLX_Datapath/RegisterFile/N23895 ) );
  AOI22_X1 U85811 ( .A1(n104869), .A2(n94598), .B1(n97454), .B2(n107677), .ZN(
        n97473) );
  OAI21_X1 U85812 ( .B1(n106197), .B2(n105348), .A(n97474), .ZN(
        \DLX_Datapath/RegisterFile/N23894 ) );
  AOI22_X1 U85813 ( .A1(n104869), .A2(n94600), .B1(n105346), .B2(n109595), 
        .ZN(n97474) );
  OAI21_X1 U85814 ( .B1(n106245), .B2(n105349), .A(n97475), .ZN(
        \DLX_Datapath/RegisterFile/N23893 ) );
  AOI22_X1 U85815 ( .A1(n97453), .A2(n94602), .B1(n105347), .B2(n108556), .ZN(
        n97475) );
  OAI21_X1 U85816 ( .B1(n106159), .B2(n105349), .A(n97476), .ZN(
        \DLX_Datapath/RegisterFile/N23892 ) );
  AOI22_X1 U85817 ( .A1(n104869), .A2(n94604), .B1(n105346), .B2(n109700), 
        .ZN(n97476) );
  OAI21_X1 U85818 ( .B1(n106115), .B2(n105348), .A(n97477), .ZN(
        \DLX_Datapath/RegisterFile/N23891 ) );
  AOI22_X1 U85819 ( .A1(n97453), .A2(n94606), .B1(n105347), .B2(n109484), .ZN(
        n97477) );
  OAI21_X1 U85820 ( .B1(n106010), .B2(n105349), .A(n97478), .ZN(
        \DLX_Datapath/RegisterFile/N23890 ) );
  AOI22_X1 U85821 ( .A1(n104870), .A2(n94608), .B1(n105346), .B2(n109021), 
        .ZN(n97478) );
  OAI21_X1 U85822 ( .B1(n106260), .B2(n105349), .A(n97479), .ZN(
        \DLX_Datapath/RegisterFile/N23889 ) );
  AOI22_X1 U85823 ( .A1(n104870), .A2(n94610), .B1(n105346), .B2(n109369), 
        .ZN(n97479) );
  OAI21_X1 U85824 ( .B1(n106044), .B2(n105348), .A(n97480), .ZN(
        \DLX_Datapath/RegisterFile/N23888 ) );
  AOI22_X1 U85825 ( .A1(n104869), .A2(n94612), .B1(n105347), .B2(n109251), 
        .ZN(n97480) );
  OAI21_X1 U85826 ( .B1(n106050), .B2(n105349), .A(n97481), .ZN(
        \DLX_Datapath/RegisterFile/N23887 ) );
  AOI22_X1 U85827 ( .A1(n104870), .A2(n94614), .B1(n105346), .B2(n109143), 
        .ZN(n97481) );
  OAI21_X1 U85828 ( .B1(n106095), .B2(n105348), .A(n97482), .ZN(
        \DLX_Datapath/RegisterFile/N23886 ) );
  AOI22_X1 U85829 ( .A1(n97453), .A2(n94616), .B1(n105347), .B2(n108678), .ZN(
        n97482) );
  OAI21_X1 U85830 ( .B1(n106055), .B2(n105349), .A(n97483), .ZN(
        \DLX_Datapath/RegisterFile/N23885 ) );
  AOI22_X1 U85831 ( .A1(n104870), .A2(n94618), .B1(n105346), .B2(n108905), 
        .ZN(n97483) );
  OAI21_X1 U85832 ( .B1(n105217), .B2(n105349), .A(n97484), .ZN(
        \DLX_Datapath/RegisterFile/N23884 ) );
  AOI22_X1 U85833 ( .A1(n97453), .A2(n94620), .B1(n105347), .B2(n108793), .ZN(
        n97484) );
  OAI21_X1 U85834 ( .B1(n106268), .B2(n105348), .A(n97485), .ZN(
        \DLX_Datapath/RegisterFile/N23883 ) );
  AOI22_X1 U85835 ( .A1(n104869), .A2(n94622), .B1(n105347), .B2(n107333), 
        .ZN(n97485) );
  NOR2_X1 U85836 ( .A1(n97486), .A2(n97487), .ZN(n97454) );
  NOR2_X1 U85837 ( .A1(n97449), .A2(n97487), .ZN(n97453) );
  NOR2_X1 U85838 ( .A1(n97451), .A2(n105089), .ZN(n97487) );
  NAND2_X1 U85839 ( .A1(n105128), .A2(n94810), .ZN(n97451) );
  OAI21_X1 U85840 ( .B1(n106041), .B2(n81651), .A(n97488), .ZN(
        \DLX_Datapath/RegisterFile/N23881 ) );
  AOI22_X1 U85841 ( .A1(n81653), .A2(n104852), .B1(n106040), .B2(n107989), 
        .ZN(n97488) );
  OAI21_X1 U85842 ( .B1(n106137), .B2(n106042), .A(n97489), .ZN(
        \DLX_Datapath/RegisterFile/N23880 ) );
  AOI22_X1 U85843 ( .A1(n104853), .A2(n81380), .B1(n106040), .B2(n107258), 
        .ZN(n97489) );
  OAI21_X1 U85844 ( .B1(n106209), .B2(n106041), .A(n97490), .ZN(
        \DLX_Datapath/RegisterFile/N23879 ) );
  AOI22_X1 U85845 ( .A1(n104853), .A2(n81377), .B1(n70209), .B2(n106039), .ZN(
        n97490) );
  OAI21_X1 U85846 ( .B1(n106203), .B2(n106041), .A(n97491), .ZN(
        \DLX_Datapath/RegisterFile/N23878 ) );
  AOI22_X1 U85847 ( .A1(n104852), .A2(n81428), .B1(n74055), .B2(n106039), .ZN(
        n97491) );
  OAI21_X1 U85848 ( .B1(n106100), .B2(n106041), .A(n97492), .ZN(
        \DLX_Datapath/RegisterFile/N23877 ) );
  AOI22_X1 U85849 ( .A1(n104853), .A2(n81410), .B1(n106040), .B2(n108097), 
        .ZN(n97492) );
  OAI21_X1 U85850 ( .B1(n106255), .B2(n106041), .A(n97493), .ZN(
        \DLX_Datapath/RegisterFile/N23876 ) );
  AOI22_X1 U85851 ( .A1(n81700), .A2(n104853), .B1(n74196), .B2(n106039), .ZN(
        n97493) );
  OAI21_X1 U85852 ( .B1(n106042), .B2(n105992), .A(n97494), .ZN(
        \DLX_Datapath/RegisterFile/N23875 ) );
  AOI22_X1 U85853 ( .A1(n81632), .A2(n104853), .B1(n74336), .B2(n106039), .ZN(
        n97494) );
  OAI21_X1 U85854 ( .B1(n106331), .B2(n106041), .A(n97495), .ZN(
        \DLX_Datapath/RegisterFile/N23874 ) );
  AOI22_X1 U85855 ( .A1(n81515), .A2(n81414), .B1(n73772), .B2(n106039), .ZN(
        n97495) );
  OAI21_X1 U85856 ( .B1(n106191), .B2(n106041), .A(n97496), .ZN(
        \DLX_Datapath/RegisterFile/N23873 ) );
  AOI22_X1 U85857 ( .A1(n104853), .A2(n81317), .B1(n73476), .B2(n106039), .ZN(
        n97496) );
  OAI21_X1 U85858 ( .B1(n106128), .B2(n106041), .A(n97497), .ZN(
        \DLX_Datapath/RegisterFile/N23872 ) );
  AOI22_X1 U85859 ( .A1(n81515), .A2(n81386), .B1(n73913), .B2(n106039), .ZN(
        n97497) );
  OAI21_X1 U85860 ( .B1(n106186), .B2(n106041), .A(n97498), .ZN(
        \DLX_Datapath/RegisterFile/N23871 ) );
  AOI22_X1 U85861 ( .A1(n104852), .A2(n81320), .B1(n73625), .B2(n106039), .ZN(
        n97498) );
  OAI21_X1 U85862 ( .B1(n106164), .B2(n106041), .A(n97499), .ZN(
        \DLX_Datapath/RegisterFile/N23870 ) );
  AOI22_X1 U85863 ( .A1(n81604), .A2(n104852), .B1(n106040), .B2(n110058), 
        .ZN(n97499) );
  OAI21_X1 U85864 ( .B1(n106105), .B2(n106041), .A(n97500), .ZN(
        \DLX_Datapath/RegisterFile/N23869 ) );
  AOI22_X1 U85865 ( .A1(n81515), .A2(n81405), .B1(n106040), .B2(n110165), .ZN(
        n97500) );
  OAI21_X1 U85866 ( .B1(n106219), .B2(n106042), .A(n97501), .ZN(
        \DLX_Datapath/RegisterFile/N23868 ) );
  AOI22_X1 U85867 ( .A1(n104852), .A2(n81402), .B1(n106040), .B2(n109949), 
        .ZN(n97501) );
  OAI21_X1 U85868 ( .B1(n106110), .B2(n106042), .A(n97502), .ZN(
        \DLX_Datapath/RegisterFile/N23867 ) );
  AOI22_X1 U85869 ( .A1(n81515), .A2(n81400), .B1(n81516), .B2(n109832), .ZN(
        n97502) );
  OAI21_X1 U85870 ( .B1(n106172), .B2(n106042), .A(n97503), .ZN(
        \DLX_Datapath/RegisterFile/N23865 ) );
  AOI22_X1 U85871 ( .A1(n104852), .A2(n81373), .B1(n106040), .B2(n108329), 
        .ZN(n97503) );
  OAI21_X1 U85872 ( .B1(n106199), .B2(n106042), .A(n97504), .ZN(
        \DLX_Datapath/RegisterFile/N23862 ) );
  AOI22_X1 U85873 ( .A1(n104853), .A2(n81313), .B1(n81516), .B2(n109596), .ZN(
        n97504) );
  OAI21_X1 U85874 ( .B1(n106159), .B2(n106042), .A(n97505), .ZN(
        \DLX_Datapath/RegisterFile/N23860 ) );
  AOI22_X1 U85875 ( .A1(n104852), .A2(n81425), .B1(n106039), .B2(n109701), 
        .ZN(n97505) );
  OAI21_X1 U85876 ( .B1(n106115), .B2(n106042), .A(n97506), .ZN(
        \DLX_Datapath/RegisterFile/N23859 ) );
  AOI22_X1 U85877 ( .A1(n81515), .A2(n81396), .B1(n81516), .B2(n109485), .ZN(
        n97506) );
  OAI21_X1 U85878 ( .B1(n106010), .B2(n106042), .A(n97507), .ZN(
        \DLX_Datapath/RegisterFile/N23858 ) );
  AOI22_X1 U85879 ( .A1(n81590), .A2(n104852), .B1(n81516), .B2(n109022), .ZN(
        n97507) );
  OAI21_X1 U85880 ( .B1(n106044), .B2(n106042), .A(n97508), .ZN(
        \DLX_Datapath/RegisterFile/N23856 ) );
  AOI22_X1 U85881 ( .A1(n81515), .A2(n81511), .B1(n106040), .B2(n109252), .ZN(
        n97508) );
  OAI21_X1 U85882 ( .B1(n106095), .B2(n106042), .A(n97509), .ZN(
        \DLX_Datapath/RegisterFile/N23854 ) );
  AOI22_X1 U85883 ( .A1(n104853), .A2(n81417), .B1(n81516), .B2(n108679), .ZN(
        n97509) );
  OAI21_X1 U85884 ( .B1(n106268), .B2(n106042), .A(n97510), .ZN(
        \DLX_Datapath/RegisterFile/N23851 ) );
  AOI22_X1 U85885 ( .A1(n104852), .A2(n81327), .B1(n106039), .B2(n107334), 
        .ZN(n97510) );
  NOR2_X1 U85886 ( .A1(n97486), .A2(n97511), .ZN(n81516) );
  NOR2_X1 U85887 ( .A1(n97449), .A2(n104695), .ZN(n81515) );
  NOR2_X1 U85888 ( .A1(n81513), .A2(n105092), .ZN(n97511) );
  NAND2_X1 U85889 ( .A1(n105127), .A2(n94853), .ZN(n81513) );
  OAI21_X1 U85890 ( .B1(n106148), .B2(n105345), .A(n97513), .ZN(
        \DLX_Datapath/RegisterFile/N23850 ) );
  AOI22_X1 U85891 ( .A1(n105343), .A2(n94667), .B1(n97515), .B2(n70354), .ZN(
        n97513) );
  OAI21_X1 U85892 ( .B1(n105971), .B2(n105345), .A(n97516), .ZN(
        \DLX_Datapath/RegisterFile/N23849 ) );
  AOI22_X1 U85893 ( .A1(n97514), .A2(n94670), .B1(n105341), .B2(n70496), .ZN(
        n97516) );
  OAI21_X1 U85894 ( .B1(n106137), .B2(n105344), .A(n97517), .ZN(
        \DLX_Datapath/RegisterFile/N23848 ) );
  AOI22_X1 U85895 ( .A1(n105343), .A2(n94672), .B1(n97515), .B2(n69549), .ZN(
        n97517) );
  OAI21_X1 U85896 ( .B1(n106209), .B2(n105344), .A(n97518), .ZN(
        \DLX_Datapath/RegisterFile/N23847 ) );
  AOI22_X1 U85897 ( .A1(n97514), .A2(n94674), .B1(n105341), .B2(n70210), .ZN(
        n97518) );
  OAI21_X1 U85898 ( .B1(n106206), .B2(n105344), .A(n97519), .ZN(
        \DLX_Datapath/RegisterFile/N23846 ) );
  AOI22_X1 U85899 ( .A1(n105343), .A2(n94676), .B1(n97515), .B2(n74056), .ZN(
        n97519) );
  OAI21_X1 U85900 ( .B1(n106100), .B2(n105345), .A(n97520), .ZN(
        \DLX_Datapath/RegisterFile/N23845 ) );
  AOI22_X1 U85901 ( .A1(n105342), .A2(n94678), .B1(n105341), .B2(n70643), .ZN(
        n97520) );
  OAI21_X1 U85902 ( .B1(n106255), .B2(n105344), .A(n97521), .ZN(
        \DLX_Datapath/RegisterFile/N23844 ) );
  AOI22_X1 U85903 ( .A1(n105343), .A2(n94680), .B1(n97515), .B2(n74197), .ZN(
        n97521) );
  OAI21_X1 U85904 ( .B1(n105992), .B2(n105344), .A(n97522), .ZN(
        \DLX_Datapath/RegisterFile/N23843 ) );
  AOI22_X1 U85905 ( .A1(n97514), .A2(n94682), .B1(n105341), .B2(n74337), .ZN(
        n97522) );
  OAI21_X1 U85906 ( .B1(n106330), .B2(n105345), .A(n97523), .ZN(
        \DLX_Datapath/RegisterFile/N23842 ) );
  AOI22_X1 U85907 ( .A1(n97514), .A2(n94684), .B1(n105341), .B2(n73773), .ZN(
        n97523) );
  OAI21_X1 U85908 ( .B1(n106191), .B2(n105345), .A(n97524), .ZN(
        \DLX_Datapath/RegisterFile/N23841 ) );
  AOI22_X1 U85909 ( .A1(n105342), .A2(n94686), .B1(n105340), .B2(n73477), .ZN(
        n97524) );
  OAI21_X1 U85910 ( .B1(n106130), .B2(n105345), .A(n97525), .ZN(
        \DLX_Datapath/RegisterFile/N23840 ) );
  AOI22_X1 U85911 ( .A1(n105342), .A2(n94688), .B1(n105340), .B2(n73914), .ZN(
        n97525) );
  OAI21_X1 U85912 ( .B1(n106186), .B2(n105345), .A(n97526), .ZN(
        \DLX_Datapath/RegisterFile/N23839 ) );
  AOI22_X1 U85913 ( .A1(n105342), .A2(n94690), .B1(n105340), .B2(n73626), .ZN(
        n97526) );
  OAI21_X1 U85914 ( .B1(n106164), .B2(n105345), .A(n97527), .ZN(
        \DLX_Datapath/RegisterFile/N23838 ) );
  AOI22_X1 U85915 ( .A1(n105342), .A2(n94692), .B1(n105340), .B2(n73188), .ZN(
        n97527) );
  OAI21_X1 U85916 ( .B1(n106105), .B2(n105345), .A(n97528), .ZN(
        \DLX_Datapath/RegisterFile/N23837 ) );
  AOI22_X1 U85917 ( .A1(n105342), .A2(n94694), .B1(n105340), .B2(n73330), .ZN(
        n97528) );
  OAI21_X1 U85918 ( .B1(n106219), .B2(n105345), .A(n97529), .ZN(
        \DLX_Datapath/RegisterFile/N23836 ) );
  AOI22_X1 U85919 ( .A1(n105342), .A2(n94696), .B1(n105340), .B2(n73046), .ZN(
        n97529) );
  OAI21_X1 U85920 ( .B1(n106110), .B2(n105345), .A(n97530), .ZN(
        \DLX_Datapath/RegisterFile/N23835 ) );
  AOI22_X1 U85921 ( .A1(n105342), .A2(n94698), .B1(n105340), .B2(n72896), .ZN(
        n97530) );
  OAI21_X1 U85922 ( .B1(n106233), .B2(n105345), .A(n97531), .ZN(
        \DLX_Datapath/RegisterFile/N23834 ) );
  AOI22_X1 U85923 ( .A1(n105342), .A2(n94700), .B1(n105340), .B2(n70792), .ZN(
        n97531) );
  OAI21_X1 U85924 ( .B1(n106172), .B2(n105345), .A(n97532), .ZN(
        \DLX_Datapath/RegisterFile/N23833 ) );
  AOI22_X1 U85925 ( .A1(n105342), .A2(n94702), .B1(n105340), .B2(n70951), .ZN(
        n97532) );
  OAI21_X1 U85926 ( .B1(n81281), .B2(n105345), .A(n97533), .ZN(
        \DLX_Datapath/RegisterFile/N23832 ) );
  AOI22_X1 U85927 ( .A1(n105342), .A2(n94704), .B1(n105340), .B2(n71096), .ZN(
        n97533) );
  OAI21_X1 U85928 ( .B1(n106071), .B2(n105345), .A(n97534), .ZN(
        \DLX_Datapath/RegisterFile/N23831 ) );
  AOI22_X1 U85929 ( .A1(n105342), .A2(n94706), .B1(n105340), .B2(n70057), .ZN(
        n97534) );
  OAI21_X1 U85930 ( .B1(n106198), .B2(n105345), .A(n97535), .ZN(
        \DLX_Datapath/RegisterFile/N23830 ) );
  AOI22_X1 U85931 ( .A1(n105342), .A2(n94708), .B1(n105341), .B2(n72586), .ZN(
        n97535) );
  OAI21_X1 U85932 ( .B1(n106245), .B2(n105344), .A(n97536), .ZN(
        \DLX_Datapath/RegisterFile/N23829 ) );
  AOI22_X1 U85933 ( .A1(n105343), .A2(n94710), .B1(n97515), .B2(n71245), .ZN(
        n97536) );
  OAI21_X1 U85934 ( .B1(n106159), .B2(n105344), .A(n97537), .ZN(
        \DLX_Datapath/RegisterFile/N23828 ) );
  AOI22_X1 U85935 ( .A1(n105342), .A2(n94712), .B1(n105341), .B2(n72728), .ZN(
        n97537) );
  OAI21_X1 U85936 ( .B1(n106115), .B2(n105344), .A(n97538), .ZN(
        \DLX_Datapath/RegisterFile/N23827 ) );
  AOI22_X1 U85937 ( .A1(n105343), .A2(n94714), .B1(n97515), .B2(n72438), .ZN(
        n97538) );
  OAI21_X1 U85938 ( .B1(n106010), .B2(n105344), .A(n97539), .ZN(
        \DLX_Datapath/RegisterFile/N23826 ) );
  AOI22_X1 U85939 ( .A1(n97514), .A2(n81259), .B1(n105341), .B2(n71838), .ZN(
        n97539) );
  OAI21_X1 U85940 ( .B1(n106260), .B2(n105344), .A(n97540), .ZN(
        \DLX_Datapath/RegisterFile/N23825 ) );
  AOI22_X1 U85941 ( .A1(n105343), .A2(n94717), .B1(n105340), .B2(n72287), .ZN(
        n97540) );
  OAI21_X1 U85942 ( .B1(n106045), .B2(n105344), .A(n97541), .ZN(
        \DLX_Datapath/RegisterFile/N23824 ) );
  AOI22_X1 U85943 ( .A1(n97514), .A2(n94719), .B1(n105341), .B2(n72136), .ZN(
        n97541) );
  OAI21_X1 U85944 ( .B1(n106050), .B2(n105344), .A(n97542), .ZN(
        \DLX_Datapath/RegisterFile/N23823 ) );
  AOI22_X1 U85945 ( .A1(n105343), .A2(n94721), .B1(n97515), .B2(n71992), .ZN(
        n97542) );
  OAI21_X1 U85946 ( .B1(n106095), .B2(n105344), .A(n97543), .ZN(
        \DLX_Datapath/RegisterFile/N23822 ) );
  AOI22_X1 U85947 ( .A1(n105343), .A2(n94723), .B1(n105341), .B2(n71394), .ZN(
        n97543) );
  OAI21_X1 U85948 ( .B1(n106055), .B2(n105344), .A(n97544), .ZN(
        \DLX_Datapath/RegisterFile/N23821 ) );
  AOI22_X1 U85949 ( .A1(n105343), .A2(n94725), .B1(n97515), .B2(n71689), .ZN(
        n97544) );
  OAI21_X1 U85950 ( .B1(n105217), .B2(n105344), .A(n97545), .ZN(
        \DLX_Datapath/RegisterFile/N23820 ) );
  AOI22_X1 U85951 ( .A1(n105343), .A2(n94727), .B1(n105341), .B2(n71545), .ZN(
        n97545) );
  OAI21_X1 U85952 ( .B1(n106268), .B2(n105344), .A(n97546), .ZN(
        \DLX_Datapath/RegisterFile/N23819 ) );
  AOI22_X1 U85953 ( .A1(n97514), .A2(n94729), .B1(n105341), .B2(n69654), .ZN(
        n97546) );
  NOR2_X1 U85954 ( .A1(n97486), .A2(n97547), .ZN(n97515) );
  AOI21_X1 U85955 ( .B1(n105205), .B2(n97449), .A(n94663), .ZN(n97486) );
  NOR2_X1 U85956 ( .A1(n97449), .A2(n97547), .ZN(n97514) );
  NOR2_X1 U85957 ( .A1(n97512), .A2(n105091), .ZN(n97547) );
  OR2_X1 U85958 ( .A1(n97061), .A2(n94848), .ZN(n97449) );
  OR2_X1 U85959 ( .A1(n95411), .A2(n96488), .ZN(n97061) );
  NAND2_X1 U85960 ( .A1(n106763), .A2(n94852), .ZN(n95411) );
  NAND2_X1 U85961 ( .A1(n94892), .A2(n105128), .ZN(n97512) );
  NOR2_X1 U85962 ( .A1(n97033), .A2(n95412), .ZN(n97062) );
  OR2_X1 U85963 ( .A1(n96530), .A2(n94895), .ZN(n97033) );
  OAI21_X1 U85964 ( .B1(n106180), .B2(n106147), .A(n97548), .ZN(
        \DLX_Datapath/RegisterFile/N23818 ) );
  AOI22_X1 U85965 ( .A1(n81360), .A2(n81338), .B1(n70355), .B2(n81339), .ZN(
        n97548) );
  OAI21_X1 U85966 ( .B1(n106180), .B2(n105969), .A(n97549), .ZN(
        \DLX_Datapath/RegisterFile/N23817 ) );
  AOI22_X1 U85967 ( .A1(n94511), .A2(n81338), .B1(n70497), .B2(n106176), .ZN(
        n97549) );
  OAI21_X1 U85968 ( .B1(n106179), .B2(n81378), .A(n97550), .ZN(
        \DLX_Datapath/RegisterFile/N23816 ) );
  AOI22_X1 U85969 ( .A1(n81539), .A2(n106178), .B1(n106176), .B2(n107259), 
        .ZN(n97550) );
  OAI21_X1 U85970 ( .B1(n106203), .B2(n106179), .A(n97551), .ZN(
        \DLX_Datapath/RegisterFile/N23814 ) );
  AOI22_X1 U85971 ( .A1(n106178), .A2(n81308), .B1(n74057), .B2(n81339), .ZN(
        n97551) );
  OAI21_X1 U85972 ( .B1(n106180), .B2(n81408), .A(n97552), .ZN(
        \DLX_Datapath/RegisterFile/N23813 ) );
  AOI22_X1 U85973 ( .A1(n94516), .A2(n106178), .B1(n106175), .B2(n108098), 
        .ZN(n97552) );
  OAI21_X1 U85974 ( .B1(n106255), .B2(n106179), .A(n97553), .ZN(
        \DLX_Datapath/RegisterFile/N23812 ) );
  AOI22_X1 U85975 ( .A1(n106177), .A2(n81272), .B1(n106175), .B2(n110797), 
        .ZN(n97553) );
  OAI21_X1 U85976 ( .B1(n106179), .B2(n81629), .A(n97554), .ZN(
        \DLX_Datapath/RegisterFile/N23811 ) );
  AOI22_X1 U85977 ( .A1(n94519), .A2(n106178), .B1(n74338), .B2(n81339), .ZN(
        n97554) );
  OAI21_X1 U85978 ( .B1(n106331), .B2(n106179), .A(n97555), .ZN(
        \DLX_Datapath/RegisterFile/N23810 ) );
  AOI22_X1 U85979 ( .A1(n106177), .A2(n80192), .B1(n106175), .B2(n110490), 
        .ZN(n97555) );
  OAI21_X1 U85980 ( .B1(n106191), .B2(n106179), .A(n97556), .ZN(
        \DLX_Datapath/RegisterFile/N23809 ) );
  AOI22_X1 U85981 ( .A1(n81474), .A2(n81338), .B1(n106175), .B2(n110273), .ZN(
        n97556) );
  OAI21_X1 U85982 ( .B1(n106180), .B2(n106128), .A(n97557), .ZN(
        \DLX_Datapath/RegisterFile/N23808 ) );
  AOI22_X1 U85983 ( .A1(n94523), .A2(n81338), .B1(n106175), .B2(n110591), .ZN(
        n97557) );
  OAI21_X1 U85984 ( .B1(n106186), .B2(n106180), .A(n97558), .ZN(
        \DLX_Datapath/RegisterFile/N23807 ) );
  AOI22_X1 U85985 ( .A1(n106060), .A2(n81338), .B1(n73627), .B2(n81339), .ZN(
        n97558) );
  OAI21_X1 U85986 ( .B1(n106180), .B2(n106106), .A(n97559), .ZN(
        \DLX_Datapath/RegisterFile/N23805 ) );
  AOI22_X1 U85987 ( .A1(n94527), .A2(n81338), .B1(n106175), .B2(n110166), .ZN(
        n97559) );
  OAI21_X1 U85988 ( .B1(n106180), .B2(n81398), .A(n97560), .ZN(
        \DLX_Datapath/RegisterFile/N23803 ) );
  AOI22_X1 U85989 ( .A1(n94530), .A2(n106177), .B1(n106175), .B2(n109833), 
        .ZN(n97560) );
  OAI21_X1 U85990 ( .B1(n106179), .B2(n81451), .A(n97561), .ZN(
        \DLX_Datapath/RegisterFile/N23799 ) );
  AOI22_X1 U85991 ( .A1(n81453), .A2(n106177), .B1(n106175), .B2(n107679), 
        .ZN(n97561) );
  OAI21_X1 U85992 ( .B1(n106200), .B2(n106179), .A(n97562), .ZN(
        \DLX_Datapath/RegisterFile/N23798 ) );
  AOI22_X1 U85993 ( .A1(n105626), .A2(n106177), .B1(n106175), .B2(n109597), 
        .ZN(n97562) );
  OAI21_X1 U85994 ( .B1(n106245), .B2(n106179), .A(n97563), .ZN(
        \DLX_Datapath/RegisterFile/N23797 ) );
  AOI22_X1 U85995 ( .A1(n106177), .A2(n106240), .B1(n106176), .B2(n108558), 
        .ZN(n97563) );
  OAI21_X1 U85996 ( .B1(n106179), .B2(n81394), .A(n97564), .ZN(
        \DLX_Datapath/RegisterFile/N23795 ) );
  AOI22_X1 U85997 ( .A1(n106019), .A2(n106177), .B1(n106176), .B2(n109486), 
        .ZN(n97564) );
  OAI21_X1 U85998 ( .B1(n106010), .B2(n106180), .A(n97565), .ZN(
        \DLX_Datapath/RegisterFile/N23794 ) );
  AOI22_X1 U85999 ( .A1(n94541), .A2(n106177), .B1(n106176), .B2(n109023), 
        .ZN(n97565) );
  OAI21_X1 U86000 ( .B1(n106260), .B2(n106180), .A(n97566), .ZN(
        \DLX_Datapath/RegisterFile/N23793 ) );
  AOI22_X1 U86001 ( .A1(n106178), .A2(n81269), .B1(n106176), .B2(n109371), 
        .ZN(n97566) );
  OAI21_X1 U86002 ( .B1(n106179), .B2(n81509), .A(n97567), .ZN(
        \DLX_Datapath/RegisterFile/N23792 ) );
  AOI22_X1 U86003 ( .A1(n105623), .A2(n106177), .B1(n106176), .B2(n109253), 
        .ZN(n97567) );
  OAI21_X1 U86004 ( .B1(n106179), .B2(n81501), .A(n97568), .ZN(
        \DLX_Datapath/RegisterFile/N23791 ) );
  AOI22_X1 U86005 ( .A1(n105622), .A2(n106177), .B1(n106176), .B2(n109145), 
        .ZN(n97568) );
  OAI21_X1 U86006 ( .B1(n106179), .B2(n81415), .A(n97569), .ZN(
        \DLX_Datapath/RegisterFile/N23790 ) );
  AOI22_X1 U86007 ( .A1(n105621), .A2(n106177), .B1(n106176), .B2(n108680), 
        .ZN(n97569) );
  OAI21_X1 U86008 ( .B1(n106179), .B2(n81498), .A(n97570), .ZN(
        \DLX_Datapath/RegisterFile/N23789 ) );
  AOI22_X1 U86009 ( .A1(n105911), .A2(n106177), .B1(n106176), .B2(n108907), 
        .ZN(n97570) );
  OAI21_X1 U86010 ( .B1(n106268), .B2(n106180), .A(n97571), .ZN(
        \DLX_Datapath/RegisterFile/N23787 ) );
  AOI22_X1 U86011 ( .A1(n106178), .A2(n81265), .B1(n81339), .B2(n107335), .ZN(
        n97571) );
  AOI21_X1 U86012 ( .B1(n97572), .B2(n94258), .A(n97573), .ZN(n81339) );
  NOR2_X1 U86013 ( .A1(n97574), .A2(n104687), .ZN(n81338) );
  NOR2_X1 U86014 ( .A1(n81336), .A2(n105092), .ZN(n97573) );
  NAND2_X1 U86015 ( .A1(n105126), .A2(n94934), .ZN(n81336) );
  OAI21_X1 U86016 ( .B1(n106148), .B2(n105339), .A(n97577), .ZN(
        \DLX_Datapath/RegisterFile/N23786 ) );
  AOI22_X1 U86017 ( .A1(n105337), .A2(n107896), .B1(n105335), .B2(n94559), 
        .ZN(n97577) );
  OAI21_X1 U86018 ( .B1(n105969), .B2(n105339), .A(n97580), .ZN(
        \DLX_Datapath/RegisterFile/N23785 ) );
  AOI22_X1 U86019 ( .A1(n97578), .A2(n107990), .B1(n105335), .B2(n94562), .ZN(
        n97580) );
  OAI21_X1 U86020 ( .B1(n106137), .B2(n105339), .A(n97581), .ZN(
        \DLX_Datapath/RegisterFile/N23784 ) );
  AOI22_X1 U86021 ( .A1(n105337), .A2(n107260), .B1(n105335), .B2(n94564), 
        .ZN(n97581) );
  OAI21_X1 U86022 ( .B1(n106209), .B2(n105339), .A(n97582), .ZN(
        \DLX_Datapath/RegisterFile/N23783 ) );
  AOI22_X1 U86023 ( .A1(n97578), .A2(n107797), .B1(n105335), .B2(n94566), .ZN(
        n97582) );
  OAI21_X1 U86024 ( .B1(n106203), .B2(n105339), .A(n97583), .ZN(
        \DLX_Datapath/RegisterFile/N23782 ) );
  AOI22_X1 U86025 ( .A1(n105337), .A2(n110697), .B1(n105335), .B2(n94568), 
        .ZN(n97583) );
  OAI21_X1 U86026 ( .B1(n106100), .B2(n105339), .A(n97584), .ZN(
        \DLX_Datapath/RegisterFile/N23781 ) );
  AOI22_X1 U86027 ( .A1(n97578), .A2(n108099), .B1(n105335), .B2(n94570), .ZN(
        n97584) );
  OAI21_X1 U86028 ( .B1(n106255), .B2(n105339), .A(n97585), .ZN(
        \DLX_Datapath/RegisterFile/N23780 ) );
  AOI22_X1 U86029 ( .A1(n105337), .A2(n110798), .B1(n105335), .B2(n94572), 
        .ZN(n97585) );
  OAI21_X1 U86030 ( .B1(n105991), .B2(n105339), .A(n97586), .ZN(
        \DLX_Datapath/RegisterFile/N23779 ) );
  AOI22_X1 U86031 ( .A1(n105336), .A2(n110896), .B1(n105335), .B2(n94574), 
        .ZN(n97586) );
  OAI21_X1 U86032 ( .B1(n106331), .B2(n105339), .A(n97587), .ZN(
        \DLX_Datapath/RegisterFile/N23778 ) );
  AOI22_X1 U86033 ( .A1(n105336), .A2(n110491), .B1(n105335), .B2(n94576), 
        .ZN(n97587) );
  OAI21_X1 U86034 ( .B1(n106191), .B2(n105338), .A(n97588), .ZN(
        \DLX_Datapath/RegisterFile/N23777 ) );
  AOI22_X1 U86035 ( .A1(n105336), .A2(n110274), .B1(n105334), .B2(n94578), 
        .ZN(n97588) );
  OAI21_X1 U86036 ( .B1(n106131), .B2(n105338), .A(n97589), .ZN(
        \DLX_Datapath/RegisterFile/N23776 ) );
  AOI22_X1 U86037 ( .A1(n105336), .A2(n110592), .B1(n97579), .B2(n94580), .ZN(
        n97589) );
  OAI21_X1 U86038 ( .B1(n106186), .B2(n105338), .A(n97590), .ZN(
        \DLX_Datapath/RegisterFile/N23775 ) );
  AOI22_X1 U86039 ( .A1(n105336), .A2(n110382), .B1(n105335), .B2(n94582), 
        .ZN(n97590) );
  OAI21_X1 U86040 ( .B1(n106164), .B2(n105338), .A(n97591), .ZN(
        \DLX_Datapath/RegisterFile/N23774 ) );
  AOI22_X1 U86041 ( .A1(n105336), .A2(n110060), .B1(n97579), .B2(n94584), .ZN(
        n97591) );
  OAI21_X1 U86042 ( .B1(n106105), .B2(n105338), .A(n97592), .ZN(
        \DLX_Datapath/RegisterFile/N23773 ) );
  AOI22_X1 U86043 ( .A1(n105336), .A2(n110167), .B1(n97579), .B2(n94586), .ZN(
        n97592) );
  OAI21_X1 U86044 ( .B1(n106219), .B2(n105338), .A(n97593), .ZN(
        \DLX_Datapath/RegisterFile/N23772 ) );
  AOI22_X1 U86045 ( .A1(n105336), .A2(n109951), .B1(n97579), .B2(n94588), .ZN(
        n97593) );
  OAI21_X1 U86046 ( .B1(n106110), .B2(n105338), .A(n97594), .ZN(
        \DLX_Datapath/RegisterFile/N23771 ) );
  AOI22_X1 U86047 ( .A1(n105336), .A2(n109834), .B1(n97579), .B2(n94590), .ZN(
        n97594) );
  OAI21_X1 U86048 ( .B1(n106230), .B2(n105338), .A(n97595), .ZN(
        \DLX_Datapath/RegisterFile/N23770 ) );
  AOI22_X1 U86049 ( .A1(n105336), .A2(n108208), .B1(n105335), .B2(n94592), 
        .ZN(n97595) );
  OAI21_X1 U86050 ( .B1(n106172), .B2(n105338), .A(n97596), .ZN(
        \DLX_Datapath/RegisterFile/N23769 ) );
  AOI22_X1 U86051 ( .A1(n105336), .A2(n108331), .B1(n105335), .B2(n94594), 
        .ZN(n97596) );
  OAI21_X1 U86052 ( .B1(n106237), .B2(n105338), .A(n97597), .ZN(
        \DLX_Datapath/RegisterFile/N23768 ) );
  AOI22_X1 U86053 ( .A1(n105336), .A2(n108442), .B1(n105335), .B2(n94596), 
        .ZN(n97597) );
  OAI21_X1 U86054 ( .B1(n106069), .B2(n105338), .A(n97598), .ZN(
        \DLX_Datapath/RegisterFile/N23767 ) );
  AOI22_X1 U86055 ( .A1(n105336), .A2(n107680), .B1(n97579), .B2(n94598), .ZN(
        n97598) );
  OAI21_X1 U86056 ( .B1(n106199), .B2(n105338), .A(n97599), .ZN(
        \DLX_Datapath/RegisterFile/N23766 ) );
  AOI22_X1 U86057 ( .A1(n97578), .A2(n109598), .B1(n105334), .B2(n94600), .ZN(
        n97599) );
  OAI21_X1 U86058 ( .B1(n106245), .B2(n105339), .A(n97600), .ZN(
        \DLX_Datapath/RegisterFile/N23765 ) );
  AOI22_X1 U86059 ( .A1(n105337), .A2(n108559), .B1(n105334), .B2(n94602), 
        .ZN(n97600) );
  OAI21_X1 U86060 ( .B1(n106159), .B2(n105339), .A(n97601), .ZN(
        \DLX_Datapath/RegisterFile/N23764 ) );
  AOI22_X1 U86061 ( .A1(n97578), .A2(n109703), .B1(n105334), .B2(n94604), .ZN(
        n97601) );
  OAI21_X1 U86062 ( .B1(n106115), .B2(n105338), .A(n97602), .ZN(
        \DLX_Datapath/RegisterFile/N23763 ) );
  AOI22_X1 U86063 ( .A1(n105337), .A2(n109487), .B1(n105334), .B2(n94606), 
        .ZN(n97602) );
  OAI21_X1 U86064 ( .B1(n106010), .B2(n105339), .A(n97603), .ZN(
        \DLX_Datapath/RegisterFile/N23762 ) );
  AOI22_X1 U86065 ( .A1(n97578), .A2(n109024), .B1(n105334), .B2(n94608), .ZN(
        n97603) );
  OAI21_X1 U86066 ( .B1(n106260), .B2(n105339), .A(n97604), .ZN(
        \DLX_Datapath/RegisterFile/N23761 ) );
  AOI22_X1 U86067 ( .A1(n105337), .A2(n109372), .B1(n105334), .B2(n94610), 
        .ZN(n97604) );
  OAI21_X1 U86068 ( .B1(n106044), .B2(n105338), .A(n97605), .ZN(
        \DLX_Datapath/RegisterFile/N23760 ) );
  AOI22_X1 U86069 ( .A1(n97578), .A2(n109254), .B1(n105334), .B2(n94612), .ZN(
        n97605) );
  OAI21_X1 U86070 ( .B1(n106051), .B2(n105339), .A(n97606), .ZN(
        \DLX_Datapath/RegisterFile/N23759 ) );
  AOI22_X1 U86071 ( .A1(n105337), .A2(n109146), .B1(n105334), .B2(n94614), 
        .ZN(n97606) );
  OAI21_X1 U86072 ( .B1(n106095), .B2(n105338), .A(n97607), .ZN(
        \DLX_Datapath/RegisterFile/N23758 ) );
  AOI22_X1 U86073 ( .A1(n97578), .A2(n108681), .B1(n105334), .B2(n94616), .ZN(
        n97607) );
  OAI21_X1 U86074 ( .B1(n106053), .B2(n105339), .A(n97608), .ZN(
        \DLX_Datapath/RegisterFile/N23757 ) );
  AOI22_X1 U86075 ( .A1(n105337), .A2(n108908), .B1(n105334), .B2(n94618), 
        .ZN(n97608) );
  OAI21_X1 U86076 ( .B1(n105217), .B2(n105339), .A(n97609), .ZN(
        \DLX_Datapath/RegisterFile/N23756 ) );
  AOI22_X1 U86077 ( .A1(n105337), .A2(n108796), .B1(n105334), .B2(n94620), 
        .ZN(n97609) );
  OAI21_X1 U86078 ( .B1(n106268), .B2(n105338), .A(n97610), .ZN(
        \DLX_Datapath/RegisterFile/N23755 ) );
  AOI22_X1 U86079 ( .A1(n105337), .A2(n107336), .B1(n105334), .B2(n94622), 
        .ZN(n97610) );
  NOR2_X1 U86080 ( .A1(n97574), .A2(n97611), .ZN(n97579) );
  NOR2_X1 U86081 ( .A1(n97611), .A2(n97612), .ZN(n97578) );
  NOR2_X1 U86082 ( .A1(n97576), .A2(n105095), .ZN(n97611) );
  NAND2_X1 U86083 ( .A1(n94296), .A2(n105125), .ZN(n97576) );
  OAI21_X1 U86084 ( .B1(n106148), .B2(n106144), .A(n97613), .ZN(
        \DLX_Datapath/RegisterFile/N23754 ) );
  AOI22_X1 U86085 ( .A1(n81369), .A2(n107897), .B1(n81521), .B2(n81370), .ZN(
        n97613) );
  OAI21_X1 U86086 ( .B1(n106144), .B2(n81651), .A(n97614), .ZN(
        \DLX_Datapath/RegisterFile/N23753 ) );
  AOI22_X1 U86087 ( .A1(n106143), .A2(n107991), .B1(n81653), .B2(n106141), 
        .ZN(n97614) );
  OAI21_X1 U86088 ( .B1(n106205), .B2(n106144), .A(n97615), .ZN(
        \DLX_Datapath/RegisterFile/N23750 ) );
  AOI22_X1 U86089 ( .A1(n81369), .A2(n110698), .B1(n81428), .B2(n81370), .ZN(
        n97615) );
  OAI21_X1 U86090 ( .B1(n106144), .B2(n106098), .A(n97616), .ZN(
        \DLX_Datapath/RegisterFile/N23749 ) );
  AOI22_X1 U86091 ( .A1(n106143), .A2(n108100), .B1(n81410), .B2(n81370), .ZN(
        n97616) );
  OAI21_X1 U86092 ( .B1(n106255), .B2(n106145), .A(n97617), .ZN(
        \DLX_Datapath/RegisterFile/N23748 ) );
  AOI22_X1 U86093 ( .A1(n81369), .A2(n110799), .B1(n81700), .B2(n106141), .ZN(
        n97617) );
  OAI21_X1 U86094 ( .B1(n106144), .B2(n81629), .A(n97618), .ZN(
        \DLX_Datapath/RegisterFile/N23747 ) );
  AOI22_X1 U86095 ( .A1(n106143), .A2(n110897), .B1(n81632), .B2(n106141), 
        .ZN(n97618) );
  OAI21_X1 U86096 ( .B1(n106331), .B2(n106145), .A(n97619), .ZN(
        \DLX_Datapath/RegisterFile/N23746 ) );
  AOI22_X1 U86097 ( .A1(n81369), .A2(n110492), .B1(n81414), .B2(n106140), .ZN(
        n97619) );
  OAI21_X1 U86098 ( .B1(n106191), .B2(n106145), .A(n97620), .ZN(
        \DLX_Datapath/RegisterFile/N23745 ) );
  AOI22_X1 U86099 ( .A1(n106143), .A2(n110275), .B1(n106140), .B2(n81317), 
        .ZN(n97620) );
  OAI21_X1 U86100 ( .B1(n106145), .B2(n106131), .A(n97621), .ZN(
        \DLX_Datapath/RegisterFile/N23744 ) );
  AOI22_X1 U86101 ( .A1(n81369), .A2(n110593), .B1(n81386), .B2(n81370), .ZN(
        n97621) );
  OAI21_X1 U86102 ( .B1(n106186), .B2(n106145), .A(n97622), .ZN(
        \DLX_Datapath/RegisterFile/N23743 ) );
  AOI22_X1 U86103 ( .A1(n106143), .A2(n110383), .B1(n106141), .B2(n81320), 
        .ZN(n97622) );
  OAI21_X1 U86104 ( .B1(n106164), .B2(n106145), .A(n97623), .ZN(
        \DLX_Datapath/RegisterFile/N23742 ) );
  AOI22_X1 U86105 ( .A1(n81369), .A2(n110061), .B1(n81604), .B2(n106141), .ZN(
        n97623) );
  OAI21_X1 U86106 ( .B1(n106145), .B2(n106103), .A(n97624), .ZN(
        \DLX_Datapath/RegisterFile/N23741 ) );
  AOI22_X1 U86107 ( .A1(n106142), .A2(n110168), .B1(n81405), .B2(n81370), .ZN(
        n97624) );
  OAI21_X1 U86108 ( .B1(n106219), .B2(n106145), .A(n97625), .ZN(
        \DLX_Datapath/RegisterFile/N23740 ) );
  AOI22_X1 U86109 ( .A1(n106142), .A2(n109952), .B1(n81402), .B2(n106140), 
        .ZN(n97625) );
  OAI21_X1 U86110 ( .B1(n106145), .B2(n81398), .A(n97626), .ZN(
        \DLX_Datapath/RegisterFile/N23739 ) );
  AOI22_X1 U86111 ( .A1(n106142), .A2(n109835), .B1(n81400), .B2(n106140), 
        .ZN(n97626) );
  OAI21_X1 U86112 ( .B1(n106145), .B2(n81451), .A(n97627), .ZN(
        \DLX_Datapath/RegisterFile/N23735 ) );
  AOI22_X1 U86113 ( .A1(n106142), .A2(n107681), .B1(n81506), .B2(n81370), .ZN(
        n97627) );
  OAI21_X1 U86114 ( .B1(n106159), .B2(n106145), .A(n97628), .ZN(
        \DLX_Datapath/RegisterFile/N23732 ) );
  AOI22_X1 U86115 ( .A1(n106142), .A2(n109704), .B1(n81425), .B2(n106141), 
        .ZN(n97628) );
  OAI21_X1 U86116 ( .B1(n106144), .B2(n81394), .A(n97629), .ZN(
        \DLX_Datapath/RegisterFile/N23731 ) );
  AOI22_X1 U86117 ( .A1(n106142), .A2(n109488), .B1(n81396), .B2(n81370), .ZN(
        n97629) );
  OAI21_X1 U86118 ( .B1(n106010), .B2(n106145), .A(n97630), .ZN(
        \DLX_Datapath/RegisterFile/N23730 ) );
  AOI22_X1 U86119 ( .A1(n106142), .A2(n109025), .B1(n81590), .B2(n106140), 
        .ZN(n97630) );
  OAI21_X1 U86120 ( .B1(n106260), .B2(n106145), .A(n97631), .ZN(
        \DLX_Datapath/RegisterFile/N23729 ) );
  AOI22_X1 U86121 ( .A1(n106142), .A2(n109373), .B1(n81423), .B2(n106141), 
        .ZN(n97631) );
  OAI21_X1 U86122 ( .B1(n106144), .B2(n81509), .A(n97632), .ZN(
        \DLX_Datapath/RegisterFile/N23728 ) );
  AOI22_X1 U86123 ( .A1(n106142), .A2(n109255), .B1(n81511), .B2(n106141), 
        .ZN(n97632) );
  OAI21_X1 U86124 ( .B1(n106144), .B2(n81501), .A(n97633), .ZN(
        \DLX_Datapath/RegisterFile/N23727 ) );
  AOI22_X1 U86125 ( .A1(n106142), .A2(n109147), .B1(n81503), .B2(n106140), 
        .ZN(n97633) );
  OAI21_X1 U86126 ( .B1(n106145), .B2(n106093), .A(n97634), .ZN(
        \DLX_Datapath/RegisterFile/N23726 ) );
  AOI22_X1 U86127 ( .A1(n106142), .A2(n108682), .B1(n81417), .B2(n81370), .ZN(
        n97634) );
  OAI21_X1 U86128 ( .B1(n106145), .B2(n81498), .A(n97635), .ZN(
        \DLX_Datapath/RegisterFile/N23725 ) );
  AOI22_X1 U86129 ( .A1(n106142), .A2(n108909), .B1(n81500), .B2(n106140), 
        .ZN(n97635) );
  OAI21_X1 U86130 ( .B1(n106268), .B2(n106144), .A(n97636), .ZN(
        \DLX_Datapath/RegisterFile/N23723 ) );
  AOI22_X1 U86131 ( .A1(n106142), .A2(n107337), .B1(n106141), .B2(n81327), 
        .ZN(n97636) );
  NOR2_X1 U86132 ( .A1(n97574), .A2(n97637), .ZN(n81370) );
  NOR2_X1 U86133 ( .A1(n97612), .A2(n97637), .ZN(n81369) );
  NOR2_X1 U86134 ( .A1(n81367), .A2(n105092), .ZN(n97637) );
  NAND2_X1 U86135 ( .A1(n94331), .A2(n105126), .ZN(n81367) );
  OAI21_X1 U86136 ( .B1(n106148), .B2(n105333), .A(n97639), .ZN(
        \DLX_Datapath/RegisterFile/N23722 ) );
  AOI22_X1 U86137 ( .A1(n105332), .A2(n94667), .B1(n105329), .B2(n70358), .ZN(
        n97639) );
  OAI21_X1 U86138 ( .B1(n105969), .B2(n105333), .A(n97642), .ZN(
        \DLX_Datapath/RegisterFile/N23721 ) );
  AOI22_X1 U86139 ( .A1(n105331), .A2(n94670), .B1(n105328), .B2(n70500), .ZN(
        n97642) );
  OAI21_X1 U86140 ( .B1(n106137), .B2(n105333), .A(n97643), .ZN(
        \DLX_Datapath/RegisterFile/N23720 ) );
  AOI22_X1 U86141 ( .A1(n105332), .A2(n94672), .B1(n105329), .B2(n69553), .ZN(
        n97643) );
  OAI21_X1 U86142 ( .B1(n106209), .B2(n105333), .A(n97644), .ZN(
        \DLX_Datapath/RegisterFile/N23719 ) );
  AOI22_X1 U86143 ( .A1(n105331), .A2(n94674), .B1(n105328), .B2(n70214), .ZN(
        n97644) );
  OAI21_X1 U86144 ( .B1(n106203), .B2(n105333), .A(n97645), .ZN(
        \DLX_Datapath/RegisterFile/N23718 ) );
  AOI22_X1 U86145 ( .A1(n105332), .A2(n94676), .B1(n105329), .B2(n74060), .ZN(
        n97645) );
  OAI21_X1 U86146 ( .B1(n106100), .B2(n105333), .A(n97646), .ZN(
        \DLX_Datapath/RegisterFile/N23717 ) );
  AOI22_X1 U86147 ( .A1(n105331), .A2(n94678), .B1(n105328), .B2(n70647), .ZN(
        n97646) );
  OAI21_X1 U86148 ( .B1(n106255), .B2(n105333), .A(n97647), .ZN(
        \DLX_Datapath/RegisterFile/N23716 ) );
  AOI22_X1 U86149 ( .A1(n105332), .A2(n94680), .B1(n105329), .B2(n74201), .ZN(
        n97647) );
  OAI21_X1 U86150 ( .B1(n81629), .B2(n105333), .A(n97648), .ZN(
        \DLX_Datapath/RegisterFile/N23715 ) );
  AOI22_X1 U86151 ( .A1(n105331), .A2(n94682), .B1(n105328), .B2(n74341), .ZN(
        n97648) );
  OAI21_X1 U86152 ( .B1(n106331), .B2(n105333), .A(n97649), .ZN(
        \DLX_Datapath/RegisterFile/N23714 ) );
  AOI22_X1 U86153 ( .A1(n105331), .A2(n94684), .B1(n105328), .B2(n73777), .ZN(
        n97649) );
  OAI21_X1 U86154 ( .B1(n106191), .B2(n105333), .A(n97650), .ZN(
        \DLX_Datapath/RegisterFile/N23713 ) );
  AOI22_X1 U86155 ( .A1(n105330), .A2(n94686), .B1(n105327), .B2(n73481), .ZN(
        n97650) );
  OAI21_X1 U86156 ( .B1(n106131), .B2(n105333), .A(n97651), .ZN(
        \DLX_Datapath/RegisterFile/N23712 ) );
  AOI22_X1 U86157 ( .A1(n105330), .A2(n94688), .B1(n105327), .B2(n73918), .ZN(
        n97651) );
  OAI21_X1 U86158 ( .B1(n106186), .B2(n105333), .A(n97652), .ZN(
        \DLX_Datapath/RegisterFile/N23711 ) );
  AOI22_X1 U86159 ( .A1(n105330), .A2(n94690), .B1(n105327), .B2(n73630), .ZN(
        n97652) );
  OAI21_X1 U86160 ( .B1(n106164), .B2(n105333), .A(n97653), .ZN(
        \DLX_Datapath/RegisterFile/N23710 ) );
  AOI22_X1 U86161 ( .A1(n105330), .A2(n94692), .B1(n105327), .B2(n73192), .ZN(
        n97653) );
  OAI21_X1 U86162 ( .B1(n106105), .B2(n105333), .A(n97654), .ZN(
        \DLX_Datapath/RegisterFile/N23709 ) );
  AOI22_X1 U86163 ( .A1(n105330), .A2(n94694), .B1(n105327), .B2(n73334), .ZN(
        n97654) );
  OAI21_X1 U86164 ( .B1(n106219), .B2(n105333), .A(n97655), .ZN(
        \DLX_Datapath/RegisterFile/N23708 ) );
  AOI22_X1 U86165 ( .A1(n105330), .A2(n94696), .B1(n105327), .B2(n73050), .ZN(
        n97655) );
  OAI21_X1 U86166 ( .B1(n106110), .B2(n105333), .A(n97656), .ZN(
        \DLX_Datapath/RegisterFile/N23707 ) );
  AOI22_X1 U86167 ( .A1(n105330), .A2(n94698), .B1(n105327), .B2(n72900), .ZN(
        n97656) );
  OAI21_X1 U86168 ( .B1(n106232), .B2(n105333), .A(n97657), .ZN(
        \DLX_Datapath/RegisterFile/N23706 ) );
  AOI22_X1 U86169 ( .A1(n105330), .A2(n94700), .B1(n105327), .B2(n70796), .ZN(
        n97657) );
  OAI21_X1 U86170 ( .B1(n106172), .B2(n105333), .A(n97658), .ZN(
        \DLX_Datapath/RegisterFile/N23705 ) );
  AOI22_X1 U86171 ( .A1(n105330), .A2(n94702), .B1(n105327), .B2(n70955), .ZN(
        n97658) );
  OAI21_X1 U86172 ( .B1(n106237), .B2(n105333), .A(n97659), .ZN(
        \DLX_Datapath/RegisterFile/N23704 ) );
  AOI22_X1 U86173 ( .A1(n105330), .A2(n94704), .B1(n105327), .B2(n71100), .ZN(
        n97659) );
  OAI21_X1 U86174 ( .B1(n106069), .B2(n105333), .A(n97660), .ZN(
        \DLX_Datapath/RegisterFile/N23703 ) );
  AOI22_X1 U86175 ( .A1(n105330), .A2(n94706), .B1(n105327), .B2(n70061), .ZN(
        n97660) );
  OAI21_X1 U86176 ( .B1(n106197), .B2(n105333), .A(n97661), .ZN(
        \DLX_Datapath/RegisterFile/N23702 ) );
  AOI22_X1 U86177 ( .A1(n105331), .A2(n94708), .B1(n105328), .B2(n72590), .ZN(
        n97661) );
  OAI21_X1 U86178 ( .B1(n106246), .B2(n97638), .A(n97662), .ZN(
        \DLX_Datapath/RegisterFile/N23701 ) );
  AOI22_X1 U86179 ( .A1(n105332), .A2(n94710), .B1(n105329), .B2(n71249), .ZN(
        n97662) );
  OAI21_X1 U86180 ( .B1(n106159), .B2(n97638), .A(n97663), .ZN(
        \DLX_Datapath/RegisterFile/N23700 ) );
  AOI22_X1 U86181 ( .A1(n105331), .A2(n94712), .B1(n105328), .B2(n72732), .ZN(
        n97663) );
  OAI21_X1 U86182 ( .B1(n106115), .B2(n97638), .A(n97664), .ZN(
        \DLX_Datapath/RegisterFile/N23699 ) );
  AOI22_X1 U86183 ( .A1(n105332), .A2(n94714), .B1(n105329), .B2(n72442), .ZN(
        n97664) );
  OAI21_X1 U86184 ( .B1(n106010), .B2(n97638), .A(n97665), .ZN(
        \DLX_Datapath/RegisterFile/N23698 ) );
  AOI22_X1 U86185 ( .A1(n105331), .A2(n81259), .B1(n105328), .B2(n71842), .ZN(
        n97665) );
  OAI21_X1 U86186 ( .B1(n106260), .B2(n97638), .A(n97666), .ZN(
        \DLX_Datapath/RegisterFile/N23697 ) );
  AOI22_X1 U86187 ( .A1(n105332), .A2(n94717), .B1(n105329), .B2(n72291), .ZN(
        n97666) );
  OAI21_X1 U86188 ( .B1(n106045), .B2(n97638), .A(n97667), .ZN(
        \DLX_Datapath/RegisterFile/N23696 ) );
  AOI22_X1 U86189 ( .A1(n105331), .A2(n94719), .B1(n105328), .B2(n72140), .ZN(
        n97667) );
  OAI21_X1 U86190 ( .B1(n106050), .B2(n97638), .A(n97668), .ZN(
        \DLX_Datapath/RegisterFile/N23695 ) );
  AOI22_X1 U86191 ( .A1(n105332), .A2(n94721), .B1(n105329), .B2(n71996), .ZN(
        n97668) );
  OAI21_X1 U86192 ( .B1(n106095), .B2(n97638), .A(n97669), .ZN(
        \DLX_Datapath/RegisterFile/N23694 ) );
  AOI22_X1 U86193 ( .A1(n105331), .A2(n94723), .B1(n105328), .B2(n71398), .ZN(
        n97669) );
  OAI21_X1 U86194 ( .B1(n106055), .B2(n97638), .A(n97670), .ZN(
        \DLX_Datapath/RegisterFile/N23693 ) );
  AOI22_X1 U86195 ( .A1(n105332), .A2(n94725), .B1(n105329), .B2(n71693), .ZN(
        n97670) );
  OAI21_X1 U86196 ( .B1(n105217), .B2(n105333), .A(n97671), .ZN(
        \DLX_Datapath/RegisterFile/N23692 ) );
  AOI22_X1 U86197 ( .A1(n105332), .A2(n94727), .B1(n105329), .B2(n71549), .ZN(
        n97671) );
  OAI21_X1 U86198 ( .B1(n106268), .B2(n105333), .A(n97672), .ZN(
        \DLX_Datapath/RegisterFile/N23691 ) );
  AOI22_X1 U86199 ( .A1(n105331), .A2(n94729), .B1(n105328), .B2(n69658), .ZN(
        n97672) );
  NOR2_X1 U86200 ( .A1(n97612), .A2(n97673), .ZN(n97641) );
  AOI21_X1 U86201 ( .B1(n105205), .B2(n97574), .A(n105601), .ZN(n97612) );
  NOR2_X1 U86203 ( .A1(n97638), .A2(n105094), .ZN(n97673) );
  OR2_X1 U86204 ( .A1(n97674), .A2(n94999), .ZN(n97574) );
  NAND2_X1 U86205 ( .A1(n94367), .A2(n105125), .ZN(n97638) );
  OAI21_X1 U86206 ( .B1(n106148), .B2(n105326), .A(n97676), .ZN(
        \DLX_Datapath/RegisterFile/N23690 ) );
  AOI22_X1 U86207 ( .A1(n105324), .A2(n107898), .B1(n105321), .B2(n81360), 
        .ZN(n97676) );
  OAI21_X1 U86208 ( .B1(n105969), .B2(n105326), .A(n97679), .ZN(
        \DLX_Datapath/RegisterFile/N23689 ) );
  AOI22_X1 U86209 ( .A1(n105325), .A2(n107992), .B1(n105322), .B2(n94511), 
        .ZN(n97679) );
  OAI21_X1 U86210 ( .B1(n106137), .B2(n105326), .A(n97680), .ZN(
        \DLX_Datapath/RegisterFile/N23688 ) );
  AOI22_X1 U86211 ( .A1(n105325), .A2(n107262), .B1(n105322), .B2(n81539), 
        .ZN(n97680) );
  OAI21_X1 U86212 ( .B1(n106209), .B2(n105326), .A(n97681), .ZN(
        \DLX_Datapath/RegisterFile/N23687 ) );
  AOI22_X1 U86213 ( .A1(n105324), .A2(n107799), .B1(n105321), .B2(n81301), 
        .ZN(n97681) );
  OAI21_X1 U86214 ( .B1(n106205), .B2(n105326), .A(n97682), .ZN(
        \DLX_Datapath/RegisterFile/N23686 ) );
  AOI22_X1 U86215 ( .A1(n105325), .A2(n74061), .B1(n105322), .B2(n81308), .ZN(
        n97682) );
  OAI21_X1 U86216 ( .B1(n106100), .B2(n105326), .A(n97683), .ZN(
        \DLX_Datapath/RegisterFile/N23685 ) );
  AOI22_X1 U86217 ( .A1(n105324), .A2(n108101), .B1(n105321), .B2(n94516), 
        .ZN(n97683) );
  OAI21_X1 U86218 ( .B1(n106255), .B2(n105326), .A(n97684), .ZN(
        \DLX_Datapath/RegisterFile/N23684 ) );
  AOI22_X1 U86219 ( .A1(n105324), .A2(n110800), .B1(n105321), .B2(n81272), 
        .ZN(n97684) );
  OAI21_X1 U86220 ( .B1(n105990), .B2(n105326), .A(n97685), .ZN(
        \DLX_Datapath/RegisterFile/N23683 ) );
  AOI22_X1 U86221 ( .A1(n105325), .A2(n74342), .B1(n105322), .B2(n94519), .ZN(
        n97685) );
  OAI21_X1 U86222 ( .B1(n106331), .B2(n105326), .A(n97686), .ZN(
        \DLX_Datapath/RegisterFile/N23682 ) );
  AOI22_X1 U86223 ( .A1(n105324), .A2(n110493), .B1(n105322), .B2(n80192), 
        .ZN(n97686) );
  OAI21_X1 U86224 ( .B1(n106191), .B2(n105326), .A(n97687), .ZN(
        \DLX_Datapath/RegisterFile/N23681 ) );
  AOI22_X1 U86225 ( .A1(n105323), .A2(n110276), .B1(n105320), .B2(n81474), 
        .ZN(n97687) );
  OAI21_X1 U86226 ( .B1(n106128), .B2(n105326), .A(n97688), .ZN(
        \DLX_Datapath/RegisterFile/N23680 ) );
  AOI22_X1 U86227 ( .A1(n105323), .A2(n110594), .B1(n105320), .B2(n94523), 
        .ZN(n97688) );
  OAI21_X1 U86228 ( .B1(n106186), .B2(n105326), .A(n97689), .ZN(
        \DLX_Datapath/RegisterFile/N23679 ) );
  AOI22_X1 U86229 ( .A1(n105323), .A2(n110384), .B1(n105320), .B2(n106061), 
        .ZN(n97689) );
  OAI21_X1 U86230 ( .B1(n106164), .B2(n105326), .A(n97690), .ZN(
        \DLX_Datapath/RegisterFile/N23678 ) );
  AOI22_X1 U86231 ( .A1(n105323), .A2(n110062), .B1(n105320), .B2(n81347), 
        .ZN(n97690) );
  OAI21_X1 U86232 ( .B1(n106105), .B2(n97675), .A(n97691), .ZN(
        \DLX_Datapath/RegisterFile/N23677 ) );
  AOI22_X1 U86233 ( .A1(n105323), .A2(n110169), .B1(n105320), .B2(n94527), 
        .ZN(n97691) );
  OAI21_X1 U86234 ( .B1(n106219), .B2(n97675), .A(n97692), .ZN(
        \DLX_Datapath/RegisterFile/N23676 ) );
  AOI22_X1 U86235 ( .A1(n105323), .A2(n109953), .B1(n105321), .B2(n81297), 
        .ZN(n97692) );
  OAI21_X1 U86236 ( .B1(n106110), .B2(n97675), .A(n97693), .ZN(
        \DLX_Datapath/RegisterFile/N23675 ) );
  AOI22_X1 U86237 ( .A1(n105323), .A2(n109836), .B1(n105320), .B2(n94530), 
        .ZN(n97693) );
  OAI21_X1 U86238 ( .B1(n106232), .B2(n97675), .A(n97694), .ZN(
        \DLX_Datapath/RegisterFile/N23674 ) );
  AOI22_X1 U86239 ( .A1(n105323), .A2(n108210), .B1(n105320), .B2(n81286), 
        .ZN(n97694) );
  OAI21_X1 U86240 ( .B1(n106172), .B2(n97675), .A(n97695), .ZN(
        \DLX_Datapath/RegisterFile/N23673 ) );
  AOI22_X1 U86241 ( .A1(n105323), .A2(n108333), .B1(n105320), .B2(n106168), 
        .ZN(n97695) );
  OAI21_X1 U86242 ( .B1(n106237), .B2(n97675), .A(n97696), .ZN(
        \DLX_Datapath/RegisterFile/N23672 ) );
  AOI22_X1 U86243 ( .A1(n105323), .A2(n108444), .B1(n105320), .B2(n81283), 
        .ZN(n97696) );
  OAI21_X1 U86244 ( .B1(n106069), .B2(n97675), .A(n97697), .ZN(
        \DLX_Datapath/RegisterFile/N23671 ) );
  AOI22_X1 U86245 ( .A1(n105323), .A2(n107682), .B1(n105320), .B2(n81453), 
        .ZN(n97697) );
  OAI21_X1 U86246 ( .B1(n106198), .B2(n97675), .A(n97698), .ZN(
        \DLX_Datapath/RegisterFile/N23670 ) );
  AOI22_X1 U86247 ( .A1(n105324), .A2(n109600), .B1(n105322), .B2(n94536), 
        .ZN(n97698) );
  OAI21_X1 U86248 ( .B1(n106246), .B2(n105326), .A(n97699), .ZN(
        \DLX_Datapath/RegisterFile/N23669 ) );
  AOI22_X1 U86249 ( .A1(n105325), .A2(n108561), .B1(n105322), .B2(n106241), 
        .ZN(n97699) );
  OAI21_X1 U86250 ( .B1(n106159), .B2(n105326), .A(n97700), .ZN(
        \DLX_Datapath/RegisterFile/N23668 ) );
  AOI22_X1 U86251 ( .A1(n105324), .A2(n109705), .B1(n105321), .B2(n81351), 
        .ZN(n97700) );
  OAI21_X1 U86252 ( .B1(n106115), .B2(n105326), .A(n97701), .ZN(
        \DLX_Datapath/RegisterFile/N23667 ) );
  AOI22_X1 U86253 ( .A1(n105325), .A2(n109489), .B1(n105322), .B2(n106020), 
        .ZN(n97701) );
  OAI21_X1 U86254 ( .B1(n106010), .B2(n105326), .A(n97702), .ZN(
        \DLX_Datapath/RegisterFile/N23666 ) );
  AOI22_X1 U86255 ( .A1(n105324), .A2(n109026), .B1(n105321), .B2(n94541), 
        .ZN(n97702) );
  OAI21_X1 U86256 ( .B1(n106261), .B2(n105326), .A(n97703), .ZN(
        \DLX_Datapath/RegisterFile/N23665 ) );
  AOI22_X1 U86257 ( .A1(n105325), .A2(n109374), .B1(n105321), .B2(n81269), 
        .ZN(n97703) );
  OAI21_X1 U86258 ( .B1(n106045), .B2(n105326), .A(n97704), .ZN(
        \DLX_Datapath/RegisterFile/N23664 ) );
  AOI22_X1 U86259 ( .A1(n105324), .A2(n109256), .B1(n105322), .B2(n105624), 
        .ZN(n97704) );
  OAI21_X1 U86260 ( .B1(n106050), .B2(n105326), .A(n97705), .ZN(
        \DLX_Datapath/RegisterFile/N23663 ) );
  AOI22_X1 U86261 ( .A1(n105325), .A2(n71997), .B1(n105321), .B2(n94546), .ZN(
        n97705) );
  OAI21_X1 U86262 ( .B1(n106095), .B2(n105326), .A(n97706), .ZN(
        \DLX_Datapath/RegisterFile/N23662 ) );
  AOI22_X1 U86263 ( .A1(n105324), .A2(n108683), .B1(n105322), .B2(n94548), 
        .ZN(n97706) );
  OAI21_X1 U86264 ( .B1(n106055), .B2(n105326), .A(n97707), .ZN(
        \DLX_Datapath/RegisterFile/N23661 ) );
  AOI22_X1 U86265 ( .A1(n105325), .A2(n108910), .B1(n105322), .B2(n81783), 
        .ZN(n97707) );
  OAI21_X1 U86266 ( .B1(n105217), .B2(n105326), .A(n97708), .ZN(
        \DLX_Datapath/RegisterFile/N23660 ) );
  AOI22_X1 U86267 ( .A1(n105325), .A2(n108798), .B1(n105321), .B2(n80188), 
        .ZN(n97708) );
  OAI21_X1 U86268 ( .B1(n106268), .B2(n105326), .A(n97709), .ZN(
        \DLX_Datapath/RegisterFile/N23659 ) );
  AOI22_X1 U86269 ( .A1(n105324), .A2(n107338), .B1(n105321), .B2(n81265), 
        .ZN(n97709) );
  AOI21_X1 U86271 ( .B1(n97572), .B2(n94398), .A(n97711), .ZN(n97677) );
  NOR2_X1 U86272 ( .A1(n97675), .A2(n105090), .ZN(n97711) );
  NAND2_X1 U86273 ( .A1(n105125), .A2(n94399), .ZN(n97675) );
  OAI21_X1 U86274 ( .B1(n106148), .B2(n105319), .A(n97713), .ZN(
        \DLX_Datapath/RegisterFile/N23658 ) );
  AOI22_X1 U86275 ( .A1(n105317), .A2(n70360), .B1(n105315), .B2(n94559), .ZN(
        n97713) );
  OAI21_X1 U86276 ( .B1(n105969), .B2(n105319), .A(n97716), .ZN(
        \DLX_Datapath/RegisterFile/N23657 ) );
  AOI22_X1 U86277 ( .A1(n105316), .A2(n70502), .B1(n105315), .B2(n94562), .ZN(
        n97716) );
  OAI21_X1 U86278 ( .B1(n106137), .B2(n105319), .A(n97717), .ZN(
        \DLX_Datapath/RegisterFile/N23656 ) );
  AOI22_X1 U86279 ( .A1(n105317), .A2(n69555), .B1(n105315), .B2(n94564), .ZN(
        n97717) );
  OAI21_X1 U86280 ( .B1(n106209), .B2(n105319), .A(n97718), .ZN(
        \DLX_Datapath/RegisterFile/N23655 ) );
  AOI22_X1 U86281 ( .A1(n105316), .A2(n70216), .B1(n105315), .B2(n94566), .ZN(
        n97718) );
  OAI21_X1 U86282 ( .B1(n106204), .B2(n105319), .A(n97719), .ZN(
        \DLX_Datapath/RegisterFile/N23654 ) );
  AOI22_X1 U86283 ( .A1(n105317), .A2(n74062), .B1(n105315), .B2(n94568), .ZN(
        n97719) );
  OAI21_X1 U86284 ( .B1(n106100), .B2(n105319), .A(n97720), .ZN(
        \DLX_Datapath/RegisterFile/N23653 ) );
  AOI22_X1 U86285 ( .A1(n105316), .A2(n70649), .B1(n105315), .B2(n94570), .ZN(
        n97720) );
  OAI21_X1 U86286 ( .B1(n106255), .B2(n105319), .A(n97721), .ZN(
        \DLX_Datapath/RegisterFile/N23652 ) );
  AOI22_X1 U86287 ( .A1(n105317), .A2(n74203), .B1(n105315), .B2(n94572), .ZN(
        n97721) );
  OAI21_X1 U86288 ( .B1(n105992), .B2(n105319), .A(n97722), .ZN(
        \DLX_Datapath/RegisterFile/N23651 ) );
  AOI22_X1 U86289 ( .A1(n105316), .A2(n74343), .B1(n105315), .B2(n94574), .ZN(
        n97722) );
  OAI21_X1 U86290 ( .B1(n106331), .B2(n105319), .A(n97723), .ZN(
        \DLX_Datapath/RegisterFile/N23650 ) );
  AOI22_X1 U86291 ( .A1(n105316), .A2(n73779), .B1(n105315), .B2(n94576), .ZN(
        n97723) );
  OAI21_X1 U86292 ( .B1(n106191), .B2(n105318), .A(n97724), .ZN(
        \DLX_Datapath/RegisterFile/N23649 ) );
  AOI22_X1 U86293 ( .A1(n97714), .A2(n73483), .B1(n105315), .B2(n94578), .ZN(
        n97724) );
  OAI21_X1 U86294 ( .B1(n106129), .B2(n105318), .A(n97725), .ZN(
        \DLX_Datapath/RegisterFile/N23648 ) );
  AOI22_X1 U86295 ( .A1(n97714), .A2(n73920), .B1(n105314), .B2(n94580), .ZN(
        n97725) );
  OAI21_X1 U86296 ( .B1(n106187), .B2(n105318), .A(n97726), .ZN(
        \DLX_Datapath/RegisterFile/N23647 ) );
  AOI22_X1 U86297 ( .A1(n97714), .A2(n73632), .B1(n97715), .B2(n94582), .ZN(
        n97726) );
  OAI21_X1 U86298 ( .B1(n106164), .B2(n105318), .A(n97727), .ZN(
        \DLX_Datapath/RegisterFile/N23646 ) );
  AOI22_X1 U86299 ( .A1(n97714), .A2(n73194), .B1(n105315), .B2(n94584), .ZN(
        n97727) );
  OAI21_X1 U86300 ( .B1(n106105), .B2(n105318), .A(n97728), .ZN(
        \DLX_Datapath/RegisterFile/N23645 ) );
  AOI22_X1 U86301 ( .A1(n105316), .A2(n73336), .B1(n97715), .B2(n94586), .ZN(
        n97728) );
  OAI21_X1 U86302 ( .B1(n106219), .B2(n105318), .A(n97729), .ZN(
        \DLX_Datapath/RegisterFile/N23644 ) );
  AOI22_X1 U86303 ( .A1(n97714), .A2(n73052), .B1(n97715), .B2(n94588), .ZN(
        n97729) );
  OAI21_X1 U86304 ( .B1(n106110), .B2(n105318), .A(n97730), .ZN(
        \DLX_Datapath/RegisterFile/N23643 ) );
  AOI22_X1 U86305 ( .A1(n97714), .A2(n72902), .B1(n97715), .B2(n94590), .ZN(
        n97730) );
  OAI21_X1 U86306 ( .B1(n106232), .B2(n105318), .A(n97731), .ZN(
        \DLX_Datapath/RegisterFile/N23642 ) );
  AOI22_X1 U86307 ( .A1(n97714), .A2(n70798), .B1(n97715), .B2(n94592), .ZN(
        n97731) );
  OAI21_X1 U86308 ( .B1(n106172), .B2(n105318), .A(n97732), .ZN(
        \DLX_Datapath/RegisterFile/N23641 ) );
  AOI22_X1 U86309 ( .A1(n105317), .A2(n70957), .B1(n105315), .B2(n94594), .ZN(
        n97732) );
  OAI21_X1 U86310 ( .B1(n106237), .B2(n105318), .A(n97733), .ZN(
        \DLX_Datapath/RegisterFile/N23640 ) );
  AOI22_X1 U86311 ( .A1(n105316), .A2(n71102), .B1(n105315), .B2(n94596), .ZN(
        n97733) );
  OAI21_X1 U86312 ( .B1(n106069), .B2(n105318), .A(n97734), .ZN(
        \DLX_Datapath/RegisterFile/N23639 ) );
  AOI22_X1 U86313 ( .A1(n97714), .A2(n70063), .B1(n97715), .B2(n94598), .ZN(
        n97734) );
  OAI21_X1 U86314 ( .B1(n106200), .B2(n105318), .A(n97735), .ZN(
        \DLX_Datapath/RegisterFile/N23638 ) );
  AOI22_X1 U86315 ( .A1(n105316), .A2(n72592), .B1(n105314), .B2(n94600), .ZN(
        n97735) );
  OAI21_X1 U86316 ( .B1(n106246), .B2(n105319), .A(n97736), .ZN(
        \DLX_Datapath/RegisterFile/N23637 ) );
  AOI22_X1 U86317 ( .A1(n105317), .A2(n71251), .B1(n105314), .B2(n94602), .ZN(
        n97736) );
  OAI21_X1 U86318 ( .B1(n106159), .B2(n105319), .A(n97737), .ZN(
        \DLX_Datapath/RegisterFile/N23636 ) );
  AOI22_X1 U86319 ( .A1(n105316), .A2(n72734), .B1(n105314), .B2(n94604), .ZN(
        n97737) );
  OAI21_X1 U86320 ( .B1(n106115), .B2(n105318), .A(n97738), .ZN(
        \DLX_Datapath/RegisterFile/N23635 ) );
  AOI22_X1 U86321 ( .A1(n105317), .A2(n72444), .B1(n105314), .B2(n94606), .ZN(
        n97738) );
  OAI21_X1 U86322 ( .B1(n106010), .B2(n105319), .A(n97739), .ZN(
        \DLX_Datapath/RegisterFile/N23634 ) );
  AOI22_X1 U86323 ( .A1(n105316), .A2(n71844), .B1(n105314), .B2(n94608), .ZN(
        n97739) );
  OAI21_X1 U86324 ( .B1(n106261), .B2(n105319), .A(n97740), .ZN(
        \DLX_Datapath/RegisterFile/N23633 ) );
  AOI22_X1 U86325 ( .A1(n105317), .A2(n72293), .B1(n105314), .B2(n94610), .ZN(
        n97740) );
  OAI21_X1 U86326 ( .B1(n106045), .B2(n105318), .A(n97741), .ZN(
        \DLX_Datapath/RegisterFile/N23632 ) );
  AOI22_X1 U86327 ( .A1(n105316), .A2(n72142), .B1(n105314), .B2(n94612), .ZN(
        n97741) );
  OAI21_X1 U86328 ( .B1(n106050), .B2(n105319), .A(n97742), .ZN(
        \DLX_Datapath/RegisterFile/N23631 ) );
  AOI22_X1 U86329 ( .A1(n105317), .A2(n71998), .B1(n105314), .B2(n94614), .ZN(
        n97742) );
  OAI21_X1 U86330 ( .B1(n106095), .B2(n105318), .A(n97743), .ZN(
        \DLX_Datapath/RegisterFile/N23630 ) );
  AOI22_X1 U86331 ( .A1(n105316), .A2(n71400), .B1(n105314), .B2(n94616), .ZN(
        n97743) );
  OAI21_X1 U86332 ( .B1(n106055), .B2(n105319), .A(n97744), .ZN(
        \DLX_Datapath/RegisterFile/N23629 ) );
  AOI22_X1 U86333 ( .A1(n105317), .A2(n71695), .B1(n105314), .B2(n94618), .ZN(
        n97744) );
  OAI21_X1 U86334 ( .B1(n105217), .B2(n105319), .A(n97745), .ZN(
        \DLX_Datapath/RegisterFile/N23628 ) );
  AOI22_X1 U86335 ( .A1(n105317), .A2(n71551), .B1(n105314), .B2(n94620), .ZN(
        n97745) );
  OAI21_X1 U86336 ( .B1(n106268), .B2(n105318), .A(n97746), .ZN(
        \DLX_Datapath/RegisterFile/N23627 ) );
  AOI22_X1 U86337 ( .A1(n105316), .A2(n69660), .B1(n105314), .B2(n94622), .ZN(
        n97746) );
  NOR2_X1 U86338 ( .A1(n97710), .A2(n97747), .ZN(n97715) );
  NOR2_X1 U86339 ( .A1(n97747), .A2(n97748), .ZN(n97714) );
  NOR2_X1 U86340 ( .A1(n97712), .A2(n105092), .ZN(n97747) );
  NAND2_X1 U86341 ( .A1(n94434), .A2(n105126), .ZN(n97712) );
  OAI21_X1 U86342 ( .B1(n106148), .B2(n106134), .A(n97749), .ZN(
        \DLX_Datapath/RegisterFile/N23626 ) );
  AOI22_X1 U86343 ( .A1(n81521), .A2(n106127), .B1(n81387), .B2(n107899), .ZN(
        n97749) );
  OAI21_X1 U86344 ( .B1(n106133), .B2(n105968), .A(n97750), .ZN(
        \DLX_Datapath/RegisterFile/N23625 ) );
  AOI22_X1 U86345 ( .A1(n81653), .A2(n106127), .B1(n81387), .B2(n107993), .ZN(
        n97750) );
  OAI21_X1 U86346 ( .B1(n106137), .B2(n106134), .A(n97751), .ZN(
        \DLX_Datapath/RegisterFile/N23624 ) );
  AOI22_X1 U86347 ( .A1(n106126), .A2(n81380), .B1(n81387), .B2(n107263), .ZN(
        n97751) );
  OAI21_X1 U86348 ( .B1(n106210), .B2(n106134), .A(n97752), .ZN(
        \DLX_Datapath/RegisterFile/N23623 ) );
  AOI22_X1 U86349 ( .A1(n106127), .A2(n81377), .B1(n81387), .B2(n107800), .ZN(
        n97752) );
  OAI21_X1 U86350 ( .B1(n106206), .B2(n106134), .A(n97753), .ZN(
        \DLX_Datapath/RegisterFile/N23622 ) );
  AOI22_X1 U86351 ( .A1(n81428), .A2(n106126), .B1(n81387), .B2(n110699), .ZN(
        n97753) );
  OAI21_X1 U86352 ( .B1(n106134), .B2(n81408), .A(n97754), .ZN(
        \DLX_Datapath/RegisterFile/N23621 ) );
  AOI22_X1 U86353 ( .A1(n81410), .A2(n106127), .B1(n106125), .B2(n108102), 
        .ZN(n97754) );
  OAI21_X1 U86354 ( .B1(n106255), .B2(n106134), .A(n97755), .ZN(
        \DLX_Datapath/RegisterFile/N23620 ) );
  AOI22_X1 U86355 ( .A1(n81700), .A2(n81385), .B1(n81387), .B2(n110801), .ZN(
        n97755) );
  OAI21_X1 U86356 ( .B1(n106134), .B2(n81629), .A(n97756), .ZN(
        \DLX_Datapath/RegisterFile/N23619 ) );
  AOI22_X1 U86357 ( .A1(n81632), .A2(n106126), .B1(n106125), .B2(n110898), 
        .ZN(n97756) );
  OAI21_X1 U86358 ( .B1(n106331), .B2(n106134), .A(n97757), .ZN(
        \DLX_Datapath/RegisterFile/N23618 ) );
  AOI22_X1 U86359 ( .A1(n81414), .A2(n106126), .B1(n73780), .B2(n106125), .ZN(
        n97757) );
  OAI21_X1 U86360 ( .B1(n106191), .B2(n106133), .A(n97758), .ZN(
        \DLX_Datapath/RegisterFile/N23617 ) );
  AOI22_X1 U86361 ( .A1(n106126), .A2(n81317), .B1(n73484), .B2(n106125), .ZN(
        n97758) );
  OAI21_X1 U86362 ( .B1(n106187), .B2(n106133), .A(n97759), .ZN(
        \DLX_Datapath/RegisterFile/N23615 ) );
  AOI22_X1 U86363 ( .A1(n106127), .A2(n81320), .B1(n81387), .B2(n110385), .ZN(
        n97759) );
  OAI21_X1 U86364 ( .B1(n106164), .B2(n106134), .A(n97760), .ZN(
        \DLX_Datapath/RegisterFile/N23614 ) );
  AOI22_X1 U86365 ( .A1(n81604), .A2(n106127), .B1(n106124), .B2(n110063), 
        .ZN(n97760) );
  OAI21_X1 U86366 ( .B1(n106133), .B2(n106104), .A(n97761), .ZN(
        \DLX_Datapath/RegisterFile/N23613 ) );
  AOI22_X1 U86367 ( .A1(n81405), .A2(n81385), .B1(n106124), .B2(n110170), .ZN(
        n97761) );
  OAI21_X1 U86368 ( .B1(n106219), .B2(n106133), .A(n97762), .ZN(
        \DLX_Datapath/RegisterFile/N23612 ) );
  AOI22_X1 U86369 ( .A1(n81402), .A2(n81385), .B1(n106124), .B2(n109954), .ZN(
        n97762) );
  OAI21_X1 U86370 ( .B1(n106134), .B2(n106111), .A(n97763), .ZN(
        \DLX_Datapath/RegisterFile/N23611 ) );
  AOI22_X1 U86371 ( .A1(n81400), .A2(n106127), .B1(n106124), .B2(n109837), 
        .ZN(n97763) );
  OAI21_X1 U86372 ( .B1(n106232), .B2(n106133), .A(n97764), .ZN(
        \DLX_Datapath/RegisterFile/N23610 ) );
  AOI22_X1 U86373 ( .A1(n81385), .A2(n81332), .B1(n106124), .B2(n108211), .ZN(
        n97764) );
  OAI21_X1 U86374 ( .B1(n106173), .B2(n106133), .A(n97765), .ZN(
        \DLX_Datapath/RegisterFile/N23609 ) );
  AOI22_X1 U86375 ( .A1(n106126), .A2(n81373), .B1(n106124), .B2(n108334), 
        .ZN(n97765) );
  OAI21_X1 U86376 ( .B1(n106237), .B2(n106133), .A(n97766), .ZN(
        \DLX_Datapath/RegisterFile/N23608 ) );
  AOI22_X1 U86377 ( .A1(n106127), .A2(n81322), .B1(n106124), .B2(n108445), 
        .ZN(n97766) );
  OAI21_X1 U86378 ( .B1(n106134), .B2(n81451), .A(n97767), .ZN(
        \DLX_Datapath/RegisterFile/N23607 ) );
  AOI22_X1 U86379 ( .A1(n81506), .A2(n106126), .B1(n106124), .B2(n107683), 
        .ZN(n97767) );
  OAI21_X1 U86380 ( .B1(n106199), .B2(n106133), .A(n97768), .ZN(
        \DLX_Datapath/RegisterFile/N23606 ) );
  AOI22_X1 U86381 ( .A1(n81385), .A2(n81313), .B1(n106124), .B2(n109601), .ZN(
        n97768) );
  OAI21_X1 U86382 ( .B1(n106246), .B2(n106133), .A(n97769), .ZN(
        \DLX_Datapath/RegisterFile/N23605 ) );
  AOI22_X1 U86383 ( .A1(n106126), .A2(n81330), .B1(n106124), .B2(n108562), 
        .ZN(n97769) );
  OAI21_X1 U86384 ( .B1(n106159), .B2(n106133), .A(n97770), .ZN(
        \DLX_Datapath/RegisterFile/N23604 ) );
  AOI22_X1 U86385 ( .A1(n81425), .A2(n81385), .B1(n106124), .B2(n109706), .ZN(
        n97770) );
  OAI21_X1 U86386 ( .B1(n106134), .B2(n106116), .A(n97771), .ZN(
        \DLX_Datapath/RegisterFile/N23603 ) );
  AOI22_X1 U86387 ( .A1(n81396), .A2(n106126), .B1(n106125), .B2(n109490), 
        .ZN(n97771) );
  OAI21_X1 U86388 ( .B1(n106010), .B2(n106133), .A(n97772), .ZN(
        \DLX_Datapath/RegisterFile/N23602 ) );
  AOI22_X1 U86389 ( .A1(n81590), .A2(n106127), .B1(n106125), .B2(n109027), 
        .ZN(n97772) );
  OAI21_X1 U86390 ( .B1(n106261), .B2(n106133), .A(n97773), .ZN(
        \DLX_Datapath/RegisterFile/N23601 ) );
  AOI22_X1 U86391 ( .A1(n81423), .A2(n106126), .B1(n106125), .B2(n109375), 
        .ZN(n97773) );
  OAI21_X1 U86392 ( .B1(n106133), .B2(n81509), .A(n97774), .ZN(
        \DLX_Datapath/RegisterFile/N23600 ) );
  AOI22_X1 U86393 ( .A1(n81511), .A2(n106126), .B1(n106125), .B2(n109257), 
        .ZN(n97774) );
  OAI21_X1 U86394 ( .B1(n106134), .B2(n81501), .A(n97775), .ZN(
        \DLX_Datapath/RegisterFile/N23599 ) );
  AOI22_X1 U86395 ( .A1(n81503), .A2(n106127), .B1(n106125), .B2(n109148), 
        .ZN(n97775) );
  OAI21_X1 U86396 ( .B1(n106133), .B2(n81415), .A(n97776), .ZN(
        \DLX_Datapath/RegisterFile/N23598 ) );
  AOI22_X1 U86397 ( .A1(n81417), .A2(n106126), .B1(n106125), .B2(n108684), 
        .ZN(n97776) );
  OAI21_X1 U86398 ( .B1(n106133), .B2(n81498), .A(n97777), .ZN(
        \DLX_Datapath/RegisterFile/N23597 ) );
  AOI22_X1 U86399 ( .A1(n81500), .A2(n106127), .B1(n106125), .B2(n108911), 
        .ZN(n97777) );
  OAI21_X1 U86400 ( .B1(n105217), .B2(n106134), .A(n97778), .ZN(
        \DLX_Datapath/RegisterFile/N23596 ) );
  AOI22_X1 U86401 ( .A1(n81385), .A2(n81335), .B1(n106125), .B2(n108799), .ZN(
        n97778) );
  OAI21_X1 U86402 ( .B1(n106269), .B2(n106134), .A(n97779), .ZN(
        \DLX_Datapath/RegisterFile/N23595 ) );
  AOI22_X1 U86403 ( .A1(n81385), .A2(n81327), .B1(n106124), .B2(n107339), .ZN(
        n97779) );
  NOR2_X1 U86404 ( .A1(n97748), .A2(n97780), .ZN(n81387) );
  NOR2_X1 U86405 ( .A1(n97710), .A2(n97780), .ZN(n81385) );
  NOR2_X1 U86406 ( .A1(n81382), .A2(n105094), .ZN(n97780) );
  NAND2_X1 U86407 ( .A1(n105126), .A2(n95132), .ZN(n81382) );
  OAI21_X1 U86408 ( .B1(n106148), .B2(n105313), .A(n97782), .ZN(
        \DLX_Datapath/RegisterFile/N23594 ) );
  AOI22_X1 U86409 ( .A1(n105311), .A2(n94667), .B1(n105309), .B2(n107900), 
        .ZN(n97782) );
  OAI21_X1 U86410 ( .B1(n105969), .B2(n105313), .A(n97785), .ZN(
        \DLX_Datapath/RegisterFile/N23593 ) );
  AOI22_X1 U86411 ( .A1(n97783), .A2(n94670), .B1(n97784), .B2(n107994), .ZN(
        n97785) );
  OAI21_X1 U86412 ( .B1(n106137), .B2(n105313), .A(n97786), .ZN(
        \DLX_Datapath/RegisterFile/N23592 ) );
  AOI22_X1 U86413 ( .A1(n105311), .A2(n94672), .B1(n105309), .B2(n107264), 
        .ZN(n97786) );
  OAI21_X1 U86414 ( .B1(n106210), .B2(n105313), .A(n97787), .ZN(
        \DLX_Datapath/RegisterFile/N23591 ) );
  AOI22_X1 U86415 ( .A1(n97783), .A2(n94674), .B1(n97784), .B2(n107801), .ZN(
        n97787) );
  OAI21_X1 U86416 ( .B1(n106205), .B2(n105313), .A(n97788), .ZN(
        \DLX_Datapath/RegisterFile/N23590 ) );
  AOI22_X1 U86417 ( .A1(n105311), .A2(n94676), .B1(n105309), .B2(n110700), 
        .ZN(n97788) );
  OAI21_X1 U86418 ( .B1(n106100), .B2(n105313), .A(n97789), .ZN(
        \DLX_Datapath/RegisterFile/N23589 ) );
  AOI22_X1 U86419 ( .A1(n97783), .A2(n94678), .B1(n97784), .B2(n108103), .ZN(
        n97789) );
  OAI21_X1 U86420 ( .B1(n106256), .B2(n105313), .A(n97790), .ZN(
        \DLX_Datapath/RegisterFile/N23588 ) );
  AOI22_X1 U86421 ( .A1(n105311), .A2(n94680), .B1(n105309), .B2(n110802), 
        .ZN(n97790) );
  OAI21_X1 U86422 ( .B1(n105991), .B2(n105313), .A(n97791), .ZN(
        \DLX_Datapath/RegisterFile/N23587 ) );
  AOI22_X1 U86423 ( .A1(n105310), .A2(n94682), .B1(n105308), .B2(n110899), 
        .ZN(n97791) );
  OAI21_X1 U86424 ( .B1(n106331), .B2(n105313), .A(n97792), .ZN(
        \DLX_Datapath/RegisterFile/N23586 ) );
  AOI22_X1 U86425 ( .A1(n105310), .A2(n94684), .B1(n105308), .B2(n110494), 
        .ZN(n97792) );
  OAI21_X1 U86426 ( .B1(n106191), .B2(n105312), .A(n97793), .ZN(
        \DLX_Datapath/RegisterFile/N23585 ) );
  AOI22_X1 U86427 ( .A1(n105310), .A2(n94686), .B1(n105308), .B2(n110277), 
        .ZN(n97793) );
  OAI21_X1 U86428 ( .B1(n106130), .B2(n105312), .A(n97794), .ZN(
        \DLX_Datapath/RegisterFile/N23584 ) );
  AOI22_X1 U86429 ( .A1(n105310), .A2(n94688), .B1(n105308), .B2(n110596), 
        .ZN(n97794) );
  OAI21_X1 U86430 ( .B1(n106187), .B2(n105312), .A(n97795), .ZN(
        \DLX_Datapath/RegisterFile/N23583 ) );
  AOI22_X1 U86431 ( .A1(n105310), .A2(n94690), .B1(n105308), .B2(n110386), 
        .ZN(n97795) );
  OAI21_X1 U86432 ( .B1(n106164), .B2(n105312), .A(n97796), .ZN(
        \DLX_Datapath/RegisterFile/N23582 ) );
  AOI22_X1 U86433 ( .A1(n105310), .A2(n94692), .B1(n105308), .B2(n110064), 
        .ZN(n97796) );
  OAI21_X1 U86434 ( .B1(n106105), .B2(n105312), .A(n97797), .ZN(
        \DLX_Datapath/RegisterFile/N23581 ) );
  AOI22_X1 U86435 ( .A1(n105310), .A2(n94694), .B1(n105308), .B2(n110171), 
        .ZN(n97797) );
  OAI21_X1 U86436 ( .B1(n106220), .B2(n105312), .A(n97798), .ZN(
        \DLX_Datapath/RegisterFile/N23580 ) );
  AOI22_X1 U86437 ( .A1(n105310), .A2(n94696), .B1(n105308), .B2(n109955), 
        .ZN(n97798) );
  OAI21_X1 U86438 ( .B1(n106110), .B2(n105312), .A(n97799), .ZN(
        \DLX_Datapath/RegisterFile/N23579 ) );
  AOI22_X1 U86439 ( .A1(n105310), .A2(n94698), .B1(n105308), .B2(n109838), 
        .ZN(n97799) );
  OAI21_X1 U86440 ( .B1(n106232), .B2(n105312), .A(n97800), .ZN(
        \DLX_Datapath/RegisterFile/N23578 ) );
  AOI22_X1 U86441 ( .A1(n105310), .A2(n94700), .B1(n105308), .B2(n108212), 
        .ZN(n97800) );
  OAI21_X1 U86442 ( .B1(n106173), .B2(n105312), .A(n97801), .ZN(
        \DLX_Datapath/RegisterFile/N23577 ) );
  AOI22_X1 U86443 ( .A1(n105310), .A2(n94702), .B1(n105308), .B2(n108335), 
        .ZN(n97801) );
  OAI21_X1 U86444 ( .B1(n106237), .B2(n105312), .A(n97802), .ZN(
        \DLX_Datapath/RegisterFile/N23576 ) );
  AOI22_X1 U86445 ( .A1(n105310), .A2(n94704), .B1(n105308), .B2(n108446), 
        .ZN(n97802) );
  OAI21_X1 U86446 ( .B1(n106069), .B2(n105312), .A(n97803), .ZN(
        \DLX_Datapath/RegisterFile/N23575 ) );
  AOI22_X1 U86447 ( .A1(n105310), .A2(n94706), .B1(n105308), .B2(n107684), 
        .ZN(n97803) );
  OAI21_X1 U86448 ( .B1(n106199), .B2(n105312), .A(n97804), .ZN(
        \DLX_Datapath/RegisterFile/N23574 ) );
  AOI22_X1 U86449 ( .A1(n97783), .A2(n94708), .B1(n97784), .B2(n109602), .ZN(
        n97804) );
  OAI21_X1 U86450 ( .B1(n106246), .B2(n105313), .A(n97805), .ZN(
        \DLX_Datapath/RegisterFile/N23573 ) );
  AOI22_X1 U86451 ( .A1(n105311), .A2(n94710), .B1(n105309), .B2(n108563), 
        .ZN(n97805) );
  OAI21_X1 U86452 ( .B1(n106160), .B2(n105313), .A(n97806), .ZN(
        \DLX_Datapath/RegisterFile/N23572 ) );
  AOI22_X1 U86453 ( .A1(n97783), .A2(n94712), .B1(n97784), .B2(n109707), .ZN(
        n97806) );
  OAI21_X1 U86454 ( .B1(n106115), .B2(n105312), .A(n97807), .ZN(
        \DLX_Datapath/RegisterFile/N23571 ) );
  AOI22_X1 U86455 ( .A1(n105311), .A2(n94714), .B1(n105309), .B2(n109491), 
        .ZN(n97807) );
  OAI21_X1 U86456 ( .B1(n106010), .B2(n105313), .A(n97808), .ZN(
        \DLX_Datapath/RegisterFile/N23570 ) );
  AOI22_X1 U86457 ( .A1(n97783), .A2(n81259), .B1(n97784), .B2(n109028), .ZN(
        n97808) );
  OAI21_X1 U86458 ( .B1(n106261), .B2(n105313), .A(n97809), .ZN(
        \DLX_Datapath/RegisterFile/N23569 ) );
  AOI22_X1 U86459 ( .A1(n105311), .A2(n94717), .B1(n105309), .B2(n109376), 
        .ZN(n97809) );
  OAI21_X1 U86460 ( .B1(n106044), .B2(n105312), .A(n97810), .ZN(
        \DLX_Datapath/RegisterFile/N23568 ) );
  AOI22_X1 U86461 ( .A1(n97783), .A2(n94719), .B1(n97784), .B2(n109258), .ZN(
        n97810) );
  OAI21_X1 U86462 ( .B1(n106048), .B2(n105313), .A(n97811), .ZN(
        \DLX_Datapath/RegisterFile/N23567 ) );
  AOI22_X1 U86463 ( .A1(n105311), .A2(n94721), .B1(n105309), .B2(n109149), 
        .ZN(n97811) );
  OAI21_X1 U86464 ( .B1(n106095), .B2(n105312), .A(n97812), .ZN(
        \DLX_Datapath/RegisterFile/N23566 ) );
  AOI22_X1 U86465 ( .A1(n97783), .A2(n94723), .B1(n97784), .B2(n108685), .ZN(
        n97812) );
  OAI21_X1 U86466 ( .B1(n106056), .B2(n105313), .A(n97813), .ZN(
        \DLX_Datapath/RegisterFile/N23565 ) );
  AOI22_X1 U86467 ( .A1(n105311), .A2(n94725), .B1(n105309), .B2(n108912), 
        .ZN(n97813) );
  OAI21_X1 U86468 ( .B1(n105217), .B2(n105313), .A(n97814), .ZN(
        \DLX_Datapath/RegisterFile/N23564 ) );
  AOI22_X1 U86469 ( .A1(n105311), .A2(n94727), .B1(n105309), .B2(n108800), 
        .ZN(n97814) );
  OAI21_X1 U86470 ( .B1(n106269), .B2(n105312), .A(n97815), .ZN(
        \DLX_Datapath/RegisterFile/N23563 ) );
  AOI22_X1 U86471 ( .A1(n105311), .A2(n94729), .B1(n105309), .B2(n107340), 
        .ZN(n97815) );
  NOR2_X1 U86472 ( .A1(n97748), .A2(n97816), .ZN(n97784) );
  AOI21_X1 U86473 ( .B1(n105205), .B2(n97710), .A(n94663), .ZN(n97748) );
  NOR2_X1 U86474 ( .A1(n97710), .A2(n97816), .ZN(n97783) );
  NOR2_X1 U86475 ( .A1(n97781), .A2(n105093), .ZN(n97816) );
  OR2_X1 U86476 ( .A1(n97674), .A2(n95131), .ZN(n97710) );
  NAND2_X1 U86477 ( .A1(n105125), .A2(n94505), .ZN(n97781) );
  OAI21_X1 U86478 ( .B1(n106155), .B2(n105971), .A(n97817), .ZN(
        \DLX_Datapath/RegisterFile/N23561 ) );
  AOI22_X1 U86479 ( .A1(n106153), .A2(n107995), .B1(n94511), .B2(n106151), 
        .ZN(n97817) );
  OAI21_X1 U86480 ( .B1(n106156), .B2(n106137), .A(n97818), .ZN(
        \DLX_Datapath/RegisterFile/N23560 ) );
  AOI22_X1 U86481 ( .A1(n81355), .A2(n107265), .B1(n81539), .B2(n106152), .ZN(
        n97818) );
  OAI21_X1 U86482 ( .B1(n106205), .B2(n106155), .A(n97819), .ZN(
        \DLX_Datapath/RegisterFile/N23558 ) );
  AOI22_X1 U86483 ( .A1(n74065), .A2(n106154), .B1(n106151), .B2(n81308), .ZN(
        n97819) );
  OAI21_X1 U86484 ( .B1(n106156), .B2(n106098), .A(n97820), .ZN(
        \DLX_Datapath/RegisterFile/N23557 ) );
  AOI22_X1 U86485 ( .A1(n70652), .A2(n106154), .B1(n94516), .B2(n106152), .ZN(
        n97820) );
  OAI21_X1 U86486 ( .B1(n106256), .B2(n106155), .A(n97821), .ZN(
        \DLX_Datapath/RegisterFile/N23556 ) );
  AOI22_X1 U86487 ( .A1(n74206), .A2(n106154), .B1(n106151), .B2(n81272), .ZN(
        n97821) );
  OAI21_X1 U86488 ( .B1(n106156), .B2(n81629), .A(n97822), .ZN(
        \DLX_Datapath/RegisterFile/N23555 ) );
  AOI22_X1 U86489 ( .A1(n106153), .A2(n111037), .B1(n94519), .B2(n106152), 
        .ZN(n97822) );
  OAI21_X1 U86490 ( .B1(n106331), .B2(n106155), .A(n97823), .ZN(
        \DLX_Datapath/RegisterFile/N23554 ) );
  AOI22_X1 U86491 ( .A1(n106153), .A2(n111036), .B1(n106151), .B2(n80192), 
        .ZN(n97823) );
  OAI21_X1 U86492 ( .B1(n106192), .B2(n106155), .A(n97824), .ZN(
        \DLX_Datapath/RegisterFile/N23553 ) );
  AOI22_X1 U86493 ( .A1(n106153), .A2(n110278), .B1(n81474), .B2(n81356), .ZN(
        n97824) );
  OAI21_X1 U86494 ( .B1(n106155), .B2(n106128), .A(n97825), .ZN(
        \DLX_Datapath/RegisterFile/N23552 ) );
  AOI22_X1 U86495 ( .A1(n106153), .A2(n110597), .B1(n94523), .B2(n81356), .ZN(
        n97825) );
  OAI21_X1 U86496 ( .B1(n106187), .B2(n106155), .A(n97826), .ZN(
        \DLX_Datapath/RegisterFile/N23551 ) );
  AOI22_X1 U86497 ( .A1(n106153), .A2(n110387), .B1(n106062), .B2(n81356), 
        .ZN(n97826) );
  OAI21_X1 U86498 ( .B1(n106164), .B2(n106155), .A(n97827), .ZN(
        \DLX_Datapath/RegisterFile/N23550 ) );
  AOI22_X1 U86499 ( .A1(n106153), .A2(n110065), .B1(n106151), .B2(n81347), 
        .ZN(n97827) );
  OAI21_X1 U86500 ( .B1(n106156), .B2(n81403), .A(n97828), .ZN(
        \DLX_Datapath/RegisterFile/N23549 ) );
  AOI22_X1 U86501 ( .A1(n106153), .A2(n110172), .B1(n94527), .B2(n106152), 
        .ZN(n97828) );
  OAI21_X1 U86502 ( .B1(n106220), .B2(n106155), .A(n97829), .ZN(
        \DLX_Datapath/RegisterFile/N23548 ) );
  AOI22_X1 U86503 ( .A1(n106153), .A2(n109956), .B1(n106151), .B2(n81297), 
        .ZN(n97829) );
  OAI21_X1 U86504 ( .B1(n106156), .B2(n81398), .A(n97830), .ZN(
        \DLX_Datapath/RegisterFile/N23547 ) );
  AOI22_X1 U86505 ( .A1(n106153), .A2(n109839), .B1(n94530), .B2(n106152), 
        .ZN(n97830) );
  OAI21_X1 U86506 ( .B1(n106156), .B2(n106069), .A(n97831), .ZN(
        \DLX_Datapath/RegisterFile/N23543 ) );
  AOI22_X1 U86507 ( .A1(n106154), .A2(n107685), .B1(n81453), .B2(n81356), .ZN(
        n97831) );
  OAI21_X1 U86508 ( .B1(n106199), .B2(n106155), .A(n97832), .ZN(
        \DLX_Datapath/RegisterFile/N23542 ) );
  AOI22_X1 U86509 ( .A1(n106154), .A2(n109603), .B1(n94536), .B2(n81356), .ZN(
        n97832) );
  OAI21_X1 U86510 ( .B1(n106155), .B2(n106113), .A(n97833), .ZN(
        \DLX_Datapath/RegisterFile/N23539 ) );
  AOI22_X1 U86511 ( .A1(n106154), .A2(n109492), .B1(n106021), .B2(n106151), 
        .ZN(n97833) );
  OAI21_X1 U86512 ( .B1(n106010), .B2(n106155), .A(n97834), .ZN(
        \DLX_Datapath/RegisterFile/N23538 ) );
  AOI22_X1 U86513 ( .A1(n106154), .A2(n109029), .B1(n94541), .B2(n106151), 
        .ZN(n97834) );
  OAI21_X1 U86514 ( .B1(n106156), .B2(n81509), .A(n97835), .ZN(
        \DLX_Datapath/RegisterFile/N23536 ) );
  AOI22_X1 U86515 ( .A1(n106154), .A2(n109259), .B1(n105625), .B2(n106151), 
        .ZN(n97835) );
  OAI21_X1 U86516 ( .B1(n106155), .B2(n81501), .A(n97836), .ZN(
        \DLX_Datapath/RegisterFile/N23535 ) );
  AOI22_X1 U86517 ( .A1(n106154), .A2(n109150), .B1(n94546), .B2(n106151), 
        .ZN(n97836) );
  OAI21_X1 U86518 ( .B1(n106155), .B2(n106095), .A(n97837), .ZN(
        \DLX_Datapath/RegisterFile/N23534 ) );
  AOI22_X1 U86519 ( .A1(n106154), .A2(n108686), .B1(n94548), .B2(n106151), 
        .ZN(n97837) );
  OAI21_X1 U86520 ( .B1(n106155), .B2(n81498), .A(n97838), .ZN(
        \DLX_Datapath/RegisterFile/N23533 ) );
  AOI22_X1 U86521 ( .A1(n106154), .A2(n108913), .B1(n81783), .B2(n106151), 
        .ZN(n97838) );
  OAI21_X1 U86522 ( .B1(n106269), .B2(n106156), .A(n97839), .ZN(
        \DLX_Datapath/RegisterFile/N23531 ) );
  AOI22_X1 U86523 ( .A1(n81355), .A2(n107341), .B1(n106152), .B2(n81265), .ZN(
        n97839) );
  NOR2_X1 U86524 ( .A1(n97840), .A2(n97841), .ZN(n81356) );
  AOI21_X1 U86525 ( .B1(n97572), .B2(n94554), .A(n97841), .ZN(n81355) );
  NOR2_X1 U86526 ( .A1(n81353), .A2(n105091), .ZN(n97841) );
  NAND2_X1 U86527 ( .A1(n105126), .A2(n94555), .ZN(n81353) );
  OAI21_X1 U86528 ( .B1(n106148), .B2(n105307), .A(n97843), .ZN(
        \DLX_Datapath/RegisterFile/N23530 ) );
  AOI22_X1 U86529 ( .A1(n105305), .A2(n70364), .B1(n105303), .B2(n94559), .ZN(
        n97843) );
  OAI21_X1 U86530 ( .B1(n105969), .B2(n105307), .A(n97846), .ZN(
        \DLX_Datapath/RegisterFile/N23529 ) );
  AOI22_X1 U86531 ( .A1(n97844), .A2(n70506), .B1(n105302), .B2(n94562), .ZN(
        n97846) );
  OAI21_X1 U86532 ( .B1(n106137), .B2(n105307), .A(n97847), .ZN(
        \DLX_Datapath/RegisterFile/N23528 ) );
  AOI22_X1 U86533 ( .A1(n105305), .A2(n107266), .B1(n105303), .B2(n94564), 
        .ZN(n97847) );
  OAI21_X1 U86534 ( .B1(n106210), .B2(n105307), .A(n97848), .ZN(
        \DLX_Datapath/RegisterFile/N23527 ) );
  AOI22_X1 U86535 ( .A1(n97844), .A2(n107803), .B1(n105302), .B2(n94566), .ZN(
        n97848) );
  OAI21_X1 U86536 ( .B1(n106205), .B2(n105307), .A(n97849), .ZN(
        \DLX_Datapath/RegisterFile/N23526 ) );
  AOI22_X1 U86537 ( .A1(n105305), .A2(n110701), .B1(n105303), .B2(n94568), 
        .ZN(n97849) );
  OAI21_X1 U86538 ( .B1(n106100), .B2(n105307), .A(n97850), .ZN(
        \DLX_Datapath/RegisterFile/N23525 ) );
  AOI22_X1 U86539 ( .A1(n97844), .A2(n108104), .B1(n105302), .B2(n94570), .ZN(
        n97850) );
  OAI21_X1 U86540 ( .B1(n106256), .B2(n105307), .A(n97851), .ZN(
        \DLX_Datapath/RegisterFile/N23524 ) );
  AOI22_X1 U86541 ( .A1(n105305), .A2(n110803), .B1(n105303), .B2(n94572), 
        .ZN(n97851) );
  OAI21_X1 U86542 ( .B1(n81629), .B2(n105307), .A(n97852), .ZN(
        \DLX_Datapath/RegisterFile/N23523 ) );
  AOI22_X1 U86543 ( .A1(n105304), .A2(n110900), .B1(n105302), .B2(n94574), 
        .ZN(n97852) );
  OAI21_X1 U86544 ( .B1(n106331), .B2(n105307), .A(n97853), .ZN(
        \DLX_Datapath/RegisterFile/N23522 ) );
  AOI22_X1 U86545 ( .A1(n97844), .A2(n110495), .B1(n105302), .B2(n94576), .ZN(
        n97853) );
  OAI21_X1 U86546 ( .B1(n106192), .B2(n105306), .A(n97854), .ZN(
        \DLX_Datapath/RegisterFile/N23521 ) );
  AOI22_X1 U86547 ( .A1(n105304), .A2(n110279), .B1(n97845), .B2(n94578), .ZN(
        n97854) );
  OAI21_X1 U86548 ( .B1(n106131), .B2(n105306), .A(n97855), .ZN(
        \DLX_Datapath/RegisterFile/N23520 ) );
  AOI22_X1 U86549 ( .A1(n105304), .A2(n110598), .B1(n97845), .B2(n94580), .ZN(
        n97855) );
  OAI21_X1 U86550 ( .B1(n106187), .B2(n105306), .A(n97856), .ZN(
        \DLX_Datapath/RegisterFile/N23519 ) );
  AOI22_X1 U86551 ( .A1(n105304), .A2(n110388), .B1(n97845), .B2(n94582), .ZN(
        n97856) );
  OAI21_X1 U86552 ( .B1(n106165), .B2(n105306), .A(n97857), .ZN(
        \DLX_Datapath/RegisterFile/N23518 ) );
  AOI22_X1 U86553 ( .A1(n105304), .A2(n110066), .B1(n105303), .B2(n94584), 
        .ZN(n97857) );
  OAI21_X1 U86554 ( .B1(n106106), .B2(n105306), .A(n97858), .ZN(
        \DLX_Datapath/RegisterFile/N23517 ) );
  AOI22_X1 U86555 ( .A1(n105304), .A2(n110173), .B1(n97845), .B2(n94586), .ZN(
        n97858) );
  OAI21_X1 U86556 ( .B1(n106220), .B2(n105306), .A(n97859), .ZN(
        \DLX_Datapath/RegisterFile/N23516 ) );
  AOI22_X1 U86557 ( .A1(n105304), .A2(n109957), .B1(n97845), .B2(n94588), .ZN(
        n97859) );
  OAI21_X1 U86558 ( .B1(n106110), .B2(n105306), .A(n97860), .ZN(
        \DLX_Datapath/RegisterFile/N23515 ) );
  AOI22_X1 U86559 ( .A1(n105304), .A2(n109840), .B1(n97845), .B2(n94590), .ZN(
        n97860) );
  OAI21_X1 U86560 ( .B1(n106232), .B2(n105306), .A(n97861), .ZN(
        \DLX_Datapath/RegisterFile/N23514 ) );
  AOI22_X1 U86561 ( .A1(n105304), .A2(n108214), .B1(n97845), .B2(n94592), .ZN(
        n97861) );
  OAI21_X1 U86562 ( .B1(n106173), .B2(n105306), .A(n97862), .ZN(
        \DLX_Datapath/RegisterFile/N23513 ) );
  AOI22_X1 U86563 ( .A1(n105304), .A2(n108337), .B1(n105302), .B2(n94594), 
        .ZN(n97862) );
  OAI21_X1 U86564 ( .B1(n106237), .B2(n105306), .A(n97863), .ZN(
        \DLX_Datapath/RegisterFile/N23512 ) );
  AOI22_X1 U86565 ( .A1(n105304), .A2(n108448), .B1(n105302), .B2(n94596), 
        .ZN(n97863) );
  OAI21_X1 U86566 ( .B1(n106069), .B2(n105306), .A(n97864), .ZN(
        \DLX_Datapath/RegisterFile/N23511 ) );
  AOI22_X1 U86567 ( .A1(n105304), .A2(n107686), .B1(n97845), .B2(n94598), .ZN(
        n97864) );
  OAI21_X1 U86568 ( .B1(n106199), .B2(n105306), .A(n97865), .ZN(
        \DLX_Datapath/RegisterFile/N23510 ) );
  AOI22_X1 U86569 ( .A1(n97844), .A2(n109604), .B1(n105302), .B2(n94600), .ZN(
        n97865) );
  OAI21_X1 U86570 ( .B1(n106246), .B2(n105307), .A(n97866), .ZN(
        \DLX_Datapath/RegisterFile/N23509 ) );
  AOI22_X1 U86571 ( .A1(n105305), .A2(n108565), .B1(n105303), .B2(n94602), 
        .ZN(n97866) );
  OAI21_X1 U86572 ( .B1(n106160), .B2(n105307), .A(n97867), .ZN(
        \DLX_Datapath/RegisterFile/N23508 ) );
  AOI22_X1 U86573 ( .A1(n97844), .A2(n109709), .B1(n105302), .B2(n94604), .ZN(
        n97867) );
  OAI21_X1 U86574 ( .B1(n106115), .B2(n105306), .A(n97868), .ZN(
        \DLX_Datapath/RegisterFile/N23507 ) );
  AOI22_X1 U86575 ( .A1(n105305), .A2(n109493), .B1(n105303), .B2(n94606), 
        .ZN(n97868) );
  OAI21_X1 U86576 ( .B1(n106011), .B2(n105307), .A(n97869), .ZN(
        \DLX_Datapath/RegisterFile/N23506 ) );
  AOI22_X1 U86577 ( .A1(n97844), .A2(n109030), .B1(n105302), .B2(n94608), .ZN(
        n97869) );
  OAI21_X1 U86578 ( .B1(n106261), .B2(n105307), .A(n97870), .ZN(
        \DLX_Datapath/RegisterFile/N23505 ) );
  AOI22_X1 U86579 ( .A1(n105305), .A2(n109378), .B1(n105303), .B2(n94610), 
        .ZN(n97870) );
  OAI21_X1 U86580 ( .B1(n106045), .B2(n105306), .A(n97871), .ZN(
        \DLX_Datapath/RegisterFile/N23504 ) );
  AOI22_X1 U86581 ( .A1(n105304), .A2(n109260), .B1(n105302), .B2(n94612), 
        .ZN(n97871) );
  OAI21_X1 U86582 ( .B1(n106050), .B2(n105307), .A(n97872), .ZN(
        \DLX_Datapath/RegisterFile/N23503 ) );
  AOI22_X1 U86583 ( .A1(n105305), .A2(n109151), .B1(n105303), .B2(n94614), 
        .ZN(n97872) );
  OAI21_X1 U86584 ( .B1(n106096), .B2(n105306), .A(n97873), .ZN(
        \DLX_Datapath/RegisterFile/N23502 ) );
  AOI22_X1 U86585 ( .A1(n97844), .A2(n108687), .B1(n105302), .B2(n94616), .ZN(
        n97873) );
  OAI21_X1 U86586 ( .B1(n106055), .B2(n105307), .A(n97874), .ZN(
        \DLX_Datapath/RegisterFile/N23501 ) );
  AOI22_X1 U86587 ( .A1(n105305), .A2(n108914), .B1(n105303), .B2(n94618), 
        .ZN(n97874) );
  OAI21_X1 U86588 ( .B1(n105216), .B2(n105307), .A(n97875), .ZN(
        \DLX_Datapath/RegisterFile/N23500 ) );
  AOI22_X1 U86589 ( .A1(n105305), .A2(n108802), .B1(n105303), .B2(n94620), 
        .ZN(n97875) );
  OAI21_X1 U86590 ( .B1(n106269), .B2(n105306), .A(n97876), .ZN(
        \DLX_Datapath/RegisterFile/N23499 ) );
  AOI22_X1 U86591 ( .A1(n105305), .A2(n107342), .B1(n105302), .B2(n94622), 
        .ZN(n97876) );
  NOR2_X1 U86592 ( .A1(n97840), .A2(n97877), .ZN(n97845) );
  NOR2_X1 U86593 ( .A1(n97877), .A2(n97878), .ZN(n97844) );
  NOR2_X1 U86594 ( .A1(n97842), .A2(n105093), .ZN(n97877) );
  NAND2_X1 U86595 ( .A1(n94625), .A2(n105125), .ZN(n97842) );
  OAI21_X1 U86596 ( .B1(n106149), .B2(n106123), .A(n97879), .ZN(
        \DLX_Datapath/RegisterFile/N23498 ) );
  AOI22_X1 U86597 ( .A1(n70365), .A2(n106120), .B1(n81521), .B2(n106119), .ZN(
        n97879) );
  OAI21_X1 U86598 ( .B1(n106123), .B2(n81651), .A(n97880), .ZN(
        \DLX_Datapath/RegisterFile/N23497 ) );
  AOI22_X1 U86599 ( .A1(n70507), .A2(n106120), .B1(n81653), .B2(n81391), .ZN(
        n97880) );
  OAI21_X1 U86600 ( .B1(n106138), .B2(n106123), .A(n97881), .ZN(
        \DLX_Datapath/RegisterFile/N23496 ) );
  AOI22_X1 U86601 ( .A1(n69560), .A2(n106120), .B1(n106119), .B2(n81380), .ZN(
        n97881) );
  OAI21_X1 U86602 ( .B1(n106205), .B2(n106123), .A(n97882), .ZN(
        \DLX_Datapath/RegisterFile/N23494 ) );
  AOI22_X1 U86603 ( .A1(n74067), .A2(n106120), .B1(n81428), .B2(n81391), .ZN(
        n97882) );
  OAI21_X1 U86604 ( .B1(n106256), .B2(n106123), .A(n97883), .ZN(
        \DLX_Datapath/RegisterFile/N23492 ) );
  AOI22_X1 U86605 ( .A1(n74208), .A2(n106121), .B1(n81700), .B2(n81391), .ZN(
        n97883) );
  OAI21_X1 U86606 ( .B1(n106122), .B2(n81629), .A(n97884), .ZN(
        \DLX_Datapath/RegisterFile/N23491 ) );
  AOI22_X1 U86607 ( .A1(n74348), .A2(n106121), .B1(n81632), .B2(n106119), .ZN(
        n97884) );
  OAI21_X1 U86608 ( .B1(n106192), .B2(n106123), .A(n97885), .ZN(
        \DLX_Datapath/RegisterFile/N23489 ) );
  AOI22_X1 U86609 ( .A1(n73488), .A2(n81390), .B1(n106118), .B2(n81317), .ZN(
        n97885) );
  OAI21_X1 U86610 ( .B1(n106165), .B2(n106123), .A(n97886), .ZN(
        \DLX_Datapath/RegisterFile/N23486 ) );
  AOI22_X1 U86611 ( .A1(n73199), .A2(n81390), .B1(n81604), .B2(n81391), .ZN(
        n97886) );
  OAI21_X1 U86612 ( .B1(n106123), .B2(n106071), .A(n97887), .ZN(
        \DLX_Datapath/RegisterFile/N23479 ) );
  AOI22_X1 U86613 ( .A1(n70068), .A2(n81390), .B1(n81506), .B2(n81391), .ZN(
        n97887) );
  OAI21_X1 U86614 ( .B1(n106160), .B2(n106123), .A(n97888), .ZN(
        \DLX_Datapath/RegisterFile/N23476 ) );
  AOI22_X1 U86615 ( .A1(n72739), .A2(n81390), .B1(n81425), .B2(n106118), .ZN(
        n97888) );
  OAI21_X1 U86616 ( .B1(n106011), .B2(n106123), .A(n97889), .ZN(
        \DLX_Datapath/RegisterFile/N23474 ) );
  AOI22_X1 U86617 ( .A1(n71849), .A2(n81390), .B1(n81590), .B2(n106119), .ZN(
        n97889) );
  OAI21_X1 U86618 ( .B1(n106261), .B2(n106123), .A(n97890), .ZN(
        \DLX_Datapath/RegisterFile/N23473 ) );
  AOI22_X1 U86619 ( .A1(n72298), .A2(n81390), .B1(n81423), .B2(n106118), .ZN(
        n97890) );
  OAI21_X1 U86620 ( .B1(n106123), .B2(n81509), .A(n97891), .ZN(
        \DLX_Datapath/RegisterFile/N23472 ) );
  AOI22_X1 U86621 ( .A1(n72147), .A2(n106121), .B1(n81511), .B2(n81391), .ZN(
        n97891) );
  OAI21_X1 U86622 ( .B1(n106123), .B2(n81501), .A(n97892), .ZN(
        \DLX_Datapath/RegisterFile/N23471 ) );
  AOI22_X1 U86623 ( .A1(n72003), .A2(n106121), .B1(n81503), .B2(n81391), .ZN(
        n97892) );
  OAI21_X1 U86624 ( .B1(n106123), .B2(n81498), .A(n97893), .ZN(
        \DLX_Datapath/RegisterFile/N23469 ) );
  AOI22_X1 U86625 ( .A1(n71700), .A2(n106121), .B1(n81500), .B2(n106118), .ZN(
        n97893) );
  OAI21_X1 U86626 ( .B1(n106269), .B2(n106122), .A(n97894), .ZN(
        \DLX_Datapath/RegisterFile/N23467 ) );
  AOI22_X1 U86627 ( .A1(n69665), .A2(n106120), .B1(n106119), .B2(n81327), .ZN(
        n97894) );
  NOR2_X1 U86628 ( .A1(n97840), .A2(n97895), .ZN(n81391) );
  NOR2_X1 U86629 ( .A1(n97878), .A2(n97895), .ZN(n81390) );
  NOR2_X1 U86630 ( .A1(n81388), .A2(n105095), .ZN(n97895) );
  NAND2_X1 U86631 ( .A1(n105125), .A2(n94664), .ZN(n81388) );
  OAI21_X1 U86632 ( .B1(n106149), .B2(n105301), .A(n97897), .ZN(
        \DLX_Datapath/RegisterFile/N23466 ) );
  AOI22_X1 U86633 ( .A1(n105299), .A2(n94667), .B1(n105297), .B2(n70366), .ZN(
        n97897) );
  OAI21_X1 U86634 ( .B1(n105969), .B2(n105301), .A(n97900), .ZN(
        \DLX_Datapath/RegisterFile/N23465 ) );
  AOI22_X1 U86635 ( .A1(n97898), .A2(n94670), .B1(n105297), .B2(n70508), .ZN(
        n97900) );
  OAI21_X1 U86636 ( .B1(n106138), .B2(n105301), .A(n97901), .ZN(
        \DLX_Datapath/RegisterFile/N23464 ) );
  AOI22_X1 U86637 ( .A1(n105299), .A2(n94672), .B1(n105297), .B2(n69561), .ZN(
        n97901) );
  OAI21_X1 U86638 ( .B1(n106210), .B2(n105301), .A(n97902), .ZN(
        \DLX_Datapath/RegisterFile/N23463 ) );
  AOI22_X1 U86639 ( .A1(n97898), .A2(n94674), .B1(n105297), .B2(n70222), .ZN(
        n97902) );
  OAI21_X1 U86640 ( .B1(n106205), .B2(n105301), .A(n97903), .ZN(
        \DLX_Datapath/RegisterFile/N23462 ) );
  AOI22_X1 U86641 ( .A1(n105299), .A2(n94676), .B1(n105297), .B2(n74068), .ZN(
        n97903) );
  OAI21_X1 U86642 ( .B1(n106100), .B2(n105301), .A(n97904), .ZN(
        \DLX_Datapath/RegisterFile/N23461 ) );
  AOI22_X1 U86643 ( .A1(n97898), .A2(n94678), .B1(n105297), .B2(n70655), .ZN(
        n97904) );
  OAI21_X1 U86644 ( .B1(n106256), .B2(n105301), .A(n97905), .ZN(
        \DLX_Datapath/RegisterFile/N23460 ) );
  AOI22_X1 U86645 ( .A1(n105299), .A2(n94680), .B1(n105297), .B2(n74209), .ZN(
        n97905) );
  OAI21_X1 U86646 ( .B1(n81629), .B2(n105301), .A(n97906), .ZN(
        \DLX_Datapath/RegisterFile/N23459 ) );
  AOI22_X1 U86647 ( .A1(n105298), .A2(n94682), .B1(n105297), .B2(n74349), .ZN(
        n97906) );
  OAI21_X1 U86648 ( .B1(n106331), .B2(n105301), .A(n97907), .ZN(
        \DLX_Datapath/RegisterFile/N23458 ) );
  AOI22_X1 U86649 ( .A1(n97898), .A2(n94684), .B1(n105297), .B2(n73785), .ZN(
        n97907) );
  OAI21_X1 U86650 ( .B1(n106192), .B2(n105300), .A(n97908), .ZN(
        \DLX_Datapath/RegisterFile/N23457 ) );
  AOI22_X1 U86651 ( .A1(n105298), .A2(n94686), .B1(n105297), .B2(n73489), .ZN(
        n97908) );
  OAI21_X1 U86652 ( .B1(n106131), .B2(n105300), .A(n97909), .ZN(
        \DLX_Datapath/RegisterFile/N23456 ) );
  AOI22_X1 U86653 ( .A1(n105298), .A2(n94688), .B1(n97899), .B2(n73926), .ZN(
        n97909) );
  OAI21_X1 U86654 ( .B1(n106187), .B2(n105300), .A(n97910), .ZN(
        \DLX_Datapath/RegisterFile/N23455 ) );
  AOI22_X1 U86655 ( .A1(n105298), .A2(n94690), .B1(n97899), .B2(n73638), .ZN(
        n97910) );
  OAI21_X1 U86656 ( .B1(n106165), .B2(n105300), .A(n97911), .ZN(
        \DLX_Datapath/RegisterFile/N23454 ) );
  AOI22_X1 U86657 ( .A1(n105298), .A2(n94692), .B1(n105297), .B2(n73200), .ZN(
        n97911) );
  OAI21_X1 U86658 ( .B1(n106106), .B2(n105300), .A(n97912), .ZN(
        \DLX_Datapath/RegisterFile/N23453 ) );
  AOI22_X1 U86659 ( .A1(n105298), .A2(n94694), .B1(n97899), .B2(n73342), .ZN(
        n97912) );
  OAI21_X1 U86660 ( .B1(n106220), .B2(n105300), .A(n97913), .ZN(
        \DLX_Datapath/RegisterFile/N23452 ) );
  AOI22_X1 U86661 ( .A1(n105298), .A2(n94696), .B1(n97899), .B2(n73058), .ZN(
        n97913) );
  OAI21_X1 U86662 ( .B1(n106110), .B2(n105300), .A(n97914), .ZN(
        \DLX_Datapath/RegisterFile/N23451 ) );
  AOI22_X1 U86663 ( .A1(n105298), .A2(n94698), .B1(n97899), .B2(n72908), .ZN(
        n97914) );
  OAI21_X1 U86664 ( .B1(n106232), .B2(n105300), .A(n97915), .ZN(
        \DLX_Datapath/RegisterFile/N23450 ) );
  AOI22_X1 U86665 ( .A1(n105298), .A2(n94700), .B1(n105296), .B2(n70804), .ZN(
        n97915) );
  OAI21_X1 U86666 ( .B1(n106173), .B2(n105300), .A(n97916), .ZN(
        \DLX_Datapath/RegisterFile/N23449 ) );
  AOI22_X1 U86667 ( .A1(n105298), .A2(n94702), .B1(n105297), .B2(n70963), .ZN(
        n97916) );
  OAI21_X1 U86668 ( .B1(n106237), .B2(n105300), .A(n97917), .ZN(
        \DLX_Datapath/RegisterFile/N23448 ) );
  AOI22_X1 U86669 ( .A1(n105298), .A2(n94704), .B1(n105297), .B2(n71108), .ZN(
        n97917) );
  OAI21_X1 U86670 ( .B1(n106069), .B2(n105300), .A(n97918), .ZN(
        \DLX_Datapath/RegisterFile/N23447 ) );
  AOI22_X1 U86671 ( .A1(n105298), .A2(n94706), .B1(n97899), .B2(n70069), .ZN(
        n97918) );
  OAI21_X1 U86672 ( .B1(n106199), .B2(n105300), .A(n97919), .ZN(
        \DLX_Datapath/RegisterFile/N23446 ) );
  AOI22_X1 U86673 ( .A1(n97898), .A2(n94708), .B1(n105296), .B2(n72598), .ZN(
        n97919) );
  OAI21_X1 U86674 ( .B1(n106246), .B2(n105301), .A(n97920), .ZN(
        \DLX_Datapath/RegisterFile/N23445 ) );
  AOI22_X1 U86675 ( .A1(n105299), .A2(n94710), .B1(n105296), .B2(n71257), .ZN(
        n97920) );
  OAI21_X1 U86676 ( .B1(n106160), .B2(n105301), .A(n97921), .ZN(
        \DLX_Datapath/RegisterFile/N23444 ) );
  AOI22_X1 U86677 ( .A1(n97898), .A2(n94712), .B1(n105296), .B2(n72740), .ZN(
        n97921) );
  OAI21_X1 U86678 ( .B1(n106115), .B2(n105300), .A(n97922), .ZN(
        \DLX_Datapath/RegisterFile/N23443 ) );
  AOI22_X1 U86679 ( .A1(n105299), .A2(n94714), .B1(n105296), .B2(n72450), .ZN(
        n97922) );
  OAI21_X1 U86680 ( .B1(n106011), .B2(n105301), .A(n97923), .ZN(
        \DLX_Datapath/RegisterFile/N23442 ) );
  AOI22_X1 U86681 ( .A1(n97898), .A2(n81259), .B1(n105296), .B2(n71850), .ZN(
        n97923) );
  OAI21_X1 U86682 ( .B1(n106261), .B2(n105301), .A(n97924), .ZN(
        \DLX_Datapath/RegisterFile/N23441 ) );
  AOI22_X1 U86683 ( .A1(n105299), .A2(n94717), .B1(n105296), .B2(n72299), .ZN(
        n97924) );
  OAI21_X1 U86684 ( .B1(n106045), .B2(n105300), .A(n97925), .ZN(
        \DLX_Datapath/RegisterFile/N23440 ) );
  AOI22_X1 U86685 ( .A1(n105298), .A2(n94719), .B1(n105296), .B2(n72148), .ZN(
        n97925) );
  OAI21_X1 U86686 ( .B1(n106050), .B2(n105301), .A(n97926), .ZN(
        \DLX_Datapath/RegisterFile/N23439 ) );
  AOI22_X1 U86687 ( .A1(n105299), .A2(n94721), .B1(n105296), .B2(n72004), .ZN(
        n97926) );
  OAI21_X1 U86688 ( .B1(n106096), .B2(n105300), .A(n97927), .ZN(
        \DLX_Datapath/RegisterFile/N23438 ) );
  AOI22_X1 U86689 ( .A1(n97898), .A2(n94723), .B1(n105296), .B2(n71406), .ZN(
        n97927) );
  OAI21_X1 U86690 ( .B1(n106055), .B2(n105301), .A(n97928), .ZN(
        \DLX_Datapath/RegisterFile/N23437 ) );
  AOI22_X1 U86691 ( .A1(n105299), .A2(n94725), .B1(n105296), .B2(n71701), .ZN(
        n97928) );
  OAI21_X1 U86692 ( .B1(n105216), .B2(n105301), .A(n97929), .ZN(
        \DLX_Datapath/RegisterFile/N23436 ) );
  AOI22_X1 U86693 ( .A1(n105299), .A2(n94727), .B1(n105296), .B2(n71557), .ZN(
        n97929) );
  OAI21_X1 U86694 ( .B1(n106269), .B2(n105300), .A(n97930), .ZN(
        \DLX_Datapath/RegisterFile/N23435 ) );
  AOI22_X1 U86695 ( .A1(n105299), .A2(n94729), .B1(n105296), .B2(n69666), .ZN(
        n97930) );
  NOR2_X1 U86696 ( .A1(n97878), .A2(n97931), .ZN(n97899) );
  AOI21_X1 U86697 ( .B1(n105199), .B2(n97840), .A(n105601), .ZN(n97878) );
  NOR2_X1 U86698 ( .A1(n97840), .A2(n97931), .ZN(n97898) );
  NOR2_X1 U86699 ( .A1(n97896), .A2(n105091), .ZN(n97931) );
  OR2_X1 U86700 ( .A1(n97674), .A2(n86230), .ZN(n97840) );
  NAND2_X1 U86701 ( .A1(n94734), .A2(n105126), .ZN(n97896) );
  OAI21_X1 U86702 ( .B1(n106149), .B2(n105295), .A(n97933), .ZN(
        \DLX_Datapath/RegisterFile/N23434 ) );
  AOI22_X1 U86703 ( .A1(n105292), .A2(n70367), .B1(n97935), .B2(n81360), .ZN(
        n97933) );
  OAI21_X1 U86704 ( .B1(n105968), .B2(n105295), .A(n97936), .ZN(
        \DLX_Datapath/RegisterFile/N23433 ) );
  AOI22_X1 U86705 ( .A1(n105293), .A2(n107996), .B1(n97935), .B2(n94511), .ZN(
        n97936) );
  OAI21_X1 U86706 ( .B1(n106138), .B2(n105295), .A(n97937), .ZN(
        \DLX_Datapath/RegisterFile/N23432 ) );
  AOI22_X1 U86707 ( .A1(n105293), .A2(n107267), .B1(n97935), .B2(n81539), .ZN(
        n97937) );
  OAI21_X1 U86708 ( .B1(n106210), .B2(n105295), .A(n97938), .ZN(
        \DLX_Datapath/RegisterFile/N23431 ) );
  AOI22_X1 U86709 ( .A1(n105292), .A2(n107804), .B1(n97935), .B2(n81301), .ZN(
        n97938) );
  OAI21_X1 U86710 ( .B1(n106205), .B2(n105295), .A(n97939), .ZN(
        \DLX_Datapath/RegisterFile/N23430 ) );
  AOI22_X1 U86711 ( .A1(n105293), .A2(n74069), .B1(n105290), .B2(n81308), .ZN(
        n97939) );
  OAI21_X1 U86712 ( .B1(n106100), .B2(n105295), .A(n97940), .ZN(
        \DLX_Datapath/RegisterFile/N23429 ) );
  AOI22_X1 U86713 ( .A1(n105292), .A2(n70656), .B1(n97935), .B2(n94516), .ZN(
        n97940) );
  OAI21_X1 U86714 ( .B1(n106256), .B2(n105295), .A(n97941), .ZN(
        \DLX_Datapath/RegisterFile/N23428 ) );
  AOI22_X1 U86715 ( .A1(n105292), .A2(n74210), .B1(n97935), .B2(n81272), .ZN(
        n97941) );
  OAI21_X1 U86716 ( .B1(n81629), .B2(n105295), .A(n97942), .ZN(
        \DLX_Datapath/RegisterFile/N23427 ) );
  AOI22_X1 U86717 ( .A1(n105293), .A2(n110901), .B1(n105291), .B2(n94519), 
        .ZN(n97942) );
  OAI21_X1 U86718 ( .B1(n106331), .B2(n105295), .A(n97943), .ZN(
        \DLX_Datapath/RegisterFile/N23426 ) );
  AOI22_X1 U86719 ( .A1(n105292), .A2(n110496), .B1(n105291), .B2(n80192), 
        .ZN(n97943) );
  OAI21_X1 U86720 ( .B1(n106192), .B2(n105294), .A(n97944), .ZN(
        \DLX_Datapath/RegisterFile/N23425 ) );
  AOI22_X1 U86721 ( .A1(n97934), .A2(n111039), .B1(n105291), .B2(n81474), .ZN(
        n97944) );
  OAI21_X1 U86722 ( .B1(n106131), .B2(n105294), .A(n97945), .ZN(
        \DLX_Datapath/RegisterFile/N23424 ) );
  AOI22_X1 U86723 ( .A1(n97934), .A2(n110599), .B1(n105291), .B2(n94523), .ZN(
        n97945) );
  OAI21_X1 U86724 ( .B1(n106187), .B2(n105294), .A(n97946), .ZN(
        \DLX_Datapath/RegisterFile/N23423 ) );
  AOI22_X1 U86725 ( .A1(n105293), .A2(n111038), .B1(n105291), .B2(n106061), 
        .ZN(n97946) );
  OAI21_X1 U86726 ( .B1(n106165), .B2(n105294), .A(n97947), .ZN(
        \DLX_Datapath/RegisterFile/N23422 ) );
  AOI22_X1 U86727 ( .A1(n97934), .A2(n111040), .B1(n105291), .B2(n81347), .ZN(
        n97947) );
  OAI21_X1 U86728 ( .B1(n106106), .B2(n105294), .A(n97948), .ZN(
        \DLX_Datapath/RegisterFile/N23421 ) );
  AOI22_X1 U86729 ( .A1(n97934), .A2(n111035), .B1(n105291), .B2(n94527), .ZN(
        n97948) );
  OAI21_X1 U86730 ( .B1(n106220), .B2(n105294), .A(n97949), .ZN(
        \DLX_Datapath/RegisterFile/N23420 ) );
  AOI22_X1 U86731 ( .A1(n97934), .A2(n109958), .B1(n105291), .B2(n81297), .ZN(
        n97949) );
  OAI21_X1 U86732 ( .B1(n106110), .B2(n105294), .A(n97950), .ZN(
        \DLX_Datapath/RegisterFile/N23419 ) );
  AOI22_X1 U86733 ( .A1(n97934), .A2(n109841), .B1(n105291), .B2(n94530), .ZN(
        n97950) );
  OAI21_X1 U86734 ( .B1(n106232), .B2(n105294), .A(n97951), .ZN(
        \DLX_Datapath/RegisterFile/N23418 ) );
  AOI22_X1 U86735 ( .A1(n105292), .A2(n108215), .B1(n105291), .B2(n81286), 
        .ZN(n97951) );
  OAI21_X1 U86736 ( .B1(n106173), .B2(n105294), .A(n97952), .ZN(
        \DLX_Datapath/RegisterFile/N23417 ) );
  AOI22_X1 U86737 ( .A1(n105292), .A2(n108338), .B1(n105291), .B2(n106168), 
        .ZN(n97952) );
  OAI21_X1 U86738 ( .B1(n106237), .B2(n105294), .A(n97953), .ZN(
        \DLX_Datapath/RegisterFile/N23416 ) );
  AOI22_X1 U86739 ( .A1(n105292), .A2(n108449), .B1(n105291), .B2(n81283), 
        .ZN(n97953) );
  OAI21_X1 U86740 ( .B1(n106069), .B2(n105294), .A(n97954), .ZN(
        \DLX_Datapath/RegisterFile/N23415 ) );
  AOI22_X1 U86741 ( .A1(n97934), .A2(n107687), .B1(n105291), .B2(n81453), .ZN(
        n97954) );
  OAI21_X1 U86742 ( .B1(n106199), .B2(n105294), .A(n97955), .ZN(
        \DLX_Datapath/RegisterFile/N23414 ) );
  AOI22_X1 U86743 ( .A1(n105292), .A2(n109605), .B1(n105290), .B2(n94536), 
        .ZN(n97955) );
  OAI21_X1 U86744 ( .B1(n106246), .B2(n105295), .A(n97956), .ZN(
        \DLX_Datapath/RegisterFile/N23413 ) );
  AOI22_X1 U86745 ( .A1(n105293), .A2(n108566), .B1(n105290), .B2(n106241), 
        .ZN(n97956) );
  OAI21_X1 U86746 ( .B1(n106160), .B2(n105295), .A(n97957), .ZN(
        \DLX_Datapath/RegisterFile/N23412 ) );
  AOI22_X1 U86747 ( .A1(n105292), .A2(n109710), .B1(n105290), .B2(n81351), 
        .ZN(n97957) );
  OAI21_X1 U86748 ( .B1(n106115), .B2(n105294), .A(n97958), .ZN(
        \DLX_Datapath/RegisterFile/N23411 ) );
  AOI22_X1 U86749 ( .A1(n105293), .A2(n109494), .B1(n105290), .B2(n106020), 
        .ZN(n97958) );
  OAI21_X1 U86750 ( .B1(n106011), .B2(n105295), .A(n97959), .ZN(
        \DLX_Datapath/RegisterFile/N23410 ) );
  AOI22_X1 U86751 ( .A1(n105292), .A2(n109031), .B1(n105290), .B2(n94541), 
        .ZN(n97959) );
  OAI21_X1 U86752 ( .B1(n106261), .B2(n105295), .A(n97960), .ZN(
        \DLX_Datapath/RegisterFile/N23409 ) );
  AOI22_X1 U86753 ( .A1(n105293), .A2(n109379), .B1(n105290), .B2(n81269), 
        .ZN(n97960) );
  OAI21_X1 U86754 ( .B1(n106045), .B2(n105294), .A(n97961), .ZN(
        \DLX_Datapath/RegisterFile/N23408 ) );
  AOI22_X1 U86755 ( .A1(n105292), .A2(n109261), .B1(n105290), .B2(n105624), 
        .ZN(n97961) );
  OAI21_X1 U86756 ( .B1(n106050), .B2(n105295), .A(n97962), .ZN(
        \DLX_Datapath/RegisterFile/N23407 ) );
  AOI22_X1 U86757 ( .A1(n105293), .A2(n109152), .B1(n105290), .B2(n94546), 
        .ZN(n97962) );
  OAI21_X1 U86758 ( .B1(n106096), .B2(n105294), .A(n97963), .ZN(
        \DLX_Datapath/RegisterFile/N23406 ) );
  AOI22_X1 U86759 ( .A1(n105292), .A2(n108688), .B1(n105290), .B2(n94548), 
        .ZN(n97963) );
  OAI21_X1 U86760 ( .B1(n106055), .B2(n105295), .A(n97964), .ZN(
        \DLX_Datapath/RegisterFile/N23405 ) );
  AOI22_X1 U86761 ( .A1(n105293), .A2(n108915), .B1(n105290), .B2(n81783), 
        .ZN(n97964) );
  OAI21_X1 U86762 ( .B1(n105216), .B2(n105295), .A(n97965), .ZN(
        \DLX_Datapath/RegisterFile/N23404 ) );
  AOI22_X1 U86763 ( .A1(n105293), .A2(n108803), .B1(n105290), .B2(n80188), 
        .ZN(n97965) );
  OAI21_X1 U86764 ( .B1(n106269), .B2(n105294), .A(n97966), .ZN(
        \DLX_Datapath/RegisterFile/N23403 ) );
  AOI22_X1 U86765 ( .A1(n105292), .A2(n107343), .B1(n105290), .B2(n81265), 
        .ZN(n97966) );
  NOR2_X1 U86766 ( .A1(n97967), .A2(n97968), .ZN(n97935) );
  AOI21_X1 U86767 ( .B1(n97572), .B2(n94771), .A(n97968), .ZN(n97934) );
  NOR2_X1 U86768 ( .A1(n97932), .A2(n105094), .ZN(n97968) );
  NAND2_X1 U86769 ( .A1(n97674), .A2(n107022), .ZN(n97572) );
  NAND2_X1 U86770 ( .A1(n105126), .A2(n94772), .ZN(n97932) );
  OAI21_X1 U86771 ( .B1(n106149), .B2(n105289), .A(n97970), .ZN(
        \DLX_Datapath/RegisterFile/N23402 ) );
  AOI22_X1 U86772 ( .A1(n105288), .A2(n107901), .B1(n105285), .B2(n94559), 
        .ZN(n97970) );
  OAI21_X1 U86773 ( .B1(n105969), .B2(n105289), .A(n97973), .ZN(
        \DLX_Datapath/RegisterFile/N23401 ) );
  AOI22_X1 U86774 ( .A1(n105287), .A2(n107997), .B1(n105284), .B2(n94562), 
        .ZN(n97973) );
  OAI21_X1 U86775 ( .B1(n106138), .B2(n105289), .A(n97974), .ZN(
        \DLX_Datapath/RegisterFile/N23400 ) );
  AOI22_X1 U86776 ( .A1(n105288), .A2(n107268), .B1(n105285), .B2(n94564), 
        .ZN(n97974) );
  OAI21_X1 U86777 ( .B1(n106210), .B2(n105289), .A(n97975), .ZN(
        \DLX_Datapath/RegisterFile/N23399 ) );
  AOI22_X1 U86778 ( .A1(n105287), .A2(n107805), .B1(n105284), .B2(n94566), 
        .ZN(n97975) );
  OAI21_X1 U86779 ( .B1(n106205), .B2(n105289), .A(n97976), .ZN(
        \DLX_Datapath/RegisterFile/N23398 ) );
  AOI22_X1 U86780 ( .A1(n105288), .A2(n110702), .B1(n105285), .B2(n94568), 
        .ZN(n97976) );
  OAI21_X1 U86781 ( .B1(n106101), .B2(n105289), .A(n97977), .ZN(
        \DLX_Datapath/RegisterFile/N23397 ) );
  AOI22_X1 U86782 ( .A1(n105287), .A2(n108105), .B1(n105284), .B2(n94570), 
        .ZN(n97977) );
  OAI21_X1 U86783 ( .B1(n106256), .B2(n105289), .A(n97978), .ZN(
        \DLX_Datapath/RegisterFile/N23396 ) );
  AOI22_X1 U86784 ( .A1(n105288), .A2(n110804), .B1(n105285), .B2(n94572), 
        .ZN(n97978) );
  OAI21_X1 U86785 ( .B1(n81629), .B2(n105289), .A(n97979), .ZN(
        \DLX_Datapath/RegisterFile/N23395 ) );
  AOI22_X1 U86786 ( .A1(n105287), .A2(n110902), .B1(n105284), .B2(n94574), 
        .ZN(n97979) );
  OAI21_X1 U86787 ( .B1(n106330), .B2(n105289), .A(n97980), .ZN(
        \DLX_Datapath/RegisterFile/N23394 ) );
  AOI22_X1 U86788 ( .A1(n105287), .A2(n110497), .B1(n105284), .B2(n94576), 
        .ZN(n97980) );
  OAI21_X1 U86789 ( .B1(n106192), .B2(n105289), .A(n97981), .ZN(
        \DLX_Datapath/RegisterFile/N23393 ) );
  AOI22_X1 U86790 ( .A1(n105286), .A2(n110280), .B1(n105283), .B2(n94578), 
        .ZN(n97981) );
  OAI21_X1 U86791 ( .B1(n106131), .B2(n105289), .A(n97982), .ZN(
        \DLX_Datapath/RegisterFile/N23392 ) );
  AOI22_X1 U86792 ( .A1(n105286), .A2(n110600), .B1(n105283), .B2(n94580), 
        .ZN(n97982) );
  OAI21_X1 U86793 ( .B1(n106187), .B2(n105289), .A(n97983), .ZN(
        \DLX_Datapath/RegisterFile/N23391 ) );
  AOI22_X1 U86794 ( .A1(n105286), .A2(n110389), .B1(n105283), .B2(n94582), 
        .ZN(n97983) );
  OAI21_X1 U86795 ( .B1(n106165), .B2(n105289), .A(n97984), .ZN(
        \DLX_Datapath/RegisterFile/N23390 ) );
  AOI22_X1 U86796 ( .A1(n105286), .A2(n110067), .B1(n105283), .B2(n94584), 
        .ZN(n97984) );
  OAI21_X1 U86797 ( .B1(n106106), .B2(n105289), .A(n97985), .ZN(
        \DLX_Datapath/RegisterFile/N23389 ) );
  AOI22_X1 U86798 ( .A1(n105286), .A2(n110174), .B1(n105283), .B2(n94586), 
        .ZN(n97985) );
  OAI21_X1 U86799 ( .B1(n106220), .B2(n105289), .A(n97986), .ZN(
        \DLX_Datapath/RegisterFile/N23388 ) );
  AOI22_X1 U86800 ( .A1(n105286), .A2(n109959), .B1(n105283), .B2(n94588), 
        .ZN(n97986) );
  OAI21_X1 U86801 ( .B1(n106111), .B2(n105289), .A(n97987), .ZN(
        \DLX_Datapath/RegisterFile/N23387 ) );
  AOI22_X1 U86802 ( .A1(n105286), .A2(n109842), .B1(n105283), .B2(n94590), 
        .ZN(n97987) );
  OAI21_X1 U86803 ( .B1(n106232), .B2(n105289), .A(n97988), .ZN(
        \DLX_Datapath/RegisterFile/N23386 ) );
  AOI22_X1 U86804 ( .A1(n105286), .A2(n108216), .B1(n105283), .B2(n94592), 
        .ZN(n97988) );
  OAI21_X1 U86805 ( .B1(n106173), .B2(n105289), .A(n97989), .ZN(
        \DLX_Datapath/RegisterFile/N23385 ) );
  AOI22_X1 U86806 ( .A1(n105286), .A2(n108339), .B1(n105283), .B2(n94594), 
        .ZN(n97989) );
  OAI21_X1 U86807 ( .B1(n106237), .B2(n105289), .A(n97990), .ZN(
        \DLX_Datapath/RegisterFile/N23384 ) );
  AOI22_X1 U86808 ( .A1(n105286), .A2(n108450), .B1(n105283), .B2(n94596), 
        .ZN(n97990) );
  OAI21_X1 U86809 ( .B1(n106069), .B2(n105289), .A(n97991), .ZN(
        \DLX_Datapath/RegisterFile/N23383 ) );
  AOI22_X1 U86810 ( .A1(n105286), .A2(n107688), .B1(n105283), .B2(n94598), 
        .ZN(n97991) );
  OAI21_X1 U86811 ( .B1(n106199), .B2(n105289), .A(n97992), .ZN(
        \DLX_Datapath/RegisterFile/N23382 ) );
  AOI22_X1 U86812 ( .A1(n105287), .A2(n72600), .B1(n105284), .B2(n94600), .ZN(
        n97992) );
  OAI21_X1 U86813 ( .B1(n106246), .B2(n97969), .A(n97993), .ZN(
        \DLX_Datapath/RegisterFile/N23381 ) );
  AOI22_X1 U86814 ( .A1(n105288), .A2(n108567), .B1(n105285), .B2(n94602), 
        .ZN(n97993) );
  OAI21_X1 U86815 ( .B1(n106160), .B2(n97969), .A(n97994), .ZN(
        \DLX_Datapath/RegisterFile/N23380 ) );
  AOI22_X1 U86816 ( .A1(n105287), .A2(n109711), .B1(n105284), .B2(n94604), 
        .ZN(n97994) );
  OAI21_X1 U86817 ( .B1(n106116), .B2(n97969), .A(n97995), .ZN(
        \DLX_Datapath/RegisterFile/N23379 ) );
  AOI22_X1 U86818 ( .A1(n105288), .A2(n109495), .B1(n105285), .B2(n94606), 
        .ZN(n97995) );
  OAI21_X1 U86819 ( .B1(n106011), .B2(n97969), .A(n97996), .ZN(
        \DLX_Datapath/RegisterFile/N23378 ) );
  AOI22_X1 U86820 ( .A1(n105287), .A2(n109032), .B1(n105284), .B2(n94608), 
        .ZN(n97996) );
  OAI21_X1 U86821 ( .B1(n106261), .B2(n97969), .A(n97997), .ZN(
        \DLX_Datapath/RegisterFile/N23377 ) );
  AOI22_X1 U86822 ( .A1(n105288), .A2(n109380), .B1(n105285), .B2(n94610), 
        .ZN(n97997) );
  OAI21_X1 U86823 ( .B1(n106045), .B2(n105289), .A(n97998), .ZN(
        \DLX_Datapath/RegisterFile/N23376 ) );
  AOI22_X1 U86824 ( .A1(n105287), .A2(n109262), .B1(n105284), .B2(n94612), 
        .ZN(n97998) );
  OAI21_X1 U86825 ( .B1(n106050), .B2(n97969), .A(n97999), .ZN(
        \DLX_Datapath/RegisterFile/N23375 ) );
  AOI22_X1 U86826 ( .A1(n105288), .A2(n109153), .B1(n105285), .B2(n94614), 
        .ZN(n97999) );
  OAI21_X1 U86827 ( .B1(n106096), .B2(n97969), .A(n98000), .ZN(
        \DLX_Datapath/RegisterFile/N23374 ) );
  AOI22_X1 U86828 ( .A1(n105287), .A2(n108689), .B1(n105284), .B2(n94616), 
        .ZN(n98000) );
  OAI21_X1 U86829 ( .B1(n106055), .B2(n97969), .A(n98001), .ZN(
        \DLX_Datapath/RegisterFile/N23373 ) );
  AOI22_X1 U86830 ( .A1(n105288), .A2(n108916), .B1(n105285), .B2(n94618), 
        .ZN(n98001) );
  OAI21_X1 U86831 ( .B1(n105216), .B2(n105289), .A(n98002), .ZN(
        \DLX_Datapath/RegisterFile/N23372 ) );
  AOI22_X1 U86832 ( .A1(n105288), .A2(n108804), .B1(n105285), .B2(n94620), 
        .ZN(n98002) );
  OAI21_X1 U86833 ( .B1(n106269), .B2(n105289), .A(n98003), .ZN(
        \DLX_Datapath/RegisterFile/N23371 ) );
  AOI22_X1 U86834 ( .A1(n105287), .A2(n107344), .B1(n105284), .B2(n94622), 
        .ZN(n98003) );
  NOR2_X1 U86837 ( .A1(n97969), .A2(n105095), .ZN(n98004) );
  NAND2_X1 U86838 ( .A1(n105125), .A2(n94810), .ZN(n97969) );
  OAI21_X1 U86839 ( .B1(n106149), .B2(n106091), .A(n98006), .ZN(
        \DLX_Datapath/RegisterFile/N23370 ) );
  AOI22_X1 U86840 ( .A1(n70369), .A2(n81421), .B1(n81521), .B2(n81422), .ZN(
        n98006) );
  OAI21_X1 U86841 ( .B1(n106091), .B2(n81651), .A(n98007), .ZN(
        \DLX_Datapath/RegisterFile/N23369 ) );
  AOI22_X1 U86842 ( .A1(n70511), .A2(n106090), .B1(n81653), .B2(n81422), .ZN(
        n98007) );
  OAI21_X1 U86843 ( .B1(n106138), .B2(n106091), .A(n98008), .ZN(
        \DLX_Datapath/RegisterFile/N23368 ) );
  AOI22_X1 U86844 ( .A1(n69564), .A2(n106090), .B1(n106088), .B2(n81380), .ZN(
        n98008) );
  OAI21_X1 U86845 ( .B1(n106210), .B2(n106092), .A(n98009), .ZN(
        \DLX_Datapath/RegisterFile/N23367 ) );
  AOI22_X1 U86846 ( .A1(n70225), .A2(n81421), .B1(n106088), .B2(n81377), .ZN(
        n98009) );
  OAI21_X1 U86847 ( .B1(n106101), .B2(n106092), .A(n98010), .ZN(
        \DLX_Datapath/RegisterFile/N23365 ) );
  AOI22_X1 U86848 ( .A1(n70658), .A2(n106090), .B1(n106088), .B2(n81410), .ZN(
        n98010) );
  OAI21_X1 U86849 ( .B1(n106256), .B2(n106092), .A(n98011), .ZN(
        \DLX_Datapath/RegisterFile/N23364 ) );
  AOI22_X1 U86850 ( .A1(n74212), .A2(n81421), .B1(n81700), .B2(n81422), .ZN(
        n98011) );
  OAI21_X1 U86851 ( .B1(n106091), .B2(n105991), .A(n98012), .ZN(
        \DLX_Datapath/RegisterFile/N23363 ) );
  AOI22_X1 U86852 ( .A1(n106089), .A2(n110903), .B1(n81632), .B2(n106088), 
        .ZN(n98012) );
  OAI21_X1 U86853 ( .B1(n106192), .B2(n106092), .A(n98013), .ZN(
        \DLX_Datapath/RegisterFile/N23361 ) );
  AOI22_X1 U86854 ( .A1(n106089), .A2(n110281), .B1(n106088), .B2(n81317), 
        .ZN(n98013) );
  OAI21_X1 U86855 ( .B1(n106165), .B2(n106092), .A(n98014), .ZN(
        \DLX_Datapath/RegisterFile/N23358 ) );
  AOI22_X1 U86856 ( .A1(n106089), .A2(n110068), .B1(n81604), .B2(n81422), .ZN(
        n98014) );
  OAI21_X1 U86857 ( .B1(n106220), .B2(n106092), .A(n98015), .ZN(
        \DLX_Datapath/RegisterFile/N23356 ) );
  AOI22_X1 U86858 ( .A1(n106090), .A2(n109960), .B1(n106088), .B2(n81402), 
        .ZN(n98015) );
  OAI21_X1 U86859 ( .B1(n106111), .B2(n106092), .A(n98016), .ZN(
        \DLX_Datapath/RegisterFile/N23355 ) );
  AOI22_X1 U86860 ( .A1(n106090), .A2(n109843), .B1(n106088), .B2(n81400), 
        .ZN(n98016) );
  OAI21_X1 U86861 ( .B1(n106092), .B2(n106070), .A(n98017), .ZN(
        \DLX_Datapath/RegisterFile/N23351 ) );
  AOI22_X1 U86862 ( .A1(n106090), .A2(n107689), .B1(n81506), .B2(n81422), .ZN(
        n98017) );
  OAI21_X1 U86863 ( .B1(n106116), .B2(n106092), .A(n98018), .ZN(
        \DLX_Datapath/RegisterFile/N23347 ) );
  AOI22_X1 U86864 ( .A1(n106090), .A2(n109496), .B1(n106088), .B2(n81396), 
        .ZN(n98018) );
  OAI21_X1 U86865 ( .B1(n106011), .B2(n106092), .A(n98019), .ZN(
        \DLX_Datapath/RegisterFile/N23346 ) );
  AOI22_X1 U86866 ( .A1(n106090), .A2(n109033), .B1(n81590), .B2(n81422), .ZN(
        n98019) );
  OAI21_X1 U86867 ( .B1(n106091), .B2(n81509), .A(n98020), .ZN(
        \DLX_Datapath/RegisterFile/N23344 ) );
  AOI22_X1 U86868 ( .A1(n106090), .A2(n109263), .B1(n81511), .B2(n106088), 
        .ZN(n98020) );
  OAI21_X1 U86869 ( .B1(n106092), .B2(n106051), .A(n98021), .ZN(
        \DLX_Datapath/RegisterFile/N23343 ) );
  AOI22_X1 U86870 ( .A1(n106090), .A2(n109154), .B1(n81503), .B2(n81422), .ZN(
        n98021) );
  OAI21_X1 U86871 ( .B1(n106092), .B2(n81498), .A(n98022), .ZN(
        \DLX_Datapath/RegisterFile/N23341 ) );
  AOI22_X1 U86872 ( .A1(n106090), .A2(n108917), .B1(n81500), .B2(n106088), 
        .ZN(n98022) );
  OAI21_X1 U86873 ( .B1(n106269), .B2(n106092), .A(n98023), .ZN(
        \DLX_Datapath/RegisterFile/N23339 ) );
  AOI22_X1 U86874 ( .A1(n106089), .A2(n107345), .B1(n106087), .B2(n81327), 
        .ZN(n98023) );
  NOR2_X1 U86875 ( .A1(n97967), .A2(n98024), .ZN(n81422) );
  NOR2_X1 U86876 ( .A1(n98005), .A2(n98024), .ZN(n81421) );
  NOR2_X1 U86877 ( .A1(n81419), .A2(n105094), .ZN(n98024) );
  NAND2_X1 U86878 ( .A1(n105126), .A2(n94853), .ZN(n81419) );
  OAI21_X1 U86879 ( .B1(n106149), .B2(n105282), .A(n98026), .ZN(
        \DLX_Datapath/RegisterFile/N23338 ) );
  AOI22_X1 U86880 ( .A1(n105280), .A2(n94667), .B1(n105278), .B2(n107902), 
        .ZN(n98026) );
  OAI21_X1 U86881 ( .B1(n105968), .B2(n105282), .A(n98029), .ZN(
        \DLX_Datapath/RegisterFile/N23337 ) );
  AOI22_X1 U86882 ( .A1(n98027), .A2(n94670), .B1(n105277), .B2(n107998), .ZN(
        n98029) );
  OAI21_X1 U86883 ( .B1(n106138), .B2(n105282), .A(n98030), .ZN(
        \DLX_Datapath/RegisterFile/N23336 ) );
  AOI22_X1 U86884 ( .A1(n105280), .A2(n94672), .B1(n105278), .B2(n107269), 
        .ZN(n98030) );
  OAI21_X1 U86885 ( .B1(n106210), .B2(n105282), .A(n98031), .ZN(
        \DLX_Datapath/RegisterFile/N23335 ) );
  AOI22_X1 U86886 ( .A1(n98027), .A2(n94674), .B1(n105277), .B2(n107806), .ZN(
        n98031) );
  OAI21_X1 U86887 ( .B1(n106205), .B2(n105282), .A(n98032), .ZN(
        \DLX_Datapath/RegisterFile/N23334 ) );
  AOI22_X1 U86888 ( .A1(n105280), .A2(n94676), .B1(n105278), .B2(n110703), 
        .ZN(n98032) );
  OAI21_X1 U86889 ( .B1(n106101), .B2(n105282), .A(n98033), .ZN(
        \DLX_Datapath/RegisterFile/N23333 ) );
  AOI22_X1 U86890 ( .A1(n98027), .A2(n94678), .B1(n105277), .B2(n108106), .ZN(
        n98033) );
  OAI21_X1 U86891 ( .B1(n106256), .B2(n105282), .A(n98034), .ZN(
        \DLX_Datapath/RegisterFile/N23332 ) );
  AOI22_X1 U86892 ( .A1(n105280), .A2(n94680), .B1(n105278), .B2(n110805), 
        .ZN(n98034) );
  OAI21_X1 U86893 ( .B1(n105990), .B2(n105282), .A(n98035), .ZN(
        \DLX_Datapath/RegisterFile/N23331 ) );
  AOI22_X1 U86894 ( .A1(n105279), .A2(n94682), .B1(n105277), .B2(n110904), 
        .ZN(n98035) );
  OAI21_X1 U86895 ( .B1(n106330), .B2(n105282), .A(n98036), .ZN(
        \DLX_Datapath/RegisterFile/N23330 ) );
  AOI22_X1 U86896 ( .A1(n98027), .A2(n94684), .B1(n105277), .B2(n110499), .ZN(
        n98036) );
  OAI21_X1 U86897 ( .B1(n106192), .B2(n105281), .A(n98037), .ZN(
        \DLX_Datapath/RegisterFile/N23329 ) );
  AOI22_X1 U86898 ( .A1(n105279), .A2(n94686), .B1(n98028), .B2(n110282), .ZN(
        n98037) );
  OAI21_X1 U86899 ( .B1(n106131), .B2(n105281), .A(n98038), .ZN(
        \DLX_Datapath/RegisterFile/N23328 ) );
  AOI22_X1 U86900 ( .A1(n105279), .A2(n94688), .B1(n98028), .B2(n110602), .ZN(
        n98038) );
  OAI21_X1 U86901 ( .B1(n106187), .B2(n105281), .A(n98039), .ZN(
        \DLX_Datapath/RegisterFile/N23327 ) );
  AOI22_X1 U86902 ( .A1(n105279), .A2(n94690), .B1(n98028), .B2(n110391), .ZN(
        n98039) );
  OAI21_X1 U86903 ( .B1(n106165), .B2(n105281), .A(n98040), .ZN(
        \DLX_Datapath/RegisterFile/N23326 ) );
  AOI22_X1 U86904 ( .A1(n105279), .A2(n94692), .B1(n105277), .B2(n110069), 
        .ZN(n98040) );
  OAI21_X1 U86905 ( .B1(n106106), .B2(n105281), .A(n98041), .ZN(
        \DLX_Datapath/RegisterFile/N23325 ) );
  AOI22_X1 U86906 ( .A1(n105279), .A2(n94694), .B1(n98028), .B2(n110176), .ZN(
        n98041) );
  OAI21_X1 U86907 ( .B1(n106220), .B2(n105281), .A(n98042), .ZN(
        \DLX_Datapath/RegisterFile/N23324 ) );
  AOI22_X1 U86908 ( .A1(n105279), .A2(n94696), .B1(n98028), .B2(n109961), .ZN(
        n98042) );
  OAI21_X1 U86909 ( .B1(n106111), .B2(n105281), .A(n98043), .ZN(
        \DLX_Datapath/RegisterFile/N23323 ) );
  AOI22_X1 U86910 ( .A1(n105279), .A2(n94698), .B1(n98028), .B2(n109844), .ZN(
        n98043) );
  OAI21_X1 U86911 ( .B1(n106232), .B2(n105281), .A(n98044), .ZN(
        \DLX_Datapath/RegisterFile/N23322 ) );
  AOI22_X1 U86912 ( .A1(n105279), .A2(n94700), .B1(n98028), .B2(n108218), .ZN(
        n98044) );
  OAI21_X1 U86913 ( .B1(n106173), .B2(n105281), .A(n98045), .ZN(
        \DLX_Datapath/RegisterFile/N23321 ) );
  AOI22_X1 U86914 ( .A1(n105279), .A2(n94702), .B1(n98028), .B2(n108341), .ZN(
        n98045) );
  OAI21_X1 U86915 ( .B1(n106237), .B2(n105281), .A(n98046), .ZN(
        \DLX_Datapath/RegisterFile/N23320 ) );
  AOI22_X1 U86916 ( .A1(n105279), .A2(n94704), .B1(n105278), .B2(n108452), 
        .ZN(n98046) );
  OAI21_X1 U86917 ( .B1(n81451), .B2(n105281), .A(n98047), .ZN(
        \DLX_Datapath/RegisterFile/N23319 ) );
  AOI22_X1 U86918 ( .A1(n105279), .A2(n94706), .B1(n105277), .B2(n107690), 
        .ZN(n98047) );
  OAI21_X1 U86919 ( .B1(n106199), .B2(n105281), .A(n98048), .ZN(
        \DLX_Datapath/RegisterFile/N23318 ) );
  AOI22_X1 U86920 ( .A1(n98027), .A2(n94708), .B1(n105277), .B2(n109607), .ZN(
        n98048) );
  OAI21_X1 U86921 ( .B1(n106246), .B2(n105282), .A(n98049), .ZN(
        \DLX_Datapath/RegisterFile/N23317 ) );
  AOI22_X1 U86922 ( .A1(n105280), .A2(n94710), .B1(n105278), .B2(n108569), 
        .ZN(n98049) );
  OAI21_X1 U86923 ( .B1(n106160), .B2(n105282), .A(n98050), .ZN(
        \DLX_Datapath/RegisterFile/N23316 ) );
  AOI22_X1 U86924 ( .A1(n98027), .A2(n94712), .B1(n105277), .B2(n109713), .ZN(
        n98050) );
  OAI21_X1 U86925 ( .B1(n106116), .B2(n105281), .A(n98051), .ZN(
        \DLX_Datapath/RegisterFile/N23315 ) );
  AOI22_X1 U86926 ( .A1(n105280), .A2(n94714), .B1(n105278), .B2(n109497), 
        .ZN(n98051) );
  OAI21_X1 U86927 ( .B1(n106011), .B2(n105282), .A(n98052), .ZN(
        \DLX_Datapath/RegisterFile/N23314 ) );
  AOI22_X1 U86928 ( .A1(n98027), .A2(n81259), .B1(n105277), .B2(n109034), .ZN(
        n98052) );
  OAI21_X1 U86929 ( .B1(n106261), .B2(n105282), .A(n98053), .ZN(
        \DLX_Datapath/RegisterFile/N23313 ) );
  AOI22_X1 U86930 ( .A1(n105280), .A2(n94717), .B1(n105278), .B2(n109382), 
        .ZN(n98053) );
  OAI21_X1 U86931 ( .B1(n106045), .B2(n105281), .A(n98054), .ZN(
        \DLX_Datapath/RegisterFile/N23312 ) );
  AOI22_X1 U86932 ( .A1(n105279), .A2(n94719), .B1(n105277), .B2(n109264), 
        .ZN(n98054) );
  OAI21_X1 U86933 ( .B1(n106051), .B2(n105282), .A(n98055), .ZN(
        \DLX_Datapath/RegisterFile/N23311 ) );
  AOI22_X1 U86934 ( .A1(n105280), .A2(n94721), .B1(n105278), .B2(n109155), 
        .ZN(n98055) );
  OAI21_X1 U86935 ( .B1(n106096), .B2(n105281), .A(n98056), .ZN(
        \DLX_Datapath/RegisterFile/N23310 ) );
  AOI22_X1 U86936 ( .A1(n98027), .A2(n94723), .B1(n105277), .B2(n108691), .ZN(
        n98056) );
  OAI21_X1 U86937 ( .B1(n106055), .B2(n105282), .A(n98057), .ZN(
        \DLX_Datapath/RegisterFile/N23309 ) );
  AOI22_X1 U86938 ( .A1(n105280), .A2(n94725), .B1(n105278), .B2(n108918), 
        .ZN(n98057) );
  OAI21_X1 U86939 ( .B1(n105216), .B2(n105282), .A(n98058), .ZN(
        \DLX_Datapath/RegisterFile/N23308 ) );
  AOI22_X1 U86940 ( .A1(n105280), .A2(n94727), .B1(n105278), .B2(n108806), 
        .ZN(n98058) );
  OAI21_X1 U86941 ( .B1(n106269), .B2(n105281), .A(n98059), .ZN(
        \DLX_Datapath/RegisterFile/N23307 ) );
  AOI22_X1 U86942 ( .A1(n105280), .A2(n94729), .B1(n105277), .B2(n107346), 
        .ZN(n98059) );
  NOR2_X1 U86943 ( .A1(n98005), .A2(n98060), .ZN(n98028) );
  AOI21_X1 U86944 ( .B1(n105205), .B2(n97967), .A(n105601), .ZN(n98005) );
  NOR2_X1 U86945 ( .A1(n97967), .A2(n98060), .ZN(n98027) );
  NOR2_X1 U86946 ( .A1(n98025), .A2(n105093), .ZN(n98060) );
  OR2_X1 U86947 ( .A1(n97674), .A2(n94848), .ZN(n97967) );
  NAND2_X1 U86948 ( .A1(n98061), .A2(n107028), .ZN(n97674) );
  NOR2_X1 U86949 ( .A1(n96488), .A2(n106763), .ZN(n98061) );
  NAND2_X1 U86950 ( .A1(n94892), .A2(n105125), .ZN(n98025) );
  NOR2_X1 U86951 ( .A1(n95991), .A2(n104732), .ZN(n97575) );
  NAND2_X1 U86952 ( .A1(n94895), .A2(n95412), .ZN(n95991) );
  OAI21_X1 U86953 ( .B1(n106229), .B2(n81358), .A(n98062), .ZN(
        \DLX_Datapath/RegisterFile/N23306 ) );
  AOI22_X1 U86954 ( .A1(n81360), .A2(n106226), .B1(n106224), .B2(n107903), 
        .ZN(n98062) );
  OAI21_X1 U86955 ( .B1(n106229), .B2(n105971), .A(n98063), .ZN(
        \DLX_Datapath/RegisterFile/N23305 ) );
  AOI22_X1 U86956 ( .A1(n94511), .A2(n106227), .B1(n106224), .B2(n107999), 
        .ZN(n98063) );
  OAI21_X1 U86957 ( .B1(n106229), .B2(n106137), .A(n98064), .ZN(
        \DLX_Datapath/RegisterFile/N23304 ) );
  AOI22_X1 U86958 ( .A1(n81539), .A2(n106226), .B1(n106224), .B2(n107270), 
        .ZN(n98064) );
  OAI21_X1 U86959 ( .B1(n106229), .B2(n106209), .A(n98065), .ZN(
        \DLX_Datapath/RegisterFile/N23303 ) );
  AOI22_X1 U86960 ( .A1(n81301), .A2(n106228), .B1(n106225), .B2(n107807), 
        .ZN(n98065) );
  OAI21_X1 U86961 ( .B1(n106229), .B2(n106099), .A(n98066), .ZN(
        \DLX_Datapath/RegisterFile/N23301 ) );
  AOI22_X1 U86962 ( .A1(n94516), .A2(n106228), .B1(n106225), .B2(n108107), 
        .ZN(n98066) );
  OAI21_X1 U86963 ( .B1(n106229), .B2(n105990), .A(n98067), .ZN(
        \DLX_Datapath/RegisterFile/N23299 ) );
  AOI22_X1 U86964 ( .A1(n94519), .A2(n106228), .B1(n106225), .B2(n110905), 
        .ZN(n98067) );
  OAI21_X1 U86965 ( .B1(n106330), .B2(n106229), .A(n98068), .ZN(
        \DLX_Datapath/RegisterFile/N23298 ) );
  AOI22_X1 U86966 ( .A1(n106227), .A2(n80192), .B1(n106225), .B2(n110500), 
        .ZN(n98068) );
  OAI21_X1 U86967 ( .B1(n106229), .B2(n81315), .A(n98069), .ZN(
        \DLX_Datapath/RegisterFile/N23297 ) );
  AOI22_X1 U86968 ( .A1(n81474), .A2(n106227), .B1(n106225), .B2(n110283), 
        .ZN(n98069) );
  OAI21_X1 U86969 ( .B1(n106229), .B2(n106129), .A(n98070), .ZN(
        \DLX_Datapath/RegisterFile/N23296 ) );
  AOI22_X1 U86970 ( .A1(n94523), .A2(n106226), .B1(n106225), .B2(n110603), 
        .ZN(n98070) );
  OAI21_X1 U86971 ( .B1(n106229), .B2(n106185), .A(n98071), .ZN(
        \DLX_Datapath/RegisterFile/N23295 ) );
  AOI22_X1 U86972 ( .A1(n106060), .A2(n106228), .B1(n106225), .B2(n110392), 
        .ZN(n98071) );
  OAI21_X1 U86973 ( .B1(n106229), .B2(n81345), .A(n98072), .ZN(
        \DLX_Datapath/RegisterFile/N23294 ) );
  AOI22_X1 U86974 ( .A1(n81347), .A2(n106226), .B1(n106225), .B2(n110070), 
        .ZN(n98072) );
  OAI21_X1 U86975 ( .B1(n106229), .B2(n81403), .A(n98073), .ZN(
        \DLX_Datapath/RegisterFile/N23293 ) );
  AOI22_X1 U86976 ( .A1(n94527), .A2(n106226), .B1(n106225), .B2(n110177), 
        .ZN(n98073) );
  OAI21_X1 U86977 ( .B1(n106229), .B2(n106220), .A(n98074), .ZN(
        \DLX_Datapath/RegisterFile/N23292 ) );
  AOI22_X1 U86978 ( .A1(n81297), .A2(n106227), .B1(n106225), .B2(n109962), 
        .ZN(n98074) );
  OAI21_X1 U86979 ( .B1(n106229), .B2(n106110), .A(n98075), .ZN(
        \DLX_Datapath/RegisterFile/N23291 ) );
  AOI22_X1 U86980 ( .A1(n94530), .A2(n106226), .B1(n106225), .B2(n109845), 
        .ZN(n98075) );
  OAI21_X1 U86981 ( .B1(n106229), .B2(n81340), .A(n98076), .ZN(
        \DLX_Datapath/RegisterFile/N23289 ) );
  AOI22_X1 U86982 ( .A1(n106167), .A2(n106226), .B1(n106225), .B2(n108342), 
        .ZN(n98076) );
  OAI21_X1 U86983 ( .B1(n106229), .B2(n81451), .A(n98077), .ZN(
        \DLX_Datapath/RegisterFile/N23287 ) );
  AOI22_X1 U86984 ( .A1(n81453), .A2(n106228), .B1(n81291), .B2(n107691), .ZN(
        n98077) );
  OAI21_X1 U86985 ( .B1(n106229), .B2(n81310), .A(n98078), .ZN(
        \DLX_Datapath/RegisterFile/N23286 ) );
  AOI22_X1 U86986 ( .A1(n105626), .A2(n106228), .B1(n72603), .B2(n106224), 
        .ZN(n98078) );
  OAI21_X1 U86987 ( .B1(n106229), .B2(n81349), .A(n98079), .ZN(
        \DLX_Datapath/RegisterFile/N23284 ) );
  AOI22_X1 U86988 ( .A1(n81351), .A2(n106226), .B1(n72745), .B2(n106224), .ZN(
        n98079) );
  OAI21_X1 U86989 ( .B1(n106229), .B2(n81394), .A(n98080), .ZN(
        \DLX_Datapath/RegisterFile/N23283 ) );
  AOI22_X1 U86990 ( .A1(n106019), .A2(n106226), .B1(n81291), .B2(n109498), 
        .ZN(n98080) );
  OAI21_X1 U86991 ( .B1(n106011), .B2(n106229), .A(n98081), .ZN(
        \DLX_Datapath/RegisterFile/N23282 ) );
  AOI22_X1 U86992 ( .A1(n94541), .A2(n106227), .B1(n106225), .B2(n109035), 
        .ZN(n98081) );
  OAI21_X1 U86993 ( .B1(n106229), .B2(n81509), .A(n98082), .ZN(
        \DLX_Datapath/RegisterFile/N23280 ) );
  AOI22_X1 U86994 ( .A1(n105623), .A2(n106227), .B1(n81291), .B2(n109265), 
        .ZN(n98082) );
  OAI21_X1 U86995 ( .B1(n106229), .B2(n81501), .A(n98083), .ZN(
        \DLX_Datapath/RegisterFile/N23279 ) );
  AOI22_X1 U86996 ( .A1(n105622), .A2(n106228), .B1(n81291), .B2(n109156), 
        .ZN(n98083) );
  OAI21_X1 U86997 ( .B1(n106229), .B2(n81415), .A(n98084), .ZN(
        \DLX_Datapath/RegisterFile/N23278 ) );
  AOI22_X1 U86998 ( .A1(n105621), .A2(n106226), .B1(n106224), .B2(n108692), 
        .ZN(n98084) );
  OAI21_X1 U86999 ( .B1(n106229), .B2(n81498), .A(n98085), .ZN(
        \DLX_Datapath/RegisterFile/N23277 ) );
  AOI22_X1 U87000 ( .A1(n105911), .A2(n106227), .B1(n81291), .B2(n108919), 
        .ZN(n98085) );
  OAI21_X1 U87001 ( .B1(n106269), .B2(n106229), .A(n98086), .ZN(
        \DLX_Datapath/RegisterFile/N23275 ) );
  AOI22_X1 U87002 ( .A1(n106228), .A2(n81265), .B1(n106224), .B2(n107347), 
        .ZN(n98086) );
  AOI21_X1 U87003 ( .B1(n98087), .B2(n94258), .A(n98088), .ZN(n81291) );
  AOI21_X1 U87004 ( .B1(n94999), .B2(n105204), .A(n105601), .ZN(n94258) );
  NOR2_X1 U87005 ( .A1(n98089), .A2(n94999), .ZN(n81290) );
  OR2_X1 U87006 ( .A1(n98088), .A2(n98090), .ZN(n98089) );
  NOR2_X1 U87007 ( .A1(n104504), .A2(n105095), .ZN(n98088) );
  OAI21_X1 U87009 ( .B1(n106149), .B2(n105275), .A(n98093), .ZN(
        \DLX_Datapath/RegisterFile/N23274 ) );
  AOI22_X1 U87010 ( .A1(n98094), .A2(n70372), .B1(n98095), .B2(n94559), .ZN(
        n98093) );
  OAI21_X1 U87011 ( .B1(n105968), .B2(n105275), .A(n98096), .ZN(
        \DLX_Datapath/RegisterFile/N23273 ) );
  AOI22_X1 U87012 ( .A1(n98094), .A2(n70514), .B1(n98095), .B2(n94562), .ZN(
        n98096) );
  OAI21_X1 U87013 ( .B1(n106137), .B2(n105275), .A(n98097), .ZN(
        \DLX_Datapath/RegisterFile/N23272 ) );
  AOI22_X1 U87014 ( .A1(n98094), .A2(n69567), .B1(n98095), .B2(n94564), .ZN(
        n98097) );
  OAI21_X1 U87015 ( .B1(n106210), .B2(n105275), .A(n98098), .ZN(
        \DLX_Datapath/RegisterFile/N23271 ) );
  AOI22_X1 U87016 ( .A1(n98094), .A2(n70228), .B1(n98095), .B2(n94566), .ZN(
        n98098) );
  OAI21_X1 U87017 ( .B1(n106205), .B2(n105275), .A(n98099), .ZN(
        \DLX_Datapath/RegisterFile/N23270 ) );
  AOI22_X1 U87018 ( .A1(n98094), .A2(n110705), .B1(n98095), .B2(n94568), .ZN(
        n98099) );
  OAI21_X1 U87019 ( .B1(n106101), .B2(n105275), .A(n98100), .ZN(
        \DLX_Datapath/RegisterFile/N23269 ) );
  AOI22_X1 U87020 ( .A1(n98094), .A2(n108108), .B1(n98095), .B2(n94570), .ZN(
        n98100) );
  OAI21_X1 U87021 ( .B1(n106256), .B2(n105275), .A(n98101), .ZN(
        \DLX_Datapath/RegisterFile/N23268 ) );
  AOI22_X1 U87022 ( .A1(n98094), .A2(n110807), .B1(n98095), .B2(n94572), .ZN(
        n98101) );
  OAI21_X1 U87023 ( .B1(n105990), .B2(n105275), .A(n98102), .ZN(
        \DLX_Datapath/RegisterFile/N23267 ) );
  AOI22_X1 U87024 ( .A1(n98094), .A2(n110906), .B1(n98095), .B2(n94574), .ZN(
        n98102) );
  OAI21_X1 U87025 ( .B1(n106330), .B2(n105275), .A(n98103), .ZN(
        \DLX_Datapath/RegisterFile/N23266 ) );
  AOI22_X1 U87026 ( .A1(n98094), .A2(n110501), .B1(n98095), .B2(n94576), .ZN(
        n98103) );
  OAI21_X1 U87027 ( .B1(n106192), .B2(n105275), .A(n98104), .ZN(
        \DLX_Datapath/RegisterFile/N23265 ) );
  AOI22_X1 U87028 ( .A1(n98094), .A2(n110284), .B1(n98095), .B2(n94578), .ZN(
        n98104) );
  OAI21_X1 U87029 ( .B1(n106131), .B2(n105275), .A(n98105), .ZN(
        \DLX_Datapath/RegisterFile/N23264 ) );
  AOI22_X1 U87030 ( .A1(n98094), .A2(n110604), .B1(n98095), .B2(n94580), .ZN(
        n98105) );
  OAI21_X1 U87031 ( .B1(n106187), .B2(n105275), .A(n98106), .ZN(
        \DLX_Datapath/RegisterFile/N23263 ) );
  AOI22_X1 U87032 ( .A1(n98094), .A2(n110393), .B1(n98095), .B2(n94582), .ZN(
        n98106) );
  OAI21_X1 U87033 ( .B1(n106165), .B2(n105276), .A(n98107), .ZN(
        \DLX_Datapath/RegisterFile/N23262 ) );
  AOI22_X1 U87034 ( .A1(n98094), .A2(n110071), .B1(n98095), .B2(n94584), .ZN(
        n98107) );
  OAI21_X1 U87035 ( .B1(n106105), .B2(n105276), .A(n98108), .ZN(
        \DLX_Datapath/RegisterFile/N23261 ) );
  AOI22_X1 U87036 ( .A1(n98094), .A2(n110178), .B1(n98095), .B2(n94586), .ZN(
        n98108) );
  OAI21_X1 U87037 ( .B1(n106220), .B2(n105276), .A(n98109), .ZN(
        \DLX_Datapath/RegisterFile/N23260 ) );
  AOI22_X1 U87038 ( .A1(n98094), .A2(n109963), .B1(n98095), .B2(n94588), .ZN(
        n98109) );
  OAI21_X1 U87039 ( .B1(n106111), .B2(n105276), .A(n98110), .ZN(
        \DLX_Datapath/RegisterFile/N23259 ) );
  AOI22_X1 U87040 ( .A1(n98094), .A2(n109846), .B1(n98095), .B2(n94590), .ZN(
        n98110) );
  OAI21_X1 U87041 ( .B1(n106232), .B2(n105276), .A(n98111), .ZN(
        \DLX_Datapath/RegisterFile/N23258 ) );
  AOI22_X1 U87042 ( .A1(n98094), .A2(n108220), .B1(n98095), .B2(n94592), .ZN(
        n98111) );
  OAI21_X1 U87043 ( .B1(n106173), .B2(n105276), .A(n98112), .ZN(
        \DLX_Datapath/RegisterFile/N23257 ) );
  AOI22_X1 U87044 ( .A1(n98094), .A2(n108343), .B1(n98095), .B2(n94594), .ZN(
        n98112) );
  OAI21_X1 U87045 ( .B1(n106238), .B2(n105276), .A(n98113), .ZN(
        \DLX_Datapath/RegisterFile/N23256 ) );
  AOI22_X1 U87046 ( .A1(n98094), .A2(n108454), .B1(n98095), .B2(n94596), .ZN(
        n98113) );
  OAI21_X1 U87047 ( .B1(n81451), .B2(n105276), .A(n98114), .ZN(
        \DLX_Datapath/RegisterFile/N23255 ) );
  AOI22_X1 U87048 ( .A1(n98094), .A2(n107692), .B1(n98095), .B2(n94598), .ZN(
        n98114) );
  OAI21_X1 U87049 ( .B1(n106199), .B2(n105276), .A(n98115), .ZN(
        \DLX_Datapath/RegisterFile/N23254 ) );
  AOI22_X1 U87050 ( .A1(n98094), .A2(n109608), .B1(n98095), .B2(n94600), .ZN(
        n98115) );
  OAI21_X1 U87051 ( .B1(n106246), .B2(n105276), .A(n98116), .ZN(
        \DLX_Datapath/RegisterFile/N23253 ) );
  AOI22_X1 U87052 ( .A1(n98094), .A2(n108570), .B1(n98095), .B2(n94602), .ZN(
        n98116) );
  OAI21_X1 U87053 ( .B1(n106160), .B2(n105276), .A(n98117), .ZN(
        \DLX_Datapath/RegisterFile/N23252 ) );
  AOI22_X1 U87054 ( .A1(n98094), .A2(n109714), .B1(n98095), .B2(n94604), .ZN(
        n98117) );
  OAI21_X1 U87055 ( .B1(n106116), .B2(n105276), .A(n98118), .ZN(
        \DLX_Datapath/RegisterFile/N23251 ) );
  AOI22_X1 U87056 ( .A1(n98094), .A2(n109499), .B1(n98095), .B2(n94606), .ZN(
        n98118) );
  OAI21_X1 U87057 ( .B1(n106011), .B2(n105275), .A(n98119), .ZN(
        \DLX_Datapath/RegisterFile/N23250 ) );
  AOI22_X1 U87058 ( .A1(n98094), .A2(n109036), .B1(n98095), .B2(n94608), .ZN(
        n98119) );
  OAI21_X1 U87059 ( .B1(n106261), .B2(n105276), .A(n98120), .ZN(
        \DLX_Datapath/RegisterFile/N23249 ) );
  AOI22_X1 U87060 ( .A1(n98094), .A2(n109384), .B1(n98095), .B2(n94610), .ZN(
        n98120) );
  OAI21_X1 U87061 ( .B1(n106045), .B2(n105275), .A(n98121), .ZN(
        \DLX_Datapath/RegisterFile/N23248 ) );
  AOI22_X1 U87062 ( .A1(n98094), .A2(n109266), .B1(n98095), .B2(n94612), .ZN(
        n98121) );
  OAI21_X1 U87063 ( .B1(n106051), .B2(n105275), .A(n98122), .ZN(
        \DLX_Datapath/RegisterFile/N23247 ) );
  AOI22_X1 U87064 ( .A1(n98094), .A2(n109157), .B1(n98095), .B2(n94614), .ZN(
        n98122) );
  OAI21_X1 U87065 ( .B1(n106095), .B2(n105276), .A(n98123), .ZN(
        \DLX_Datapath/RegisterFile/N23246 ) );
  AOI22_X1 U87066 ( .A1(n98094), .A2(n108693), .B1(n98095), .B2(n94616), .ZN(
        n98123) );
  OAI21_X1 U87067 ( .B1(n106055), .B2(n105275), .A(n98124), .ZN(
        \DLX_Datapath/RegisterFile/N23245 ) );
  AOI22_X1 U87068 ( .A1(n98094), .A2(n108920), .B1(n98095), .B2(n94618), .ZN(
        n98124) );
  OAI21_X1 U87069 ( .B1(n105216), .B2(n105276), .A(n98125), .ZN(
        \DLX_Datapath/RegisterFile/N23244 ) );
  AOI22_X1 U87070 ( .A1(n98094), .A2(n108808), .B1(n98095), .B2(n94620), .ZN(
        n98125) );
  OAI21_X1 U87071 ( .B1(n81262), .B2(n105276), .A(n98126), .ZN(
        \DLX_Datapath/RegisterFile/N23243 ) );
  AOI22_X1 U87072 ( .A1(n98094), .A2(n107348), .B1(n98095), .B2(n94622), .ZN(
        n98126) );
  AND2_X2 U87073 ( .A1(n98127), .A2(n98128), .ZN(n98095) );
  AND2_X2 U87074 ( .A1(n98129), .A2(n98128), .ZN(n98094) );
  OR2_X1 U87075 ( .A1(n98092), .A2(n105089), .ZN(n98128) );
  NAND2_X1 U87076 ( .A1(n94296), .A2(n104871), .ZN(n98092) );
  OAI21_X1 U87077 ( .B1(n106149), .B2(n98130), .A(n98131), .ZN(
        \DLX_Datapath/RegisterFile/N23242 ) );
  AOI22_X1 U87078 ( .A1(n98132), .A2(n107905), .B1(n98133), .B2(n81521), .ZN(
        n98131) );
  OAI21_X1 U87079 ( .B1(n105968), .B2(n98130), .A(n98134), .ZN(
        \DLX_Datapath/RegisterFile/N23241 ) );
  AOI22_X1 U87080 ( .A1(n98132), .A2(n108001), .B1(n98133), .B2(n81653), .ZN(
        n98134) );
  OAI21_X1 U87081 ( .B1(n106138), .B2(n98130), .A(n98135), .ZN(
        \DLX_Datapath/RegisterFile/N23240 ) );
  AOI22_X1 U87082 ( .A1(n98132), .A2(n107272), .B1(n98133), .B2(n81380), .ZN(
        n98135) );
  OAI21_X1 U87083 ( .B1(n106210), .B2(n98130), .A(n98136), .ZN(
        \DLX_Datapath/RegisterFile/N23239 ) );
  AOI22_X1 U87084 ( .A1(n98132), .A2(n107809), .B1(n98133), .B2(n81377), .ZN(
        n98136) );
  OAI21_X1 U87085 ( .B1(n106205), .B2(n98130), .A(n98137), .ZN(
        \DLX_Datapath/RegisterFile/N23238 ) );
  AOI22_X1 U87086 ( .A1(n98132), .A2(n110706), .B1(n98133), .B2(n81428), .ZN(
        n98137) );
  OAI21_X1 U87087 ( .B1(n106101), .B2(n98130), .A(n98138), .ZN(
        \DLX_Datapath/RegisterFile/N23237 ) );
  AOI22_X1 U87088 ( .A1(n98132), .A2(n108109), .B1(n98133), .B2(n81410), .ZN(
        n98138) );
  OAI21_X1 U87089 ( .B1(n106256), .B2(n105274), .A(n98139), .ZN(
        \DLX_Datapath/RegisterFile/N23236 ) );
  AOI22_X1 U87090 ( .A1(n98132), .A2(n110808), .B1(n98133), .B2(n81700), .ZN(
        n98139) );
  OAI21_X1 U87091 ( .B1(n81629), .B2(n105274), .A(n98140), .ZN(
        \DLX_Datapath/RegisterFile/N23235 ) );
  AOI22_X1 U87092 ( .A1(n98132), .A2(n110907), .B1(n98133), .B2(n81632), .ZN(
        n98140) );
  OAI21_X1 U87093 ( .B1(n106330), .B2(n105274), .A(n98141), .ZN(
        \DLX_Datapath/RegisterFile/N23234 ) );
  AOI22_X1 U87094 ( .A1(n98132), .A2(n110502), .B1(n98133), .B2(n81414), .ZN(
        n98141) );
  OAI21_X1 U87095 ( .B1(n106192), .B2(n105274), .A(n98142), .ZN(
        \DLX_Datapath/RegisterFile/N23233 ) );
  AOI22_X1 U87096 ( .A1(n98132), .A2(n110285), .B1(n98133), .B2(n81317), .ZN(
        n98142) );
  OAI21_X1 U87097 ( .B1(n106131), .B2(n105274), .A(n98143), .ZN(
        \DLX_Datapath/RegisterFile/N23232 ) );
  AOI22_X1 U87098 ( .A1(n98132), .A2(n110605), .B1(n98133), .B2(n81386), .ZN(
        n98143) );
  OAI21_X1 U87099 ( .B1(n106187), .B2(n105274), .A(n98144), .ZN(
        \DLX_Datapath/RegisterFile/N23231 ) );
  AOI22_X1 U87100 ( .A1(n98132), .A2(n110394), .B1(n98133), .B2(n81320), .ZN(
        n98144) );
  OAI21_X1 U87101 ( .B1(n106165), .B2(n105274), .A(n98145), .ZN(
        \DLX_Datapath/RegisterFile/N23230 ) );
  AOI22_X1 U87102 ( .A1(n98132), .A2(n110072), .B1(n98133), .B2(n81604), .ZN(
        n98145) );
  OAI21_X1 U87103 ( .B1(n106106), .B2(n105274), .A(n98146), .ZN(
        \DLX_Datapath/RegisterFile/N23229 ) );
  AOI22_X1 U87104 ( .A1(n98132), .A2(n110179), .B1(n98133), .B2(n81405), .ZN(
        n98146) );
  OAI21_X1 U87105 ( .B1(n106220), .B2(n105274), .A(n98147), .ZN(
        \DLX_Datapath/RegisterFile/N23228 ) );
  AOI22_X1 U87106 ( .A1(n98132), .A2(n109964), .B1(n98133), .B2(n81402), .ZN(
        n98147) );
  OAI21_X1 U87107 ( .B1(n106111), .B2(n105274), .A(n98148), .ZN(
        \DLX_Datapath/RegisterFile/N23227 ) );
  AOI22_X1 U87108 ( .A1(n98132), .A2(n109847), .B1(n98133), .B2(n81400), .ZN(
        n98148) );
  OAI21_X1 U87109 ( .B1(n106233), .B2(n105274), .A(n98149), .ZN(
        \DLX_Datapath/RegisterFile/N23226 ) );
  AOI22_X1 U87110 ( .A1(n98132), .A2(n108221), .B1(n98133), .B2(n81332), .ZN(
        n98149) );
  OAI21_X1 U87111 ( .B1(n106173), .B2(n105274), .A(n98150), .ZN(
        \DLX_Datapath/RegisterFile/N23225 ) );
  AOI22_X1 U87112 ( .A1(n98132), .A2(n108344), .B1(n98133), .B2(n81373), .ZN(
        n98150) );
  OAI21_X1 U87113 ( .B1(n106237), .B2(n105274), .A(n98151), .ZN(
        \DLX_Datapath/RegisterFile/N23224 ) );
  AOI22_X1 U87114 ( .A1(n98132), .A2(n108455), .B1(n98133), .B2(n81322), .ZN(
        n98151) );
  OAI21_X1 U87115 ( .B1(n106071), .B2(n105274), .A(n98152), .ZN(
        \DLX_Datapath/RegisterFile/N23223 ) );
  AOI22_X1 U87116 ( .A1(n98132), .A2(n107693), .B1(n98133), .B2(n81506), .ZN(
        n98152) );
  OAI21_X1 U87117 ( .B1(n106199), .B2(n105274), .A(n98153), .ZN(
        \DLX_Datapath/RegisterFile/N23222 ) );
  AOI22_X1 U87118 ( .A1(n98132), .A2(n109609), .B1(n98133), .B2(n81313), .ZN(
        n98153) );
  OAI21_X1 U87119 ( .B1(n106244), .B2(n105274), .A(n98154), .ZN(
        \DLX_Datapath/RegisterFile/N23221 ) );
  AOI22_X1 U87120 ( .A1(n98132), .A2(n108571), .B1(n98133), .B2(n81330), .ZN(
        n98154) );
  OAI21_X1 U87121 ( .B1(n106160), .B2(n105274), .A(n98155), .ZN(
        \DLX_Datapath/RegisterFile/N23220 ) );
  AOI22_X1 U87122 ( .A1(n98132), .A2(n109715), .B1(n98133), .B2(n81425), .ZN(
        n98155) );
  OAI21_X1 U87123 ( .B1(n106116), .B2(n105274), .A(n98156), .ZN(
        \DLX_Datapath/RegisterFile/N23219 ) );
  AOI22_X1 U87124 ( .A1(n98132), .A2(n109500), .B1(n98133), .B2(n81396), .ZN(
        n98156) );
  OAI21_X1 U87125 ( .B1(n106011), .B2(n105274), .A(n98157), .ZN(
        \DLX_Datapath/RegisterFile/N23218 ) );
  AOI22_X1 U87126 ( .A1(n98132), .A2(n109037), .B1(n98133), .B2(n81590), .ZN(
        n98157) );
  OAI21_X1 U87127 ( .B1(n106262), .B2(n105274), .A(n98158), .ZN(
        \DLX_Datapath/RegisterFile/N23217 ) );
  AOI22_X1 U87128 ( .A1(n98132), .A2(n109385), .B1(n98133), .B2(n81423), .ZN(
        n98158) );
  OAI21_X1 U87129 ( .B1(n106046), .B2(n105274), .A(n98159), .ZN(
        \DLX_Datapath/RegisterFile/N23216 ) );
  AOI22_X1 U87130 ( .A1(n98132), .A2(n109267), .B1(n98133), .B2(n81511), .ZN(
        n98159) );
  OAI21_X1 U87131 ( .B1(n106051), .B2(n105274), .A(n98160), .ZN(
        \DLX_Datapath/RegisterFile/N23215 ) );
  AOI22_X1 U87132 ( .A1(n98132), .A2(n109158), .B1(n98133), .B2(n81503), .ZN(
        n98160) );
  OAI21_X1 U87133 ( .B1(n106096), .B2(n105274), .A(n98161), .ZN(
        \DLX_Datapath/RegisterFile/N23214 ) );
  AOI22_X1 U87134 ( .A1(n98132), .A2(n108694), .B1(n98133), .B2(n81417), .ZN(
        n98161) );
  OAI21_X1 U87135 ( .B1(n106056), .B2(n105274), .A(n98162), .ZN(
        \DLX_Datapath/RegisterFile/N23213 ) );
  AOI22_X1 U87136 ( .A1(n98132), .A2(n108921), .B1(n98133), .B2(n81500), .ZN(
        n98162) );
  OAI21_X1 U87137 ( .B1(n105216), .B2(n105274), .A(n98163), .ZN(
        \DLX_Datapath/RegisterFile/N23212 ) );
  AOI22_X1 U87138 ( .A1(n98132), .A2(n108809), .B1(n98133), .B2(n81335), .ZN(
        n98163) );
  OAI21_X1 U87139 ( .B1(n106269), .B2(n105274), .A(n98164), .ZN(
        \DLX_Datapath/RegisterFile/N23211 ) );
  AOI22_X1 U87140 ( .A1(n98132), .A2(n107349), .B1(n98133), .B2(n81327), .ZN(
        n98164) );
  AND2_X2 U87141 ( .A1(n98127), .A2(n98165), .ZN(n98133) );
  AND2_X2 U87142 ( .A1(n98129), .A2(n98165), .ZN(n98132) );
  OR2_X1 U87143 ( .A1(n98130), .A2(n105089), .ZN(n98165) );
  NAND2_X1 U87144 ( .A1(n94331), .A2(n105124), .ZN(n98130) );
  OAI21_X1 U87145 ( .B1(n106149), .B2(n105273), .A(n98167), .ZN(
        \DLX_Datapath/RegisterFile/N23210 ) );
  AOI22_X1 U87146 ( .A1(n98168), .A2(n94667), .B1(n98169), .B2(n107906), .ZN(
        n98167) );
  OAI21_X1 U87147 ( .B1(n105968), .B2(n105272), .A(n98170), .ZN(
        \DLX_Datapath/RegisterFile/N23209 ) );
  AOI22_X1 U87148 ( .A1(n98168), .A2(n94670), .B1(n98169), .B2(n108002), .ZN(
        n98170) );
  OAI21_X1 U87149 ( .B1(n106138), .B2(n105272), .A(n98171), .ZN(
        \DLX_Datapath/RegisterFile/N23208 ) );
  AOI22_X1 U87150 ( .A1(n98168), .A2(n94672), .B1(n98169), .B2(n107273), .ZN(
        n98171) );
  OAI21_X1 U87151 ( .B1(n106211), .B2(n105272), .A(n98172), .ZN(
        \DLX_Datapath/RegisterFile/N23207 ) );
  AOI22_X1 U87152 ( .A1(n98168), .A2(n94674), .B1(n98169), .B2(n107810), .ZN(
        n98172) );
  OAI21_X1 U87153 ( .B1(n106205), .B2(n105273), .A(n98173), .ZN(
        \DLX_Datapath/RegisterFile/N23206 ) );
  AOI22_X1 U87154 ( .A1(n98168), .A2(n94676), .B1(n98169), .B2(n110707), .ZN(
        n98173) );
  OAI21_X1 U87155 ( .B1(n106101), .B2(n105272), .A(n98174), .ZN(
        \DLX_Datapath/RegisterFile/N23205 ) );
  AOI22_X1 U87156 ( .A1(n98168), .A2(n94678), .B1(n98169), .B2(n108110), .ZN(
        n98174) );
  OAI21_X1 U87157 ( .B1(n106257), .B2(n105272), .A(n98175), .ZN(
        \DLX_Datapath/RegisterFile/N23204 ) );
  AOI22_X1 U87158 ( .A1(n98168), .A2(n94680), .B1(n98169), .B2(n110809), .ZN(
        n98175) );
  AOI22_X1 U87160 ( .A1(n98168), .A2(n94682), .B1(n98169), .B2(n110908), .ZN(
        n98176) );
  OAI21_X1 U87161 ( .B1(n106330), .B2(n105273), .A(n98177), .ZN(
        \DLX_Datapath/RegisterFile/N23202 ) );
  AOI22_X1 U87162 ( .A1(n98168), .A2(n94684), .B1(n98169), .B2(n110503), .ZN(
        n98177) );
  OAI21_X1 U87163 ( .B1(n106193), .B2(n105272), .A(n98178), .ZN(
        \DLX_Datapath/RegisterFile/N23201 ) );
  AOI22_X1 U87164 ( .A1(n98168), .A2(n94686), .B1(n98169), .B2(n110286), .ZN(
        n98178) );
  OAI21_X1 U87165 ( .B1(n106131), .B2(n105273), .A(n98179), .ZN(
        \DLX_Datapath/RegisterFile/N23200 ) );
  AOI22_X1 U87166 ( .A1(n98168), .A2(n94688), .B1(n98169), .B2(n110606), .ZN(
        n98179) );
  OAI21_X1 U87167 ( .B1(n106187), .B2(n105272), .A(n98180), .ZN(
        \DLX_Datapath/RegisterFile/N23199 ) );
  AOI22_X1 U87168 ( .A1(n98168), .A2(n94690), .B1(n98169), .B2(n110395), .ZN(
        n98180) );
  OAI21_X1 U87169 ( .B1(n106165), .B2(n105272), .A(n98181), .ZN(
        \DLX_Datapath/RegisterFile/N23198 ) );
  AOI22_X1 U87170 ( .A1(n98168), .A2(n94692), .B1(n98169), .B2(n110073), .ZN(
        n98181) );
  OAI21_X1 U87171 ( .B1(n106106), .B2(n105272), .A(n98182), .ZN(
        \DLX_Datapath/RegisterFile/N23197 ) );
  AOI22_X1 U87172 ( .A1(n98168), .A2(n94694), .B1(n98169), .B2(n110180), .ZN(
        n98182) );
  OAI21_X1 U87173 ( .B1(n106221), .B2(n105272), .A(n98183), .ZN(
        \DLX_Datapath/RegisterFile/N23196 ) );
  AOI22_X1 U87174 ( .A1(n98168), .A2(n94696), .B1(n98169), .B2(n109965), .ZN(
        n98183) );
  OAI21_X1 U87175 ( .B1(n106111), .B2(n105272), .A(n98184), .ZN(
        \DLX_Datapath/RegisterFile/N23195 ) );
  AOI22_X1 U87176 ( .A1(n98168), .A2(n94698), .B1(n98169), .B2(n109848), .ZN(
        n98184) );
  OAI21_X1 U87177 ( .B1(n106232), .B2(n105272), .A(n98185), .ZN(
        \DLX_Datapath/RegisterFile/N23194 ) );
  AOI22_X1 U87178 ( .A1(n98168), .A2(n94700), .B1(n98169), .B2(n108222), .ZN(
        n98185) );
  OAI21_X1 U87179 ( .B1(n106173), .B2(n105272), .A(n98186), .ZN(
        \DLX_Datapath/RegisterFile/N23193 ) );
  AOI22_X1 U87180 ( .A1(n98168), .A2(n94702), .B1(n98169), .B2(n108345), .ZN(
        n98186) );
  OAI21_X1 U87181 ( .B1(n106238), .B2(n105272), .A(n98187), .ZN(
        \DLX_Datapath/RegisterFile/N23192 ) );
  AOI22_X1 U87182 ( .A1(n98168), .A2(n94704), .B1(n98169), .B2(n108456), .ZN(
        n98187) );
  OAI21_X1 U87183 ( .B1(n81451), .B2(n105272), .A(n98188), .ZN(
        \DLX_Datapath/RegisterFile/N23191 ) );
  AOI22_X1 U87184 ( .A1(n98168), .A2(n94706), .B1(n98169), .B2(n107694), .ZN(
        n98188) );
  OAI21_X1 U87185 ( .B1(n106200), .B2(n105272), .A(n98189), .ZN(
        \DLX_Datapath/RegisterFile/N23190 ) );
  AOI22_X1 U87186 ( .A1(n98168), .A2(n94708), .B1(n98169), .B2(n109610), .ZN(
        n98189) );
  OAI21_X1 U87187 ( .B1(n106246), .B2(n105272), .A(n98190), .ZN(
        \DLX_Datapath/RegisterFile/N23189 ) );
  AOI22_X1 U87188 ( .A1(n98168), .A2(n94710), .B1(n98169), .B2(n108572), .ZN(
        n98190) );
  OAI21_X1 U87189 ( .B1(n106160), .B2(n105272), .A(n98191), .ZN(
        \DLX_Datapath/RegisterFile/N23188 ) );
  AOI22_X1 U87190 ( .A1(n98168), .A2(n94712), .B1(n98169), .B2(n109716), .ZN(
        n98191) );
  OAI21_X1 U87191 ( .B1(n106116), .B2(n105272), .A(n98192), .ZN(
        \DLX_Datapath/RegisterFile/N23187 ) );
  AOI22_X1 U87192 ( .A1(n98168), .A2(n94714), .B1(n98169), .B2(n109501), .ZN(
        n98192) );
  OAI21_X1 U87193 ( .B1(n106011), .B2(n105273), .A(n98193), .ZN(
        \DLX_Datapath/RegisterFile/N23186 ) );
  AOI22_X1 U87194 ( .A1(n98168), .A2(n81259), .B1(n98169), .B2(n109038), .ZN(
        n98193) );
  OAI21_X1 U87195 ( .B1(n106261), .B2(n105273), .A(n98194), .ZN(
        \DLX_Datapath/RegisterFile/N23185 ) );
  AOI22_X1 U87196 ( .A1(n98168), .A2(n94717), .B1(n98169), .B2(n109386), .ZN(
        n98194) );
  OAI21_X1 U87197 ( .B1(n106046), .B2(n105273), .A(n98195), .ZN(
        \DLX_Datapath/RegisterFile/N23184 ) );
  AOI22_X1 U87198 ( .A1(n98168), .A2(n94719), .B1(n98169), .B2(n109268), .ZN(
        n98195) );
  OAI21_X1 U87199 ( .B1(n106051), .B2(n105273), .A(n98196), .ZN(
        \DLX_Datapath/RegisterFile/N23183 ) );
  AOI22_X1 U87200 ( .A1(n98168), .A2(n94721), .B1(n98169), .B2(n109159), .ZN(
        n98196) );
  OAI21_X1 U87201 ( .B1(n106096), .B2(n105273), .A(n98197), .ZN(
        \DLX_Datapath/RegisterFile/N23182 ) );
  AOI22_X1 U87202 ( .A1(n98168), .A2(n94723), .B1(n98169), .B2(n108695), .ZN(
        n98197) );
  OAI21_X1 U87203 ( .B1(n106056), .B2(n105273), .A(n98198), .ZN(
        \DLX_Datapath/RegisterFile/N23181 ) );
  AOI22_X1 U87204 ( .A1(n98168), .A2(n94725), .B1(n98169), .B2(n108922), .ZN(
        n98198) );
  OAI21_X1 U87205 ( .B1(n105216), .B2(n105273), .A(n98199), .ZN(
        \DLX_Datapath/RegisterFile/N23180 ) );
  AOI22_X1 U87206 ( .A1(n98168), .A2(n94727), .B1(n98169), .B2(n108810), .ZN(
        n98199) );
  OAI21_X1 U87207 ( .B1(n106268), .B2(n105273), .A(n98200), .ZN(
        \DLX_Datapath/RegisterFile/N23179 ) );
  AOI22_X1 U87208 ( .A1(n98168), .A2(n94729), .B1(n98169), .B2(n107350), .ZN(
        n98200) );
  AND2_X2 U87209 ( .A1(n98129), .A2(n98201), .ZN(n98169) );
  OAI21_X1 U87210 ( .B1(n94366), .B2(n98127), .A(n105602), .ZN(n98129) );
  AND2_X2 U87211 ( .A1(n98127), .A2(n98201), .ZN(n98168) );
  OR2_X1 U87212 ( .A1(n98166), .A2(n105091), .ZN(n98201) );
  NOR2_X1 U87213 ( .A1(n94999), .A2(n98090), .ZN(n98127) );
  NAND2_X1 U87214 ( .A1(n94367), .A2(n104871), .ZN(n98166) );
  OAI21_X1 U87215 ( .B1(n106223), .B2(n81358), .A(n98202), .ZN(
        \DLX_Datapath/RegisterFile/N23178 ) );
  AOI22_X1 U87216 ( .A1(n106216), .A2(n107907), .B1(n81360), .B2(n106213), 
        .ZN(n98202) );
  OAI21_X1 U87217 ( .B1(n106223), .B2(n105969), .A(n98203), .ZN(
        \DLX_Datapath/RegisterFile/N23177 ) );
  AOI22_X1 U87218 ( .A1(n106216), .A2(n108003), .B1(n94511), .B2(n106214), 
        .ZN(n98203) );
  OAI21_X1 U87219 ( .B1(n106223), .B2(n106138), .A(n98204), .ZN(
        \DLX_Datapath/RegisterFile/N23176 ) );
  AOI22_X1 U87220 ( .A1(n106216), .A2(n107274), .B1(n81539), .B2(n106213), 
        .ZN(n98204) );
  OAI21_X1 U87221 ( .B1(n106223), .B2(n106204), .A(n98205), .ZN(
        \DLX_Datapath/RegisterFile/N23174 ) );
  AOI22_X1 U87222 ( .A1(n74077), .A2(n106216), .B1(n81308), .B2(n106215), .ZN(
        n98205) );
  OAI21_X1 U87223 ( .B1(n106223), .B2(n106100), .A(n98206), .ZN(
        \DLX_Datapath/RegisterFile/N23173 ) );
  AOI22_X1 U87224 ( .A1(n70664), .A2(n106216), .B1(n94516), .B2(n106213), .ZN(
        n98206) );
  OAI21_X1 U87225 ( .B1(n106256), .B2(n106223), .A(n98207), .ZN(
        \DLX_Datapath/RegisterFile/N23172 ) );
  AOI22_X1 U87226 ( .A1(n74218), .A2(n106216), .B1(n106215), .B2(n81272), .ZN(
        n98207) );
  OAI21_X1 U87227 ( .B1(n106223), .B2(n105992), .A(n98208), .ZN(
        \DLX_Datapath/RegisterFile/N23171 ) );
  AOI22_X1 U87228 ( .A1(n106216), .A2(n110909), .B1(n94519), .B2(n106215), 
        .ZN(n98208) );
  OAI21_X1 U87229 ( .B1(n106330), .B2(n106223), .A(n98209), .ZN(
        \DLX_Datapath/RegisterFile/N23170 ) );
  AOI22_X1 U87230 ( .A1(n106216), .A2(n110504), .B1(n106214), .B2(n80192), 
        .ZN(n98209) );
  OAI21_X1 U87231 ( .B1(n106223), .B2(n106192), .A(n98210), .ZN(
        \DLX_Datapath/RegisterFile/N23169 ) );
  AOI22_X1 U87232 ( .A1(n106217), .A2(n110287), .B1(n81474), .B2(n106214), 
        .ZN(n98210) );
  OAI21_X1 U87233 ( .B1(n106223), .B2(n81383), .A(n98211), .ZN(
        \DLX_Datapath/RegisterFile/N23168 ) );
  AOI22_X1 U87234 ( .A1(n106217), .A2(n110607), .B1(n94523), .B2(n106213), 
        .ZN(n98211) );
  OAI21_X1 U87235 ( .B1(n106223), .B2(n106187), .A(n98212), .ZN(
        \DLX_Datapath/RegisterFile/N23167 ) );
  AOI22_X1 U87236 ( .A1(n106217), .A2(n110396), .B1(n106062), .B2(n106215), 
        .ZN(n98212) );
  OAI21_X1 U87237 ( .B1(n106223), .B2(n81345), .A(n98213), .ZN(
        \DLX_Datapath/RegisterFile/N23166 ) );
  AOI22_X1 U87238 ( .A1(n106217), .A2(n110074), .B1(n81347), .B2(n106213), 
        .ZN(n98213) );
  OAI21_X1 U87239 ( .B1(n106223), .B2(n81403), .A(n98214), .ZN(
        \DLX_Datapath/RegisterFile/N23165 ) );
  AOI22_X1 U87240 ( .A1(n106217), .A2(n110181), .B1(n94527), .B2(n106213), 
        .ZN(n98214) );
  OAI21_X1 U87241 ( .B1(n106223), .B2(n106109), .A(n98215), .ZN(
        \DLX_Datapath/RegisterFile/N23163 ) );
  AOI22_X1 U87242 ( .A1(n106217), .A2(n109849), .B1(n94530), .B2(n106213), 
        .ZN(n98215) );
  OAI21_X1 U87243 ( .B1(n106233), .B2(n106223), .A(n98216), .ZN(
        \DLX_Datapath/RegisterFile/N23162 ) );
  AOI22_X1 U87244 ( .A1(n106217), .A2(n108223), .B1(n106214), .B2(n81286), 
        .ZN(n98216) );
  OAI21_X1 U87245 ( .B1(n106223), .B2(n81340), .A(n98217), .ZN(
        \DLX_Datapath/RegisterFile/N23161 ) );
  AOI22_X1 U87246 ( .A1(n106217), .A2(n108346), .B1(n106169), .B2(n106213), 
        .ZN(n98217) );
  OAI21_X1 U87247 ( .B1(n106238), .B2(n106223), .A(n98218), .ZN(
        \DLX_Datapath/RegisterFile/N23160 ) );
  AOI22_X1 U87248 ( .A1(n106217), .A2(n108457), .B1(n106215), .B2(n81283), 
        .ZN(n98218) );
  OAI21_X1 U87249 ( .B1(n106223), .B2(n106071), .A(n98219), .ZN(
        \DLX_Datapath/RegisterFile/N23159 ) );
  AOI22_X1 U87250 ( .A1(n106217), .A2(n107695), .B1(n81453), .B2(n106215), 
        .ZN(n98219) );
  OAI21_X1 U87251 ( .B1(n106223), .B2(n106199), .A(n98220), .ZN(
        \DLX_Datapath/RegisterFile/N23158 ) );
  AOI22_X1 U87252 ( .A1(n72607), .A2(n106216), .B1(n94536), .B2(n106213), .ZN(
        n98220) );
  OAI21_X1 U87253 ( .B1(n106246), .B2(n106223), .A(n98221), .ZN(
        \DLX_Datapath/RegisterFile/N23157 ) );
  AOI22_X1 U87254 ( .A1(n71266), .A2(n106216), .B1(n106214), .B2(n106241), 
        .ZN(n98221) );
  OAI21_X1 U87255 ( .B1(n106223), .B2(n81349), .A(n98222), .ZN(
        \DLX_Datapath/RegisterFile/N23156 ) );
  AOI22_X1 U87256 ( .A1(n106217), .A2(n109717), .B1(n81351), .B2(n106213), 
        .ZN(n98222) );
  AOI22_X1 U87258 ( .A1(n81296), .A2(n109502), .B1(n106021), .B2(n106215), 
        .ZN(n98223) );
  OAI21_X1 U87259 ( .B1(n106011), .B2(n106223), .A(n98224), .ZN(
        \DLX_Datapath/RegisterFile/N23154 ) );
  AOI22_X1 U87260 ( .A1(n81296), .A2(n109039), .B1(n94541), .B2(n106214), .ZN(
        n98224) );
  OAI21_X1 U87261 ( .B1(n106262), .B2(n106223), .A(n98225), .ZN(
        \DLX_Datapath/RegisterFile/N23153 ) );
  AOI22_X1 U87262 ( .A1(n81296), .A2(n109387), .B1(n106214), .B2(n81269), .ZN(
        n98225) );
  OAI21_X1 U87263 ( .B1(n106223), .B2(n81509), .A(n98226), .ZN(
        \DLX_Datapath/RegisterFile/N23152 ) );
  AOI22_X1 U87264 ( .A1(n81296), .A2(n109269), .B1(n105625), .B2(n106214), 
        .ZN(n98226) );
  OAI21_X1 U87265 ( .B1(n106223), .B2(n81501), .A(n98227), .ZN(
        \DLX_Datapath/RegisterFile/N23151 ) );
  AOI22_X1 U87266 ( .A1(n106216), .A2(n109160), .B1(n94546), .B2(n106215), 
        .ZN(n98227) );
  OAI21_X1 U87267 ( .B1(n106223), .B2(n106095), .A(n98228), .ZN(
        \DLX_Datapath/RegisterFile/N23150 ) );
  AOI22_X1 U87268 ( .A1(n81296), .A2(n108696), .B1(n94548), .B2(n106214), .ZN(
        n98228) );
  OAI21_X1 U87269 ( .B1(n106223), .B2(n106053), .A(n98229), .ZN(
        \DLX_Datapath/RegisterFile/N23149 ) );
  AOI22_X1 U87270 ( .A1(n81296), .A2(n108923), .B1(n81783), .B2(n106215), .ZN(
        n98229) );
  OAI21_X1 U87271 ( .B1(n105216), .B2(n106223), .A(n98230), .ZN(
        \DLX_Datapath/RegisterFile/N23148 ) );
  AOI22_X1 U87272 ( .A1(n81296), .A2(n108811), .B1(n106215), .B2(n80188), .ZN(
        n98230) );
  OAI21_X1 U87273 ( .B1(n81262), .B2(n106223), .A(n98231), .ZN(
        \DLX_Datapath/RegisterFile/N23147 ) );
  AOI22_X1 U87274 ( .A1(n106216), .A2(n107351), .B1(n106215), .B2(n81265), 
        .ZN(n98231) );
  OR2_X1 U87276 ( .A1(n98233), .A2(n95131), .ZN(n98232) );
  AOI21_X1 U87277 ( .B1(n98087), .B2(n94398), .A(n104779), .ZN(n81296) );
  NOR2_X1 U87278 ( .A1(n81293), .A2(n105094), .ZN(n98233) );
  AOI21_X1 U87279 ( .B1(n95131), .B2(n105204), .A(n105601), .ZN(n94398) );
  NAND2_X1 U87280 ( .A1(n104871), .A2(n94399), .ZN(n81293) );
  OAI21_X1 U87281 ( .B1(n106149), .B2(n98234), .A(n98235), .ZN(
        \DLX_Datapath/RegisterFile/N23146 ) );
  AOI22_X1 U87282 ( .A1(n98236), .A2(n94559), .B1(n98237), .B2(n70376), .ZN(
        n98235) );
  OAI21_X1 U87283 ( .B1(n105968), .B2(n98234), .A(n98238), .ZN(
        \DLX_Datapath/RegisterFile/N23145 ) );
  AOI22_X1 U87284 ( .A1(n98236), .A2(n94562), .B1(n98237), .B2(n70518), .ZN(
        n98238) );
  OAI21_X1 U87285 ( .B1(n106138), .B2(n98234), .A(n98239), .ZN(
        \DLX_Datapath/RegisterFile/N23144 ) );
  AOI22_X1 U87286 ( .A1(n98236), .A2(n94564), .B1(n98237), .B2(n69571), .ZN(
        n98239) );
  OAI21_X1 U87287 ( .B1(n106210), .B2(n98234), .A(n98240), .ZN(
        \DLX_Datapath/RegisterFile/N23143 ) );
  AOI22_X1 U87288 ( .A1(n98236), .A2(n94566), .B1(n98237), .B2(n107812), .ZN(
        n98240) );
  OAI21_X1 U87289 ( .B1(n106205), .B2(n98234), .A(n98241), .ZN(
        \DLX_Datapath/RegisterFile/N23142 ) );
  AOI22_X1 U87290 ( .A1(n98236), .A2(n94568), .B1(n98237), .B2(n110708), .ZN(
        n98241) );
  OAI21_X1 U87291 ( .B1(n106101), .B2(n98234), .A(n98242), .ZN(
        \DLX_Datapath/RegisterFile/N23141 ) );
  AOI22_X1 U87292 ( .A1(n98236), .A2(n94570), .B1(n98237), .B2(n108111), .ZN(
        n98242) );
  OAI21_X1 U87293 ( .B1(n106257), .B2(n105271), .A(n98243), .ZN(
        \DLX_Datapath/RegisterFile/N23140 ) );
  AOI22_X1 U87294 ( .A1(n98236), .A2(n94572), .B1(n98237), .B2(n110810), .ZN(
        n98243) );
  OAI21_X1 U87295 ( .B1(n81629), .B2(n105271), .A(n98244), .ZN(
        \DLX_Datapath/RegisterFile/N23139 ) );
  AOI22_X1 U87296 ( .A1(n98236), .A2(n94574), .B1(n98237), .B2(n110910), .ZN(
        n98244) );
  OAI21_X1 U87297 ( .B1(n106330), .B2(n105271), .A(n98245), .ZN(
        \DLX_Datapath/RegisterFile/N23138 ) );
  AOI22_X1 U87298 ( .A1(n98236), .A2(n94576), .B1(n98237), .B2(n110505), .ZN(
        n98245) );
  OAI21_X1 U87299 ( .B1(n106193), .B2(n105271), .A(n98246), .ZN(
        \DLX_Datapath/RegisterFile/N23137 ) );
  AOI22_X1 U87300 ( .A1(n98236), .A2(n94578), .B1(n98237), .B2(n110288), .ZN(
        n98246) );
  OAI21_X1 U87301 ( .B1(n106131), .B2(n105271), .A(n98247), .ZN(
        \DLX_Datapath/RegisterFile/N23136 ) );
  AOI22_X1 U87302 ( .A1(n98236), .A2(n94580), .B1(n98237), .B2(n110608), .ZN(
        n98247) );
  OAI21_X1 U87303 ( .B1(n106188), .B2(n105271), .A(n98248), .ZN(
        \DLX_Datapath/RegisterFile/N23135 ) );
  AOI22_X1 U87304 ( .A1(n98236), .A2(n94582), .B1(n98237), .B2(n110397), .ZN(
        n98248) );
  OAI21_X1 U87305 ( .B1(n106165), .B2(n105271), .A(n98249), .ZN(
        \DLX_Datapath/RegisterFile/N23134 ) );
  AOI22_X1 U87306 ( .A1(n98236), .A2(n94584), .B1(n98237), .B2(n110075), .ZN(
        n98249) );
  OAI21_X1 U87307 ( .B1(n106106), .B2(n105271), .A(n98250), .ZN(
        \DLX_Datapath/RegisterFile/N23133 ) );
  AOI22_X1 U87308 ( .A1(n98236), .A2(n94586), .B1(n98237), .B2(n110182), .ZN(
        n98250) );
  OAI21_X1 U87309 ( .B1(n106220), .B2(n105271), .A(n98251), .ZN(
        \DLX_Datapath/RegisterFile/N23132 ) );
  AOI22_X1 U87310 ( .A1(n98236), .A2(n94588), .B1(n98237), .B2(n109967), .ZN(
        n98251) );
  OAI21_X1 U87311 ( .B1(n106111), .B2(n105271), .A(n98252), .ZN(
        \DLX_Datapath/RegisterFile/N23131 ) );
  AOI22_X1 U87312 ( .A1(n98236), .A2(n94590), .B1(n98237), .B2(n109850), .ZN(
        n98252) );
  OAI21_X1 U87313 ( .B1(n106233), .B2(n105271), .A(n98253), .ZN(
        \DLX_Datapath/RegisterFile/N23130 ) );
  AOI22_X1 U87314 ( .A1(n98236), .A2(n94592), .B1(n98237), .B2(n108224), .ZN(
        n98253) );
  OAI21_X1 U87315 ( .B1(n106173), .B2(n105271), .A(n98254), .ZN(
        \DLX_Datapath/RegisterFile/N23129 ) );
  AOI22_X1 U87316 ( .A1(n98236), .A2(n94594), .B1(n98237), .B2(n108347), .ZN(
        n98254) );
  OAI21_X1 U87317 ( .B1(n106238), .B2(n105271), .A(n98255), .ZN(
        \DLX_Datapath/RegisterFile/N23128 ) );
  AOI22_X1 U87318 ( .A1(n98236), .A2(n94596), .B1(n98237), .B2(n108458), .ZN(
        n98255) );
  OAI21_X1 U87319 ( .B1(n106072), .B2(n105271), .A(n98256), .ZN(
        \DLX_Datapath/RegisterFile/N23127 ) );
  AOI22_X1 U87320 ( .A1(n98236), .A2(n94598), .B1(n98237), .B2(n107696), .ZN(
        n98256) );
  OAI21_X1 U87321 ( .B1(n106200), .B2(n105271), .A(n98257), .ZN(
        \DLX_Datapath/RegisterFile/N23126 ) );
  AOI22_X1 U87322 ( .A1(n98236), .A2(n94600), .B1(n98237), .B2(n109611), .ZN(
        n98257) );
  OAI21_X1 U87323 ( .B1(n106243), .B2(n105271), .A(n98258), .ZN(
        \DLX_Datapath/RegisterFile/N23125 ) );
  AOI22_X1 U87324 ( .A1(n98236), .A2(n94602), .B1(n98237), .B2(n108573), .ZN(
        n98258) );
  OAI21_X1 U87325 ( .B1(n106160), .B2(n105271), .A(n98259), .ZN(
        \DLX_Datapath/RegisterFile/N23124 ) );
  AOI22_X1 U87326 ( .A1(n98236), .A2(n94604), .B1(n98237), .B2(n109718), .ZN(
        n98259) );
  OAI21_X1 U87327 ( .B1(n106116), .B2(n105271), .A(n98260), .ZN(
        \DLX_Datapath/RegisterFile/N23123 ) );
  AOI22_X1 U87328 ( .A1(n98236), .A2(n94606), .B1(n98237), .B2(n109503), .ZN(
        n98260) );
  OAI21_X1 U87329 ( .B1(n106007), .B2(n105271), .A(n98261), .ZN(
        \DLX_Datapath/RegisterFile/N23122 ) );
  AOI22_X1 U87330 ( .A1(n98236), .A2(n94608), .B1(n98237), .B2(n109040), .ZN(
        n98261) );
  OAI21_X1 U87331 ( .B1(n106262), .B2(n105271), .A(n98262), .ZN(
        \DLX_Datapath/RegisterFile/N23121 ) );
  AOI22_X1 U87332 ( .A1(n98236), .A2(n94610), .B1(n98237), .B2(n109388), .ZN(
        n98262) );
  OAI21_X1 U87333 ( .B1(n106046), .B2(n105271), .A(n98263), .ZN(
        \DLX_Datapath/RegisterFile/N23120 ) );
  AOI22_X1 U87334 ( .A1(n98236), .A2(n94612), .B1(n98237), .B2(n109270), .ZN(
        n98263) );
  OAI21_X1 U87335 ( .B1(n106050), .B2(n105271), .A(n98264), .ZN(
        \DLX_Datapath/RegisterFile/N23119 ) );
  AOI22_X1 U87336 ( .A1(n98236), .A2(n94614), .B1(n98237), .B2(n109161), .ZN(
        n98264) );
  OAI21_X1 U87337 ( .B1(n106096), .B2(n105271), .A(n98265), .ZN(
        \DLX_Datapath/RegisterFile/N23118 ) );
  AOI22_X1 U87338 ( .A1(n98236), .A2(n94616), .B1(n98237), .B2(n108697), .ZN(
        n98265) );
  OAI21_X1 U87339 ( .B1(n106056), .B2(n105271), .A(n98266), .ZN(
        \DLX_Datapath/RegisterFile/N23117 ) );
  AOI22_X1 U87340 ( .A1(n98236), .A2(n94618), .B1(n98237), .B2(n108924), .ZN(
        n98266) );
  OAI21_X1 U87341 ( .B1(n105216), .B2(n105271), .A(n98267), .ZN(
        \DLX_Datapath/RegisterFile/N23116 ) );
  AOI22_X1 U87342 ( .A1(n98236), .A2(n94620), .B1(n98237), .B2(n108812), .ZN(
        n98267) );
  OAI21_X1 U87343 ( .B1(n81262), .B2(n105271), .A(n98268), .ZN(
        \DLX_Datapath/RegisterFile/N23115 ) );
  AOI22_X1 U87344 ( .A1(n98236), .A2(n94622), .B1(n98237), .B2(n107352), .ZN(
        n98268) );
  AND2_X2 U87345 ( .A1(n98269), .A2(n98270), .ZN(n98237) );
  AND2_X2 U87346 ( .A1(n98271), .A2(n98270), .ZN(n98236) );
  OR2_X1 U87347 ( .A1(n98234), .A2(n105089), .ZN(n98270) );
  NAND2_X1 U87348 ( .A1(n94434), .A2(n105124), .ZN(n98234) );
  OAI21_X1 U87349 ( .B1(n106202), .B2(n81358), .A(n98272), .ZN(
        \DLX_Datapath/RegisterFile/N23114 ) );
  AOI22_X1 U87350 ( .A1(n81521), .A2(n106196), .B1(n81314), .B2(n107908), .ZN(
        n98272) );
  OAI21_X1 U87351 ( .B1(n106202), .B2(n81651), .A(n98273), .ZN(
        \DLX_Datapath/RegisterFile/N23113 ) );
  AOI22_X1 U87352 ( .A1(n81653), .A2(n106195), .B1(n81314), .B2(n108004), .ZN(
        n98273) );
  OAI21_X1 U87353 ( .B1(n106202), .B2(n106136), .A(n98274), .ZN(
        \DLX_Datapath/RegisterFile/N23112 ) );
  AOI22_X1 U87354 ( .A1(n81380), .A2(n106196), .B1(n81314), .B2(n107275), .ZN(
        n98274) );
  OAI21_X1 U87355 ( .B1(n106211), .B2(n106202), .A(n98275), .ZN(
        \DLX_Datapath/RegisterFile/N23111 ) );
  AOI22_X1 U87356 ( .A1(n81377), .A2(n106195), .B1(n81314), .B2(n107813), .ZN(
        n98275) );
  OAI21_X1 U87357 ( .B1(n106206), .B2(n106202), .A(n98276), .ZN(
        \DLX_Datapath/RegisterFile/N23110 ) );
  AOI22_X1 U87358 ( .A1(n81428), .A2(n81312), .B1(n81314), .B2(n110709), .ZN(
        n98276) );
  OAI21_X1 U87359 ( .B1(n106202), .B2(n81408), .A(n98277), .ZN(
        \DLX_Datapath/RegisterFile/N23109 ) );
  AOI22_X1 U87360 ( .A1(n81410), .A2(n106195), .B1(n81314), .B2(n108112), .ZN(
        n98277) );
  OAI21_X1 U87361 ( .B1(n106257), .B2(n106202), .A(n98278), .ZN(
        \DLX_Datapath/RegisterFile/N23108 ) );
  AOI22_X1 U87362 ( .A1(n81700), .A2(n106196), .B1(n81314), .B2(n110811), .ZN(
        n98278) );
  OAI21_X1 U87363 ( .B1(n106202), .B2(n105991), .A(n98279), .ZN(
        \DLX_Datapath/RegisterFile/N23107 ) );
  AOI22_X1 U87364 ( .A1(n81632), .A2(n106196), .B1(n81314), .B2(n110911), .ZN(
        n98279) );
  OAI21_X1 U87365 ( .B1(n106330), .B2(n106202), .A(n98280), .ZN(
        \DLX_Datapath/RegisterFile/N23106 ) );
  AOI22_X1 U87366 ( .A1(n81414), .A2(n106195), .B1(n81314), .B2(n110506), .ZN(
        n98280) );
  OAI21_X1 U87367 ( .B1(n106202), .B2(n106130), .A(n98281), .ZN(
        \DLX_Datapath/RegisterFile/N23104 ) );
  AOI22_X1 U87368 ( .A1(n81386), .A2(n81312), .B1(n81314), .B2(n110609), .ZN(
        n98281) );
  OAI21_X1 U87369 ( .B1(n106202), .B2(n106163), .A(n98282), .ZN(
        \DLX_Datapath/RegisterFile/N23102 ) );
  AOI22_X1 U87370 ( .A1(n81604), .A2(n106195), .B1(n81314), .B2(n110076), .ZN(
        n98282) );
  OAI21_X1 U87371 ( .B1(n106202), .B2(n106104), .A(n98283), .ZN(
        \DLX_Datapath/RegisterFile/N23101 ) );
  AOI22_X1 U87372 ( .A1(n81405), .A2(n81312), .B1(n81314), .B2(n110183), .ZN(
        n98283) );
  OAI21_X1 U87373 ( .B1(n106221), .B2(n106202), .A(n98284), .ZN(
        \DLX_Datapath/RegisterFile/N23100 ) );
  AOI22_X1 U87374 ( .A1(n81402), .A2(n106196), .B1(n81314), .B2(n109968), .ZN(
        n98284) );
  OAI21_X1 U87375 ( .B1(n106202), .B2(n106111), .A(n98285), .ZN(
        \DLX_Datapath/RegisterFile/N23099 ) );
  AOI22_X1 U87376 ( .A1(n81400), .A2(n106196), .B1(n81314), .B2(n109851), .ZN(
        n98285) );
  OAI21_X1 U87377 ( .B1(n106233), .B2(n106202), .A(n98286), .ZN(
        \DLX_Datapath/RegisterFile/N23098 ) );
  AOI22_X1 U87378 ( .A1(n81332), .A2(n106195), .B1(n81314), .B2(n108225), .ZN(
        n98286) );
  OAI21_X1 U87379 ( .B1(n106202), .B2(n106170), .A(n98287), .ZN(
        \DLX_Datapath/RegisterFile/N23097 ) );
  AOI22_X1 U87380 ( .A1(n81373), .A2(n106195), .B1(n81314), .B2(n108348), .ZN(
        n98287) );
  OAI21_X1 U87381 ( .B1(n106202), .B2(n106069), .A(n98288), .ZN(
        \DLX_Datapath/RegisterFile/N23095 ) );
  AOI22_X1 U87382 ( .A1(n81506), .A2(n81312), .B1(n81314), .B2(n107697), .ZN(
        n98288) );
  OAI21_X1 U87383 ( .B1(n106244), .B2(n106202), .A(n98289), .ZN(
        \DLX_Datapath/RegisterFile/N23093 ) );
  AOI22_X1 U87384 ( .A1(n81330), .A2(n106196), .B1(n81314), .B2(n108574), .ZN(
        n98289) );
  OAI21_X1 U87385 ( .B1(n106202), .B2(n106157), .A(n98290), .ZN(
        \DLX_Datapath/RegisterFile/N23092 ) );
  AOI22_X1 U87386 ( .A1(n81425), .A2(n81312), .B1(n81314), .B2(n109719), .ZN(
        n98290) );
  OAI21_X1 U87387 ( .B1(n106202), .B2(n106116), .A(n98291), .ZN(
        \DLX_Datapath/RegisterFile/N23091 ) );
  AOI22_X1 U87388 ( .A1(n81396), .A2(n81312), .B1(n81314), .B2(n109504), .ZN(
        n98291) );
  OAI21_X1 U87389 ( .B1(n106007), .B2(n106202), .A(n98292), .ZN(
        \DLX_Datapath/RegisterFile/N23090 ) );
  AOI22_X1 U87390 ( .A1(n81590), .A2(n81312), .B1(n81314), .B2(n109041), .ZN(
        n98292) );
  OAI21_X1 U87391 ( .B1(n106262), .B2(n106202), .A(n98293), .ZN(
        \DLX_Datapath/RegisterFile/N23089 ) );
  AOI22_X1 U87392 ( .A1(n81423), .A2(n106195), .B1(n81314), .B2(n109389), .ZN(
        n98293) );
  OAI21_X1 U87393 ( .B1(n106202), .B2(n81509), .A(n98294), .ZN(
        \DLX_Datapath/RegisterFile/N23088 ) );
  AOI22_X1 U87394 ( .A1(n81511), .A2(n81312), .B1(n81314), .B2(n109271), .ZN(
        n98294) );
  OAI21_X1 U87395 ( .B1(n106202), .B2(n81501), .A(n98295), .ZN(
        \DLX_Datapath/RegisterFile/N23087 ) );
  AOI22_X1 U87396 ( .A1(n81503), .A2(n81312), .B1(n81314), .B2(n109162), .ZN(
        n98295) );
  OAI21_X1 U87397 ( .B1(n106202), .B2(n106096), .A(n98296), .ZN(
        \DLX_Datapath/RegisterFile/N23086 ) );
  AOI22_X1 U87398 ( .A1(n81417), .A2(n81312), .B1(n81314), .B2(n108698), .ZN(
        n98296) );
  OAI21_X1 U87399 ( .B1(n106202), .B2(n106056), .A(n98297), .ZN(
        \DLX_Datapath/RegisterFile/N23085 ) );
  AOI22_X1 U87400 ( .A1(n81500), .A2(n106196), .B1(n81314), .B2(n108925), .ZN(
        n98297) );
  OAI21_X1 U87401 ( .B1(n105216), .B2(n106202), .A(n98298), .ZN(
        \DLX_Datapath/RegisterFile/N23084 ) );
  AOI22_X1 U87402 ( .A1(n81335), .A2(n106195), .B1(n81314), .B2(n108813), .ZN(
        n98298) );
  OAI21_X1 U87403 ( .B1(n106266), .B2(n106202), .A(n98299), .ZN(
        \DLX_Datapath/RegisterFile/N23083 ) );
  AOI22_X1 U87404 ( .A1(n81327), .A2(n106196), .B1(n81314), .B2(n107353), .ZN(
        n98299) );
  AND2_X2 U87405 ( .A1(n98300), .A2(n98269), .ZN(n81314) );
  AND2_X2 U87406 ( .A1(n98271), .A2(n98300), .ZN(n81312) );
  OR2_X1 U87407 ( .A1(n81309), .A2(n105089), .ZN(n98300) );
  NAND2_X1 U87408 ( .A1(n105124), .A2(n95132), .ZN(n81309) );
  OAI21_X1 U87409 ( .B1(n106149), .B2(n105269), .A(n98302), .ZN(
        \DLX_Datapath/RegisterFile/N23082 ) );
  AOI22_X1 U87410 ( .A1(n98303), .A2(n94667), .B1(n98304), .B2(n107909), .ZN(
        n98302) );
  OAI21_X1 U87411 ( .B1(n105968), .B2(n105269), .A(n98305), .ZN(
        \DLX_Datapath/RegisterFile/N23081 ) );
  AOI22_X1 U87412 ( .A1(n98303), .A2(n94670), .B1(n105267), .B2(n108005), .ZN(
        n98305) );
  OAI21_X1 U87413 ( .B1(n106138), .B2(n105269), .A(n98306), .ZN(
        \DLX_Datapath/RegisterFile/N23080 ) );
  AOI22_X1 U87414 ( .A1(n98303), .A2(n94672), .B1(n105267), .B2(n107276), .ZN(
        n98306) );
  OAI21_X1 U87415 ( .B1(n106211), .B2(n105269), .A(n98307), .ZN(
        \DLX_Datapath/RegisterFile/N23079 ) );
  AOI22_X1 U87416 ( .A1(n98303), .A2(n94674), .B1(n105267), .B2(n107814), .ZN(
        n98307) );
  OAI21_X1 U87417 ( .B1(n106206), .B2(n105269), .A(n98308), .ZN(
        \DLX_Datapath/RegisterFile/N23078 ) );
  AOI22_X1 U87418 ( .A1(n98303), .A2(n94676), .B1(n105267), .B2(n110710), .ZN(
        n98308) );
  OAI21_X1 U87419 ( .B1(n106101), .B2(n105269), .A(n98309), .ZN(
        \DLX_Datapath/RegisterFile/N23077 ) );
  AOI22_X1 U87420 ( .A1(n98303), .A2(n94678), .B1(n105267), .B2(n108113), .ZN(
        n98309) );
  OAI21_X1 U87421 ( .B1(n106257), .B2(n105269), .A(n98310), .ZN(
        \DLX_Datapath/RegisterFile/N23076 ) );
  AOI22_X1 U87422 ( .A1(n98303), .A2(n94680), .B1(n105267), .B2(n110812), .ZN(
        n98310) );
  AOI22_X1 U87424 ( .A1(n98303), .A2(n94682), .B1(n105267), .B2(n110912), .ZN(
        n98311) );
  OAI21_X1 U87425 ( .B1(n106330), .B2(n105269), .A(n98312), .ZN(
        \DLX_Datapath/RegisterFile/N23074 ) );
  AOI22_X1 U87426 ( .A1(n98303), .A2(n94684), .B1(n105267), .B2(n110507), .ZN(
        n98312) );
  OAI21_X1 U87427 ( .B1(n106193), .B2(n105269), .A(n98313), .ZN(
        \DLX_Datapath/RegisterFile/N23073 ) );
  AOI22_X1 U87428 ( .A1(n98303), .A2(n94686), .B1(n105267), .B2(n110290), .ZN(
        n98313) );
  OAI21_X1 U87429 ( .B1(n106131), .B2(n105269), .A(n98314), .ZN(
        \DLX_Datapath/RegisterFile/N23072 ) );
  AOI22_X1 U87430 ( .A1(n98303), .A2(n94688), .B1(n105267), .B2(n110610), .ZN(
        n98314) );
  OAI21_X1 U87431 ( .B1(n106188), .B2(n105269), .A(n98315), .ZN(
        \DLX_Datapath/RegisterFile/N23071 ) );
  AOI22_X1 U87432 ( .A1(n98303), .A2(n94690), .B1(n105267), .B2(n110399), .ZN(
        n98315) );
  OAI21_X1 U87433 ( .B1(n106162), .B2(n105270), .A(n98316), .ZN(
        \DLX_Datapath/RegisterFile/N23070 ) );
  AOI22_X1 U87434 ( .A1(n98303), .A2(n94692), .B1(n98304), .B2(n110077), .ZN(
        n98316) );
  OAI21_X1 U87435 ( .B1(n106106), .B2(n105270), .A(n98317), .ZN(
        \DLX_Datapath/RegisterFile/N23069 ) );
  AOI22_X1 U87436 ( .A1(n98303), .A2(n94694), .B1(n105268), .B2(n110184), .ZN(
        n98317) );
  OAI21_X1 U87437 ( .B1(n106221), .B2(n105270), .A(n98318), .ZN(
        \DLX_Datapath/RegisterFile/N23068 ) );
  AOI22_X1 U87438 ( .A1(n98303), .A2(n94696), .B1(n98304), .B2(n109969), .ZN(
        n98318) );
  OAI21_X1 U87439 ( .B1(n106111), .B2(n105270), .A(n98319), .ZN(
        \DLX_Datapath/RegisterFile/N23067 ) );
  AOI22_X1 U87440 ( .A1(n98303), .A2(n94698), .B1(n105268), .B2(n109852), .ZN(
        n98319) );
  OAI21_X1 U87441 ( .B1(n106233), .B2(n105270), .A(n98320), .ZN(
        \DLX_Datapath/RegisterFile/N23066 ) );
  AOI22_X1 U87442 ( .A1(n98303), .A2(n94700), .B1(n98304), .B2(n108226), .ZN(
        n98320) );
  OAI21_X1 U87443 ( .B1(n106170), .B2(n105270), .A(n98321), .ZN(
        \DLX_Datapath/RegisterFile/N23065 ) );
  AOI22_X1 U87444 ( .A1(n98303), .A2(n94702), .B1(n105268), .B2(n108349), .ZN(
        n98321) );
  OAI21_X1 U87445 ( .B1(n106238), .B2(n105270), .A(n98322), .ZN(
        \DLX_Datapath/RegisterFile/N23064 ) );
  AOI22_X1 U87446 ( .A1(n98303), .A2(n94704), .B1(n98304), .B2(n108460), .ZN(
        n98322) );
  OAI21_X1 U87447 ( .B1(n81451), .B2(n105270), .A(n98323), .ZN(
        \DLX_Datapath/RegisterFile/N23063 ) );
  AOI22_X1 U87448 ( .A1(n98303), .A2(n94706), .B1(n105268), .B2(n107698), .ZN(
        n98323) );
  OAI21_X1 U87449 ( .B1(n106200), .B2(n105270), .A(n98324), .ZN(
        \DLX_Datapath/RegisterFile/N23062 ) );
  AOI22_X1 U87450 ( .A1(n98303), .A2(n94708), .B1(n105267), .B2(n109613), .ZN(
        n98324) );
  OAI21_X1 U87451 ( .B1(n106246), .B2(n105270), .A(n98325), .ZN(
        \DLX_Datapath/RegisterFile/N23061 ) );
  AOI22_X1 U87452 ( .A1(n98303), .A2(n94710), .B1(n105268), .B2(n108575), .ZN(
        n98325) );
  OAI21_X1 U87453 ( .B1(n106157), .B2(n105270), .A(n98326), .ZN(
        \DLX_Datapath/RegisterFile/N23060 ) );
  AOI22_X1 U87454 ( .A1(n98303), .A2(n94712), .B1(n98304), .B2(n109720), .ZN(
        n98326) );
  OAI21_X1 U87455 ( .B1(n106116), .B2(n105270), .A(n98327), .ZN(
        \DLX_Datapath/RegisterFile/N23059 ) );
  AOI22_X1 U87456 ( .A1(n98303), .A2(n94714), .B1(n105268), .B2(n109505), .ZN(
        n98327) );
  OAI21_X1 U87457 ( .B1(n106008), .B2(n105270), .A(n98328), .ZN(
        \DLX_Datapath/RegisterFile/N23058 ) );
  AOI22_X1 U87458 ( .A1(n98303), .A2(n81259), .B1(n98304), .B2(n109042), .ZN(
        n98328) );
  OAI21_X1 U87459 ( .B1(n106262), .B2(n105269), .A(n98329), .ZN(
        \DLX_Datapath/RegisterFile/N23057 ) );
  AOI22_X1 U87460 ( .A1(n98303), .A2(n94717), .B1(n105268), .B2(n109390), .ZN(
        n98329) );
  OAI21_X1 U87461 ( .B1(n106046), .B2(n105270), .A(n98330), .ZN(
        \DLX_Datapath/RegisterFile/N23056 ) );
  AOI22_X1 U87462 ( .A1(n98303), .A2(n94719), .B1(n98304), .B2(n109272), .ZN(
        n98330) );
  OAI21_X1 U87463 ( .B1(n106051), .B2(n105269), .A(n98331), .ZN(
        \DLX_Datapath/RegisterFile/N23055 ) );
  AOI22_X1 U87464 ( .A1(n98303), .A2(n94721), .B1(n105268), .B2(n109163), .ZN(
        n98331) );
  OAI21_X1 U87465 ( .B1(n106096), .B2(n105270), .A(n98332), .ZN(
        \DLX_Datapath/RegisterFile/N23054 ) );
  AOI22_X1 U87466 ( .A1(n98303), .A2(n94723), .B1(n98304), .B2(n108699), .ZN(
        n98332) );
  OAI21_X1 U87467 ( .B1(n106056), .B2(n105270), .A(n98333), .ZN(
        \DLX_Datapath/RegisterFile/N23053 ) );
  AOI22_X1 U87468 ( .A1(n98303), .A2(n94725), .B1(n105268), .B2(n108926), .ZN(
        n98333) );
  OAI21_X1 U87469 ( .B1(n105216), .B2(n105270), .A(n98334), .ZN(
        \DLX_Datapath/RegisterFile/N23052 ) );
  AOI22_X1 U87470 ( .A1(n98303), .A2(n94727), .B1(n105268), .B2(n108814), .ZN(
        n98334) );
  OAI21_X1 U87471 ( .B1(n81262), .B2(n105270), .A(n98335), .ZN(
        \DLX_Datapath/RegisterFile/N23051 ) );
  AOI22_X1 U87472 ( .A1(n98303), .A2(n94729), .B1(n105268), .B2(n107354), .ZN(
        n98335) );
  AND2_X2 U87473 ( .A1(n98269), .A2(n98336), .ZN(n98304) );
  OAI21_X1 U87474 ( .B1(n94366), .B2(n98271), .A(n105602), .ZN(n98269) );
  AND2_X2 U87475 ( .A1(n98271), .A2(n98336), .ZN(n98303) );
  OR2_X1 U87476 ( .A1(n98301), .A2(n105091), .ZN(n98336) );
  NOR2_X1 U87477 ( .A1(n98090), .A2(n95131), .ZN(n98271) );
  NAND2_X1 U87478 ( .A1(n104871), .A2(n94505), .ZN(n98301) );
  OAI21_X1 U87479 ( .B1(n106271), .B2(n106149), .A(n98337), .ZN(
        \DLX_Datapath/RegisterFile/N23050 ) );
  AOI22_X1 U87480 ( .A1(n106265), .A2(n107910), .B1(n81360), .B2(n104880), 
        .ZN(n98337) );
  OAI21_X1 U87481 ( .B1(n106272), .B2(n105970), .A(n98338), .ZN(
        \DLX_Datapath/RegisterFile/N23049 ) );
  AOI22_X1 U87482 ( .A1(n106265), .A2(n108006), .B1(n94511), .B2(n104880), 
        .ZN(n98338) );
  OAI21_X1 U87483 ( .B1(n106271), .B2(n106138), .A(n98339), .ZN(
        \DLX_Datapath/RegisterFile/N23048 ) );
  AOI22_X1 U87484 ( .A1(n106265), .A2(n107277), .B1(n81539), .B2(n104879), 
        .ZN(n98339) );
  OAI21_X1 U87485 ( .B1(n106272), .B2(n81299), .A(n98340), .ZN(
        \DLX_Datapath/RegisterFile/N23047 ) );
  AOI22_X1 U87486 ( .A1(n106265), .A2(n107815), .B1(n81301), .B2(n104879), 
        .ZN(n98340) );
  OAI21_X1 U87487 ( .B1(n106271), .B2(n106204), .A(n98341), .ZN(
        \DLX_Datapath/RegisterFile/N23046 ) );
  AOI22_X1 U87488 ( .A1(n106265), .A2(n110711), .B1(n81308), .B2(n81266), .ZN(
        n98341) );
  OAI21_X1 U87489 ( .B1(n106272), .B2(n106101), .A(n98342), .ZN(
        \DLX_Datapath/RegisterFile/N23045 ) );
  AOI22_X1 U87490 ( .A1(n106265), .A2(n108114), .B1(n94516), .B2(n81266), .ZN(
        n98342) );
  OAI21_X1 U87491 ( .B1(n106272), .B2(n105991), .A(n98343), .ZN(
        \DLX_Datapath/RegisterFile/N23043 ) );
  AOI22_X1 U87492 ( .A1(n106265), .A2(n110913), .B1(n94519), .B2(n104880), 
        .ZN(n98343) );
  OAI21_X1 U87493 ( .B1(n106330), .B2(n106272), .A(n98344), .ZN(
        \DLX_Datapath/RegisterFile/N23042 ) );
  AOI22_X1 U87494 ( .A1(n81264), .A2(n110508), .B1(n104879), .B2(n80192), .ZN(
        n98344) );
  OAI21_X1 U87495 ( .B1(n106272), .B2(n106191), .A(n98345), .ZN(
        \DLX_Datapath/RegisterFile/N23041 ) );
  AOI22_X1 U87496 ( .A1(n81264), .A2(n110291), .B1(n81474), .B2(n104880), .ZN(
        n98345) );
  OAI21_X1 U87497 ( .B1(n106272), .B2(n106130), .A(n98346), .ZN(
        \DLX_Datapath/RegisterFile/N23040 ) );
  AOI22_X1 U87498 ( .A1(n81264), .A2(n110611), .B1(n94523), .B2(n104879), .ZN(
        n98346) );
  OAI21_X1 U87499 ( .B1(n106271), .B2(n106186), .A(n98347), .ZN(
        \DLX_Datapath/RegisterFile/N23039 ) );
  AOI22_X1 U87500 ( .A1(n106264), .A2(n110400), .B1(n106062), .B2(n81266), 
        .ZN(n98347) );
  OAI21_X1 U87501 ( .B1(n106271), .B2(n106164), .A(n98348), .ZN(
        \DLX_Datapath/RegisterFile/N23038 ) );
  AOI22_X1 U87502 ( .A1(n81264), .A2(n110078), .B1(n81347), .B2(n104880), .ZN(
        n98348) );
  OAI21_X1 U87503 ( .B1(n106271), .B2(n106103), .A(n98349), .ZN(
        \DLX_Datapath/RegisterFile/N23037 ) );
  AOI22_X1 U87504 ( .A1(n81264), .A2(n110185), .B1(n94527), .B2(n104880), .ZN(
        n98349) );
  OAI21_X1 U87505 ( .B1(n106271), .B2(n81294), .A(n98350), .ZN(
        \DLX_Datapath/RegisterFile/N23036 ) );
  AOI22_X1 U87506 ( .A1(n106265), .A2(n109970), .B1(n81297), .B2(n104880), 
        .ZN(n98350) );
  OAI21_X1 U87507 ( .B1(n106271), .B2(n106108), .A(n98351), .ZN(
        \DLX_Datapath/RegisterFile/N23035 ) );
  AOI22_X1 U87508 ( .A1(n106265), .A2(n109853), .B1(n94530), .B2(n104879), 
        .ZN(n98351) );
  OAI21_X1 U87509 ( .B1(n106271), .B2(n106233), .A(n98352), .ZN(
        \DLX_Datapath/RegisterFile/N23034 ) );
  AOI22_X1 U87510 ( .A1(n81264), .A2(n108227), .B1(n81286), .B2(n104879), .ZN(
        n98352) );
  OAI21_X1 U87511 ( .B1(n106271), .B2(n81340), .A(n98353), .ZN(
        \DLX_Datapath/RegisterFile/N23033 ) );
  AOI22_X1 U87512 ( .A1(n106265), .A2(n108350), .B1(n106169), .B2(n104880), 
        .ZN(n98353) );
  OAI21_X1 U87513 ( .B1(n106271), .B2(n106236), .A(n98354), .ZN(
        \DLX_Datapath/RegisterFile/N23032 ) );
  AOI22_X1 U87514 ( .A1(n106264), .A2(n108461), .B1(n81283), .B2(n104880), 
        .ZN(n98354) );
  OAI21_X1 U87515 ( .B1(n106271), .B2(n106070), .A(n98355), .ZN(
        \DLX_Datapath/RegisterFile/N23031 ) );
  AOI22_X1 U87516 ( .A1(n106264), .A2(n107699), .B1(n81453), .B2(n81266), .ZN(
        n98355) );
  OAI21_X1 U87517 ( .B1(n106271), .B2(n106198), .A(n98356), .ZN(
        \DLX_Datapath/RegisterFile/N23030 ) );
  AOI22_X1 U87518 ( .A1(n106264), .A2(n109614), .B1(n94536), .B2(n104879), 
        .ZN(n98356) );
  OAI21_X1 U87519 ( .B1(n106271), .B2(n106245), .A(n98357), .ZN(
        \DLX_Datapath/RegisterFile/N23029 ) );
  AOI22_X1 U87520 ( .A1(n106264), .A2(n108576), .B1(n106242), .B2(n81266), 
        .ZN(n98357) );
  OAI21_X1 U87521 ( .B1(n106272), .B2(n106159), .A(n98358), .ZN(
        \DLX_Datapath/RegisterFile/N23028 ) );
  AOI22_X1 U87522 ( .A1(n106264), .A2(n109721), .B1(n81351), .B2(n104879), 
        .ZN(n98358) );
  OAI21_X1 U87523 ( .B1(n106272), .B2(n106115), .A(n98359), .ZN(
        \DLX_Datapath/RegisterFile/N23027 ) );
  AOI22_X1 U87524 ( .A1(n106264), .A2(n109506), .B1(n106021), .B2(n104880), 
        .ZN(n98359) );
  OAI21_X1 U87525 ( .B1(n106010), .B2(n106272), .A(n98360), .ZN(
        \DLX_Datapath/RegisterFile/N23026 ) );
  AOI22_X1 U87526 ( .A1(n106264), .A2(n109043), .B1(n94541), .B2(n81266), .ZN(
        n98360) );
  OAI21_X1 U87527 ( .B1(n106272), .B2(n81509), .A(n98361), .ZN(
        \DLX_Datapath/RegisterFile/N23024 ) );
  AOI22_X1 U87528 ( .A1(n106264), .A2(n109273), .B1(n105625), .B2(n104880), 
        .ZN(n98361) );
  OAI21_X1 U87529 ( .B1(n106272), .B2(n81501), .A(n98362), .ZN(
        \DLX_Datapath/RegisterFile/N23023 ) );
  AOI22_X1 U87530 ( .A1(n106264), .A2(n109164), .B1(n94546), .B2(n104879), 
        .ZN(n98362) );
  OAI21_X1 U87531 ( .B1(n106272), .B2(n106093), .A(n98363), .ZN(
        \DLX_Datapath/RegisterFile/N23022 ) );
  AOI22_X1 U87532 ( .A1(n106264), .A2(n108700), .B1(n94548), .B2(n81266), .ZN(
        n98363) );
  OAI21_X1 U87533 ( .B1(n106272), .B2(n106055), .A(n98364), .ZN(
        \DLX_Datapath/RegisterFile/N23021 ) );
  AOI22_X1 U87534 ( .A1(n106264), .A2(n108927), .B1(n81783), .B2(n104879), 
        .ZN(n98364) );
  OAI21_X1 U87535 ( .B1(n105215), .B2(n106272), .A(n98365), .ZN(
        \DLX_Datapath/RegisterFile/N23020 ) );
  AOI22_X1 U87536 ( .A1(n106264), .A2(n108815), .B1(n81266), .B2(n80188), .ZN(
        n98365) );
  NOR2_X1 U87537 ( .A1(n98366), .A2(n98367), .ZN(n81266) );
  AOI21_X1 U87538 ( .B1(n98087), .B2(n94554), .A(n98367), .ZN(n81264) );
  NOR2_X1 U87539 ( .A1(n81261), .A2(n105095), .ZN(n98367) );
  AND2_X2 U87540 ( .A1(n105602), .A2(n98368), .ZN(n94554) );
  NAND2_X1 U87541 ( .A1(n105124), .A2(n94555), .ZN(n81261) );
  OAI21_X1 U87543 ( .B1(n106149), .B2(n105266), .A(n98371), .ZN(
        \DLX_Datapath/RegisterFile/N23018 ) );
  AOI22_X1 U87544 ( .A1(n104830), .A2(n107911), .B1(n105264), .B2(n94559), 
        .ZN(n98371) );
  OAI21_X1 U87545 ( .B1(n105968), .B2(n105266), .A(n98374), .ZN(
        \DLX_Datapath/RegisterFile/N23017 ) );
  AOI22_X1 U87546 ( .A1(n98372), .A2(n108007), .B1(n105263), .B2(n94562), .ZN(
        n98374) );
  OAI21_X1 U87547 ( .B1(n106138), .B2(n105266), .A(n98375), .ZN(
        \DLX_Datapath/RegisterFile/N23016 ) );
  AOI22_X1 U87548 ( .A1(n98372), .A2(n107278), .B1(n105264), .B2(n94564), .ZN(
        n98375) );
  OAI21_X1 U87549 ( .B1(n106211), .B2(n105266), .A(n98376), .ZN(
        \DLX_Datapath/RegisterFile/N23015 ) );
  AOI22_X1 U87550 ( .A1(n104829), .A2(n107816), .B1(n105263), .B2(n94566), 
        .ZN(n98376) );
  OAI21_X1 U87551 ( .B1(n106206), .B2(n105266), .A(n98377), .ZN(
        \DLX_Datapath/RegisterFile/N23014 ) );
  AOI22_X1 U87552 ( .A1(n104830), .A2(n110712), .B1(n105264), .B2(n94568), 
        .ZN(n98377) );
  OAI21_X1 U87553 ( .B1(n106101), .B2(n105266), .A(n98378), .ZN(
        \DLX_Datapath/RegisterFile/N23013 ) );
  AOI22_X1 U87554 ( .A1(n104829), .A2(n108115), .B1(n105263), .B2(n94570), 
        .ZN(n98378) );
  OAI21_X1 U87555 ( .B1(n106257), .B2(n105266), .A(n98379), .ZN(
        \DLX_Datapath/RegisterFile/N23012 ) );
  AOI22_X1 U87556 ( .A1(n98372), .A2(n110814), .B1(n105264), .B2(n94572), .ZN(
        n98379) );
  OAI21_X1 U87557 ( .B1(n81629), .B2(n105266), .A(n98380), .ZN(
        \DLX_Datapath/RegisterFile/N23011 ) );
  AOI22_X1 U87558 ( .A1(n104829), .A2(n110914), .B1(n105263), .B2(n94574), 
        .ZN(n98380) );
  OAI21_X1 U87559 ( .B1(n106330), .B2(n105266), .A(n98381), .ZN(
        \DLX_Datapath/RegisterFile/N23010 ) );
  AOI22_X1 U87560 ( .A1(n104830), .A2(n110509), .B1(n105263), .B2(n94576), 
        .ZN(n98381) );
  OAI21_X1 U87561 ( .B1(n106192), .B2(n105265), .A(n98382), .ZN(
        \DLX_Datapath/RegisterFile/N23009 ) );
  AOI22_X1 U87562 ( .A1(n104829), .A2(n110292), .B1(n98373), .B2(n94578), .ZN(
        n98382) );
  OAI21_X1 U87563 ( .B1(n106131), .B2(n105265), .A(n98383), .ZN(
        \DLX_Datapath/RegisterFile/N23008 ) );
  AOI22_X1 U87564 ( .A1(n104830), .A2(n110612), .B1(n98373), .B2(n94580), .ZN(
        n98383) );
  OAI21_X1 U87565 ( .B1(n106188), .B2(n105265), .A(n98384), .ZN(
        \DLX_Datapath/RegisterFile/N23007 ) );
  AOI22_X1 U87566 ( .A1(n104830), .A2(n110401), .B1(n105264), .B2(n94582), 
        .ZN(n98384) );
  OAI21_X1 U87567 ( .B1(n106165), .B2(n105265), .A(n98385), .ZN(
        \DLX_Datapath/RegisterFile/N23006 ) );
  AOI22_X1 U87568 ( .A1(n104829), .A2(n110079), .B1(n105263), .B2(n94584), 
        .ZN(n98385) );
  OAI21_X1 U87569 ( .B1(n106106), .B2(n105265), .A(n98386), .ZN(
        \DLX_Datapath/RegisterFile/N23005 ) );
  AOI22_X1 U87570 ( .A1(n104829), .A2(n110186), .B1(n98373), .B2(n94586), .ZN(
        n98386) );
  OAI21_X1 U87571 ( .B1(n106221), .B2(n105265), .A(n98387), .ZN(
        \DLX_Datapath/RegisterFile/N23004 ) );
  AOI22_X1 U87572 ( .A1(n104829), .A2(n109971), .B1(n105263), .B2(n94588), 
        .ZN(n98387) );
  OAI21_X1 U87573 ( .B1(n106111), .B2(n105265), .A(n98388), .ZN(
        \DLX_Datapath/RegisterFile/N23003 ) );
  AOI22_X1 U87574 ( .A1(n104830), .A2(n109854), .B1(n98373), .B2(n94590), .ZN(
        n98388) );
  OAI21_X1 U87575 ( .B1(n106233), .B2(n105265), .A(n98389), .ZN(
        \DLX_Datapath/RegisterFile/N23002 ) );
  AOI22_X1 U87576 ( .A1(n98372), .A2(n108228), .B1(n98373), .B2(n94592), .ZN(
        n98389) );
  OAI21_X1 U87577 ( .B1(n106173), .B2(n105265), .A(n98390), .ZN(
        \DLX_Datapath/RegisterFile/N23001 ) );
  AOI22_X1 U87578 ( .A1(n104830), .A2(n108351), .B1(n98373), .B2(n94594), .ZN(
        n98390) );
  OAI21_X1 U87579 ( .B1(n106238), .B2(n105265), .A(n98391), .ZN(
        \DLX_Datapath/RegisterFile/N23000 ) );
  AOI22_X1 U87580 ( .A1(n104829), .A2(n108462), .B1(n98373), .B2(n94596), .ZN(
        n98391) );
  OAI21_X1 U87581 ( .B1(n106070), .B2(n105265), .A(n98392), .ZN(
        \DLX_Datapath/RegisterFile/N22999 ) );
  AOI22_X1 U87582 ( .A1(n104830), .A2(n107700), .B1(n98373), .B2(n94598), .ZN(
        n98392) );
  OAI21_X1 U87583 ( .B1(n106199), .B2(n105265), .A(n98393), .ZN(
        \DLX_Datapath/RegisterFile/N22998 ) );
  AOI22_X1 U87584 ( .A1(n98372), .A2(n109615), .B1(n105263), .B2(n94600), .ZN(
        n98393) );
  OAI21_X1 U87585 ( .B1(n106246), .B2(n105266), .A(n98394), .ZN(
        \DLX_Datapath/RegisterFile/N22997 ) );
  AOI22_X1 U87586 ( .A1(n98372), .A2(n108577), .B1(n105264), .B2(n94602), .ZN(
        n98394) );
  OAI21_X1 U87587 ( .B1(n106160), .B2(n105266), .A(n98395), .ZN(
        \DLX_Datapath/RegisterFile/N22996 ) );
  AOI22_X1 U87588 ( .A1(n98372), .A2(n109722), .B1(n105263), .B2(n94604), .ZN(
        n98395) );
  OAI21_X1 U87589 ( .B1(n106116), .B2(n105265), .A(n98396), .ZN(
        \DLX_Datapath/RegisterFile/N22995 ) );
  AOI22_X1 U87590 ( .A1(n104829), .A2(n109507), .B1(n105264), .B2(n94606), 
        .ZN(n98396) );
  OAI21_X1 U87591 ( .B1(n106007), .B2(n105266), .A(n98397), .ZN(
        \DLX_Datapath/RegisterFile/N22994 ) );
  AOI22_X1 U87592 ( .A1(n104829), .A2(n109044), .B1(n105263), .B2(n94608), 
        .ZN(n98397) );
  OAI21_X1 U87593 ( .B1(n106262), .B2(n105266), .A(n98398), .ZN(
        \DLX_Datapath/RegisterFile/N22993 ) );
  AOI22_X1 U87594 ( .A1(n104830), .A2(n109392), .B1(n105264), .B2(n94610), 
        .ZN(n98398) );
  OAI21_X1 U87595 ( .B1(n106046), .B2(n105265), .A(n98399), .ZN(
        \DLX_Datapath/RegisterFile/N22992 ) );
  AOI22_X1 U87596 ( .A1(n98372), .A2(n109274), .B1(n105263), .B2(n94612), .ZN(
        n98399) );
  OAI21_X1 U87597 ( .B1(n106051), .B2(n105266), .A(n98400), .ZN(
        \DLX_Datapath/RegisterFile/N22991 ) );
  AOI22_X1 U87598 ( .A1(n104830), .A2(n109165), .B1(n105264), .B2(n94614), 
        .ZN(n98400) );
  OAI21_X1 U87599 ( .B1(n106096), .B2(n105265), .A(n98401), .ZN(
        \DLX_Datapath/RegisterFile/N22990 ) );
  AOI22_X1 U87600 ( .A1(n104829), .A2(n108701), .B1(n105263), .B2(n94616), 
        .ZN(n98401) );
  OAI21_X1 U87601 ( .B1(n106056), .B2(n105266), .A(n98402), .ZN(
        \DLX_Datapath/RegisterFile/N22989 ) );
  AOI22_X1 U87602 ( .A1(n104830), .A2(n108928), .B1(n105264), .B2(n94618), 
        .ZN(n98402) );
  OAI21_X1 U87603 ( .B1(n105215), .B2(n105266), .A(n98403), .ZN(
        \DLX_Datapath/RegisterFile/N22988 ) );
  AOI22_X1 U87604 ( .A1(n104829), .A2(n108816), .B1(n105264), .B2(n94620), 
        .ZN(n98403) );
  OAI21_X1 U87605 ( .B1(n81262), .B2(n105265), .A(n98404), .ZN(
        \DLX_Datapath/RegisterFile/N22987 ) );
  AOI22_X1 U87606 ( .A1(n104829), .A2(n107356), .B1(n105263), .B2(n94622), 
        .ZN(n98404) );
  NOR2_X1 U87607 ( .A1(n98366), .A2(n98405), .ZN(n98373) );
  NOR2_X1 U87608 ( .A1(n98405), .A2(n98406), .ZN(n98372) );
  NOR2_X1 U87609 ( .A1(n98370), .A2(n105093), .ZN(n98405) );
  NAND2_X1 U87610 ( .A1(n94625), .A2(n104871), .ZN(n98370) );
  NOR2_X1 U87611 ( .A1(n98407), .A2(n107128), .ZN(n94625) );
  OAI21_X1 U87612 ( .B1(n106184), .B2(n106146), .A(n98408), .ZN(
        \DLX_Datapath/RegisterFile/N22986 ) );
  AOI22_X1 U87613 ( .A1(n106182), .A2(n107912), .B1(n81521), .B2(n81326), .ZN(
        n98408) );
  OAI21_X1 U87614 ( .B1(n106183), .B2(n105968), .A(n98409), .ZN(
        \DLX_Datapath/RegisterFile/N22985 ) );
  AOI22_X1 U87615 ( .A1(n81325), .A2(n108008), .B1(n81653), .B2(n104881), .ZN(
        n98409) );
  OAI21_X1 U87616 ( .B1(n106184), .B2(n106135), .A(n98410), .ZN(
        \DLX_Datapath/RegisterFile/N22984 ) );
  AOI22_X1 U87617 ( .A1(n81325), .A2(n107279), .B1(n81380), .B2(n104881), .ZN(
        n98410) );
  OAI21_X1 U87618 ( .B1(n106211), .B2(n106184), .A(n98411), .ZN(
        \DLX_Datapath/RegisterFile/N22983 ) );
  AOI22_X1 U87619 ( .A1(n106181), .A2(n107817), .B1(n81377), .B2(n81326), .ZN(
        n98411) );
  OAI21_X1 U87620 ( .B1(n106206), .B2(n106184), .A(n98412), .ZN(
        \DLX_Datapath/RegisterFile/N22982 ) );
  AOI22_X1 U87621 ( .A1(n106181), .A2(n110713), .B1(n81428), .B2(n104881), 
        .ZN(n98412) );
  OAI21_X1 U87622 ( .B1(n106183), .B2(n106100), .A(n98413), .ZN(
        \DLX_Datapath/RegisterFile/N22981 ) );
  AOI22_X1 U87623 ( .A1(n106182), .A2(n108116), .B1(n81410), .B2(n104882), 
        .ZN(n98413) );
  OAI21_X1 U87624 ( .B1(n106257), .B2(n106183), .A(n98414), .ZN(
        \DLX_Datapath/RegisterFile/N22980 ) );
  AOI22_X1 U87625 ( .A1(n106181), .A2(n110815), .B1(n81700), .B2(n104882), 
        .ZN(n98414) );
  OAI21_X1 U87626 ( .B1(n106184), .B2(n105991), .A(n98415), .ZN(
        \DLX_Datapath/RegisterFile/N22979 ) );
  AOI22_X1 U87627 ( .A1(n106182), .A2(n110915), .B1(n81632), .B2(n104882), 
        .ZN(n98415) );
  OAI21_X1 U87628 ( .B1(n80190), .B2(n106183), .A(n98416), .ZN(
        \DLX_Datapath/RegisterFile/N22978 ) );
  AOI22_X1 U87629 ( .A1(n106181), .A2(n110510), .B1(n81414), .B2(n104881), 
        .ZN(n98416) );
  OAI21_X1 U87630 ( .B1(n106193), .B2(n106183), .A(n98417), .ZN(
        \DLX_Datapath/RegisterFile/N22977 ) );
  AOI22_X1 U87631 ( .A1(n106181), .A2(n110293), .B1(n81326), .B2(n81317), .ZN(
        n98417) );
  OAI21_X1 U87632 ( .B1(n106183), .B2(n106129), .A(n98418), .ZN(
        \DLX_Datapath/RegisterFile/N22976 ) );
  AOI22_X1 U87633 ( .A1(n106182), .A2(n110613), .B1(n81386), .B2(n104882), 
        .ZN(n98418) );
  OAI21_X1 U87634 ( .B1(n106184), .B2(n106165), .A(n98419), .ZN(
        \DLX_Datapath/RegisterFile/N22974 ) );
  AOI22_X1 U87635 ( .A1(n106181), .A2(n110080), .B1(n81604), .B2(n104881), 
        .ZN(n98419) );
  OAI21_X1 U87636 ( .B1(n106184), .B2(n106105), .A(n98420), .ZN(
        \DLX_Datapath/RegisterFile/N22973 ) );
  AOI22_X1 U87637 ( .A1(n106182), .A2(n110187), .B1(n81405), .B2(n81326), .ZN(
        n98420) );
  OAI21_X1 U87638 ( .B1(n106221), .B2(n106183), .A(n98421), .ZN(
        \DLX_Datapath/RegisterFile/N22972 ) );
  AOI22_X1 U87639 ( .A1(n106181), .A2(n109972), .B1(n81402), .B2(n104881), 
        .ZN(n98421) );
  OAI21_X1 U87640 ( .B1(n106184), .B2(n106109), .A(n98422), .ZN(
        \DLX_Datapath/RegisterFile/N22971 ) );
  AOI22_X1 U87641 ( .A1(n81325), .A2(n109855), .B1(n81400), .B2(n104882), .ZN(
        n98422) );
  OAI21_X1 U87642 ( .B1(n106183), .B2(n106172), .A(n98423), .ZN(
        \DLX_Datapath/RegisterFile/N22969 ) );
  AOI22_X1 U87643 ( .A1(n106182), .A2(n108352), .B1(n81373), .B2(n104882), 
        .ZN(n98423) );
  OAI21_X1 U87644 ( .B1(n106183), .B2(n106072), .A(n98424), .ZN(
        \DLX_Datapath/RegisterFile/N22967 ) );
  AOI22_X1 U87645 ( .A1(n81325), .A2(n107701), .B1(n81506), .B2(n104881), .ZN(
        n98424) );
  OAI21_X1 U87646 ( .B1(n106200), .B2(n106183), .A(n98425), .ZN(
        \DLX_Datapath/RegisterFile/N22966 ) );
  AOI22_X1 U87647 ( .A1(n106181), .A2(n109616), .B1(n104881), .B2(n81313), 
        .ZN(n98425) );
  OAI21_X1 U87648 ( .B1(n106184), .B2(n106160), .A(n98426), .ZN(
        \DLX_Datapath/RegisterFile/N22964 ) );
  AOI22_X1 U87649 ( .A1(n106182), .A2(n109723), .B1(n81425), .B2(n81326), .ZN(
        n98426) );
  OAI21_X1 U87650 ( .B1(n106183), .B2(n106114), .A(n98427), .ZN(
        \DLX_Datapath/RegisterFile/N22963 ) );
  AOI22_X1 U87651 ( .A1(n106182), .A2(n109508), .B1(n81396), .B2(n104882), 
        .ZN(n98427) );
  OAI21_X1 U87652 ( .B1(n106009), .B2(n106184), .A(n98428), .ZN(
        \DLX_Datapath/RegisterFile/N22962 ) );
  AOI22_X1 U87653 ( .A1(n106181), .A2(n109045), .B1(n81590), .B2(n104882), 
        .ZN(n98428) );
  OAI21_X1 U87654 ( .B1(n106262), .B2(n106184), .A(n98429), .ZN(
        \DLX_Datapath/RegisterFile/N22961 ) );
  AOI22_X1 U87655 ( .A1(n106181), .A2(n109393), .B1(n81423), .B2(n104882), 
        .ZN(n98429) );
  OAI21_X1 U87656 ( .B1(n106183), .B2(n106044), .A(n98430), .ZN(
        \DLX_Datapath/RegisterFile/N22960 ) );
  AOI22_X1 U87657 ( .A1(n106182), .A2(n109275), .B1(n81511), .B2(n104881), 
        .ZN(n98430) );
  OAI21_X1 U87658 ( .B1(n106183), .B2(n81501), .A(n98431), .ZN(
        \DLX_Datapath/RegisterFile/N22959 ) );
  AOI22_X1 U87659 ( .A1(n106181), .A2(n109166), .B1(n81503), .B2(n104881), 
        .ZN(n98431) );
  OAI21_X1 U87660 ( .B1(n106183), .B2(n106094), .A(n98432), .ZN(
        \DLX_Datapath/RegisterFile/N22958 ) );
  AOI22_X1 U87661 ( .A1(n106182), .A2(n108702), .B1(n81417), .B2(n81326), .ZN(
        n98432) );
  OAI21_X1 U87662 ( .B1(n106183), .B2(n81498), .A(n98433), .ZN(
        \DLX_Datapath/RegisterFile/N22957 ) );
  AOI22_X1 U87663 ( .A1(n106182), .A2(n108929), .B1(n81500), .B2(n104882), 
        .ZN(n98433) );
  NOR2_X1 U87664 ( .A1(n98366), .A2(n98434), .ZN(n81326) );
  NOR2_X1 U87665 ( .A1(n98406), .A2(n98434), .ZN(n81325) );
  NOR2_X1 U87666 ( .A1(n81323), .A2(n105094), .ZN(n98434) );
  NAND2_X1 U87667 ( .A1(n104871), .A2(n94664), .ZN(n81323) );
  NOR2_X1 U87668 ( .A1(n98435), .A2(n107128), .ZN(n94664) );
  OAI21_X1 U87669 ( .B1(n106149), .B2(n105262), .A(n98437), .ZN(
        \DLX_Datapath/RegisterFile/N22954 ) );
  AOI22_X1 U87670 ( .A1(n104823), .A2(n94667), .B1(n105259), .B2(n70382), .ZN(
        n98437) );
  OAI21_X1 U87671 ( .B1(n81651), .B2(n105262), .A(n98440), .ZN(
        \DLX_Datapath/RegisterFile/N22953 ) );
  AOI22_X1 U87672 ( .A1(n104824), .A2(n94670), .B1(n105260), .B2(n70524), .ZN(
        n98440) );
  OAI21_X1 U87673 ( .B1(n106138), .B2(n105262), .A(n98441), .ZN(
        \DLX_Datapath/RegisterFile/N22952 ) );
  AOI22_X1 U87674 ( .A1(n104823), .A2(n94672), .B1(n105259), .B2(n69577), .ZN(
        n98441) );
  OAI21_X1 U87675 ( .B1(n106210), .B2(n105262), .A(n98442), .ZN(
        \DLX_Datapath/RegisterFile/N22951 ) );
  AOI22_X1 U87676 ( .A1(n98438), .A2(n94674), .B1(n105260), .B2(n70238), .ZN(
        n98442) );
  OAI21_X1 U87677 ( .B1(n106206), .B2(n105262), .A(n98443), .ZN(
        \DLX_Datapath/RegisterFile/N22950 ) );
  AOI22_X1 U87678 ( .A1(n104823), .A2(n94676), .B1(n105259), .B2(n74084), .ZN(
        n98443) );
  OAI21_X1 U87679 ( .B1(n106101), .B2(n105262), .A(n98444), .ZN(
        \DLX_Datapath/RegisterFile/N22949 ) );
  AOI22_X1 U87680 ( .A1(n104824), .A2(n94678), .B1(n105260), .B2(n70671), .ZN(
        n98444) );
  OAI21_X1 U87681 ( .B1(n106257), .B2(n105262), .A(n98445), .ZN(
        \DLX_Datapath/RegisterFile/N22948 ) );
  AOI22_X1 U87682 ( .A1(n104823), .A2(n94680), .B1(n105259), .B2(n74225), .ZN(
        n98445) );
  OAI21_X1 U87683 ( .B1(n105990), .B2(n105262), .A(n98446), .ZN(
        \DLX_Datapath/RegisterFile/N22947 ) );
  AOI22_X1 U87684 ( .A1(n104823), .A2(n94682), .B1(n105260), .B2(n74365), .ZN(
        n98446) );
  OAI21_X1 U87685 ( .B1(n80190), .B2(n105262), .A(n98447), .ZN(
        \DLX_Datapath/RegisterFile/N22946 ) );
  AOI22_X1 U87686 ( .A1(n104823), .A2(n94684), .B1(n105259), .B2(n73801), .ZN(
        n98447) );
  OAI21_X1 U87687 ( .B1(n106192), .B2(n105261), .A(n98448), .ZN(
        \DLX_Datapath/RegisterFile/N22945 ) );
  AOI22_X1 U87688 ( .A1(n104823), .A2(n94686), .B1(n98439), .B2(n73505), .ZN(
        n98448) );
  OAI21_X1 U87689 ( .B1(n81383), .B2(n105261), .A(n98449), .ZN(
        \DLX_Datapath/RegisterFile/N22944 ) );
  AOI22_X1 U87690 ( .A1(n104824), .A2(n94688), .B1(n105259), .B2(n73942), .ZN(
        n98449) );
  OAI21_X1 U87691 ( .B1(n106188), .B2(n105261), .A(n98450), .ZN(
        \DLX_Datapath/RegisterFile/N22943 ) );
  AOI22_X1 U87692 ( .A1(n104824), .A2(n94690), .B1(n105259), .B2(n73654), .ZN(
        n98450) );
  OAI21_X1 U87693 ( .B1(n106164), .B2(n105261), .A(n98451), .ZN(
        \DLX_Datapath/RegisterFile/N22942 ) );
  AOI22_X1 U87694 ( .A1(n98438), .A2(n94692), .B1(n98439), .B2(n73216), .ZN(
        n98451) );
  OAI21_X1 U87695 ( .B1(n106105), .B2(n105261), .A(n98452), .ZN(
        \DLX_Datapath/RegisterFile/N22941 ) );
  AOI22_X1 U87696 ( .A1(n104823), .A2(n94694), .B1(n98439), .B2(n73358), .ZN(
        n98452) );
  OAI21_X1 U87697 ( .B1(n106220), .B2(n105261), .A(n98453), .ZN(
        \DLX_Datapath/RegisterFile/N22940 ) );
  AOI22_X1 U87698 ( .A1(n104823), .A2(n94696), .B1(n98439), .B2(n73074), .ZN(
        n98453) );
  OAI21_X1 U87699 ( .B1(n106111), .B2(n105261), .A(n98454), .ZN(
        \DLX_Datapath/RegisterFile/N22939 ) );
  AOI22_X1 U87700 ( .A1(n104824), .A2(n94698), .B1(n98439), .B2(n72924), .ZN(
        n98454) );
  OAI21_X1 U87701 ( .B1(n106233), .B2(n105261), .A(n98455), .ZN(
        \DLX_Datapath/RegisterFile/N22938 ) );
  AOI22_X1 U87702 ( .A1(n98438), .A2(n94700), .B1(n98439), .B2(n70820), .ZN(
        n98455) );
  OAI21_X1 U87703 ( .B1(n81340), .B2(n105261), .A(n98456), .ZN(
        \DLX_Datapath/RegisterFile/N22937 ) );
  AOI22_X1 U87704 ( .A1(n104824), .A2(n94702), .B1(n105259), .B2(n70979), .ZN(
        n98456) );
  OAI21_X1 U87705 ( .B1(n106238), .B2(n105261), .A(n98457), .ZN(
        \DLX_Datapath/RegisterFile/N22936 ) );
  AOI22_X1 U87706 ( .A1(n104823), .A2(n94704), .B1(n98439), .B2(n71124), .ZN(
        n98457) );
  OAI21_X1 U87707 ( .B1(n81451), .B2(n105261), .A(n98458), .ZN(
        \DLX_Datapath/RegisterFile/N22935 ) );
  AOI22_X1 U87708 ( .A1(n104824), .A2(n94706), .B1(n105260), .B2(n70085), .ZN(
        n98458) );
  OAI21_X1 U87709 ( .B1(n106199), .B2(n105261), .A(n98459), .ZN(
        \DLX_Datapath/RegisterFile/N22934 ) );
  AOI22_X1 U87710 ( .A1(n98438), .A2(n94708), .B1(n105259), .B2(n72614), .ZN(
        n98459) );
  OAI21_X1 U87711 ( .B1(n106244), .B2(n105262), .A(n98460), .ZN(
        \DLX_Datapath/RegisterFile/N22933 ) );
  AOI22_X1 U87712 ( .A1(n104823), .A2(n94710), .B1(n105260), .B2(n71273), .ZN(
        n98460) );
  OAI21_X1 U87713 ( .B1(n106159), .B2(n105261), .A(n98461), .ZN(
        \DLX_Datapath/RegisterFile/N22932 ) );
  AOI22_X1 U87714 ( .A1(n104824), .A2(n94712), .B1(n105259), .B2(n72756), .ZN(
        n98461) );
  OAI21_X1 U87715 ( .B1(n106116), .B2(n105262), .A(n98462), .ZN(
        \DLX_Datapath/RegisterFile/N22931 ) );
  AOI22_X1 U87716 ( .A1(n104824), .A2(n94714), .B1(n105259), .B2(n72466), .ZN(
        n98462) );
  OAI21_X1 U87717 ( .B1(n106007), .B2(n105262), .A(n98463), .ZN(
        \DLX_Datapath/RegisterFile/N22930 ) );
  AOI22_X1 U87718 ( .A1(n98438), .A2(n81259), .B1(n105260), .B2(n71866), .ZN(
        n98463) );
  OAI21_X1 U87719 ( .B1(n106262), .B2(n105261), .A(n98464), .ZN(
        \DLX_Datapath/RegisterFile/N22929 ) );
  AOI22_X1 U87720 ( .A1(n104823), .A2(n94717), .B1(n105259), .B2(n72315), .ZN(
        n98464) );
  OAI21_X1 U87721 ( .B1(n106045), .B2(n105262), .A(n98465), .ZN(
        \DLX_Datapath/RegisterFile/N22928 ) );
  AOI22_X1 U87722 ( .A1(n104823), .A2(n94719), .B1(n105260), .B2(n72164), .ZN(
        n98465) );
  OAI21_X1 U87723 ( .B1(n106050), .B2(n105261), .A(n98466), .ZN(
        \DLX_Datapath/RegisterFile/N22927 ) );
  AOI22_X1 U87724 ( .A1(n104824), .A2(n94721), .B1(n105259), .B2(n72020), .ZN(
        n98466) );
  OAI21_X1 U87725 ( .B1(n106095), .B2(n105262), .A(n98467), .ZN(
        \DLX_Datapath/RegisterFile/N22926 ) );
  AOI22_X1 U87726 ( .A1(n104824), .A2(n94723), .B1(n105260), .B2(n71422), .ZN(
        n98467) );
  OAI21_X1 U87727 ( .B1(n106056), .B2(n105261), .A(n98468), .ZN(
        \DLX_Datapath/RegisterFile/N22925 ) );
  AOI22_X1 U87728 ( .A1(n98438), .A2(n94725), .B1(n105259), .B2(n71717), .ZN(
        n98468) );
  OAI21_X1 U87729 ( .B1(n105215), .B2(n105262), .A(n98469), .ZN(
        \DLX_Datapath/RegisterFile/N22924 ) );
  AOI22_X1 U87730 ( .A1(n98438), .A2(n94727), .B1(n105260), .B2(n71573), .ZN(
        n98469) );
  OAI21_X1 U87731 ( .B1(n81262), .B2(n105262), .A(n98470), .ZN(
        \DLX_Datapath/RegisterFile/N22923 ) );
  AOI22_X1 U87732 ( .A1(n104823), .A2(n94729), .B1(n105260), .B2(n69682), .ZN(
        n98470) );
  NOR2_X1 U87733 ( .A1(n98406), .A2(n98471), .ZN(n98439) );
  AOI21_X1 U87734 ( .B1(n105205), .B2(n98366), .A(n105601), .ZN(n98406) );
  NOR2_X1 U87735 ( .A1(n98366), .A2(n98471), .ZN(n98438) );
  NOR2_X1 U87736 ( .A1(n98436), .A2(n105093), .ZN(n98471) );
  OR2_X1 U87737 ( .A1(n86230), .A2(n98090), .ZN(n98366) );
  NAND2_X1 U87738 ( .A1(n94734), .A2(n105124), .ZN(n98436) );
  NOR2_X1 U87739 ( .A1(n98472), .A2(n107128), .ZN(n94734) );
  OAI21_X1 U87740 ( .B1(n106252), .B2(n106149), .A(n98473), .ZN(
        \DLX_Datapath/RegisterFile/N22922 ) );
  AOI22_X1 U87741 ( .A1(n70383), .A2(n106251), .B1(n81360), .B2(n81276), .ZN(
        n98473) );
  OAI21_X1 U87742 ( .B1(n106253), .B2(n105970), .A(n98474), .ZN(
        \DLX_Datapath/RegisterFile/N22921 ) );
  AOI22_X1 U87743 ( .A1(n70525), .A2(n106250), .B1(n94511), .B2(n81276), .ZN(
        n98474) );
  OAI21_X1 U87744 ( .B1(n106252), .B2(n106137), .A(n98475), .ZN(
        \DLX_Datapath/RegisterFile/N22920 ) );
  AOI22_X1 U87745 ( .A1(n69578), .A2(n81275), .B1(n81539), .B2(n106248), .ZN(
        n98475) );
  OAI21_X1 U87746 ( .B1(n106252), .B2(n106210), .A(n98476), .ZN(
        \DLX_Datapath/RegisterFile/N22919 ) );
  AOI22_X1 U87747 ( .A1(n70239), .A2(n106251), .B1(n81301), .B2(n81276), .ZN(
        n98476) );
  OAI21_X1 U87748 ( .B1(n106253), .B2(n106204), .A(n98477), .ZN(
        \DLX_Datapath/RegisterFile/N22918 ) );
  AOI22_X1 U87749 ( .A1(n74085), .A2(n106250), .B1(n81308), .B2(n81276), .ZN(
        n98477) );
  OAI21_X1 U87750 ( .B1(n106253), .B2(n106101), .A(n98478), .ZN(
        \DLX_Datapath/RegisterFile/N22917 ) );
  AOI22_X1 U87751 ( .A1(n70672), .A2(n106251), .B1(n94516), .B2(n81276), .ZN(
        n98478) );
  OAI21_X1 U87752 ( .B1(n106257), .B2(n106253), .A(n98479), .ZN(
        \DLX_Datapath/RegisterFile/N22916 ) );
  AOI22_X1 U87753 ( .A1(n74226), .A2(n106251), .B1(n106249), .B2(n81272), .ZN(
        n98479) );
  OAI21_X1 U87754 ( .B1(n106253), .B2(n105992), .A(n98480), .ZN(
        \DLX_Datapath/RegisterFile/N22915 ) );
  AOI22_X1 U87755 ( .A1(n74366), .A2(n106250), .B1(n94519), .B2(n106249), .ZN(
        n98480) );
  OAI21_X1 U87756 ( .B1(n80190), .B2(n106253), .A(n98481), .ZN(
        \DLX_Datapath/RegisterFile/N22914 ) );
  AOI22_X1 U87757 ( .A1(n73802), .A2(n106250), .B1(n106249), .B2(n80192), .ZN(
        n98481) );
  OAI21_X1 U87758 ( .B1(n106253), .B2(n106191), .A(n98482), .ZN(
        \DLX_Datapath/RegisterFile/N22913 ) );
  AOI22_X1 U87759 ( .A1(n73506), .A2(n106251), .B1(n81474), .B2(n81276), .ZN(
        n98482) );
  OAI21_X1 U87760 ( .B1(n106252), .B2(n106130), .A(n98483), .ZN(
        \DLX_Datapath/RegisterFile/N22912 ) );
  AOI22_X1 U87761 ( .A1(n73943), .A2(n81275), .B1(n94523), .B2(n81276), .ZN(
        n98483) );
  OAI21_X1 U87762 ( .B1(n106252), .B2(n106186), .A(n98484), .ZN(
        \DLX_Datapath/RegisterFile/N22911 ) );
  AOI22_X1 U87763 ( .A1(n73655), .A2(n81275), .B1(n106062), .B2(n106248), .ZN(
        n98484) );
  OAI21_X1 U87764 ( .B1(n106252), .B2(n81345), .A(n98485), .ZN(
        \DLX_Datapath/RegisterFile/N22910 ) );
  AOI22_X1 U87765 ( .A1(n73217), .A2(n106251), .B1(n81347), .B2(n106248), .ZN(
        n98485) );
  OAI21_X1 U87766 ( .B1(n106252), .B2(n106105), .A(n98486), .ZN(
        \DLX_Datapath/RegisterFile/N22909 ) );
  AOI22_X1 U87767 ( .A1(n73359), .A2(n81275), .B1(n94527), .B2(n106248), .ZN(
        n98486) );
  OAI21_X1 U87768 ( .B1(n106252), .B2(n106220), .A(n98487), .ZN(
        \DLX_Datapath/RegisterFile/N22908 ) );
  AOI22_X1 U87769 ( .A1(n73075), .A2(n81275), .B1(n81297), .B2(n106248), .ZN(
        n98487) );
  OAI21_X1 U87770 ( .B1(n106252), .B2(n106108), .A(n98488), .ZN(
        \DLX_Datapath/RegisterFile/N22907 ) );
  AOI22_X1 U87771 ( .A1(n72925), .A2(n81275), .B1(n94530), .B2(n106248), .ZN(
        n98488) );
  OAI21_X1 U87772 ( .B1(n106252), .B2(n106173), .A(n98489), .ZN(
        \DLX_Datapath/RegisterFile/N22905 ) );
  AOI22_X1 U87773 ( .A1(n70980), .A2(n106251), .B1(n106169), .B2(n106248), 
        .ZN(n98489) );
  OAI21_X1 U87774 ( .B1(n106252), .B2(n106070), .A(n98490), .ZN(
        \DLX_Datapath/RegisterFile/N22903 ) );
  AOI22_X1 U87775 ( .A1(n70086), .A2(n81275), .B1(n81453), .B2(n106248), .ZN(
        n98490) );
  OAI21_X1 U87776 ( .B1(n106252), .B2(n106198), .A(n98491), .ZN(
        \DLX_Datapath/RegisterFile/N22902 ) );
  AOI22_X1 U87777 ( .A1(n72615), .A2(n106250), .B1(n94536), .B2(n106248), .ZN(
        n98491) );
  OAI21_X1 U87778 ( .B1(n106253), .B2(n81349), .A(n98492), .ZN(
        \DLX_Datapath/RegisterFile/N22900 ) );
  AOI22_X1 U87779 ( .A1(n72757), .A2(n106250), .B1(n81351), .B2(n106248), .ZN(
        n98492) );
  OAI21_X1 U87780 ( .B1(n106252), .B2(n106115), .A(n98493), .ZN(
        \DLX_Datapath/RegisterFile/N22899 ) );
  AOI22_X1 U87781 ( .A1(n72467), .A2(n81275), .B1(n106021), .B2(n106248), .ZN(
        n98493) );
  OAI21_X1 U87782 ( .B1(n106011), .B2(n106253), .A(n98494), .ZN(
        \DLX_Datapath/RegisterFile/N22898 ) );
  AOI22_X1 U87783 ( .A1(n71867), .A2(n106251), .B1(n94541), .B2(n106249), .ZN(
        n98494) );
  OAI21_X1 U87784 ( .B1(n106253), .B2(n106044), .A(n98495), .ZN(
        \DLX_Datapath/RegisterFile/N22896 ) );
  AOI22_X1 U87785 ( .A1(n72165), .A2(n106251), .B1(n105625), .B2(n106249), 
        .ZN(n98495) );
  OAI21_X1 U87786 ( .B1(n106253), .B2(n81501), .A(n98496), .ZN(
        \DLX_Datapath/RegisterFile/N22895 ) );
  AOI22_X1 U87787 ( .A1(n72021), .A2(n106250), .B1(n94546), .B2(n106249), .ZN(
        n98496) );
  OAI21_X1 U87788 ( .B1(n106252), .B2(n106094), .A(n98497), .ZN(
        \DLX_Datapath/RegisterFile/N22894 ) );
  AOI22_X1 U87789 ( .A1(n71423), .A2(n106250), .B1(n94548), .B2(n106248), .ZN(
        n98497) );
  OAI21_X1 U87790 ( .B1(n106252), .B2(n106055), .A(n98498), .ZN(
        \DLX_Datapath/RegisterFile/N22893 ) );
  AOI22_X1 U87791 ( .A1(n71718), .A2(n106250), .B1(n81783), .B2(n81276), .ZN(
        n98498) );
  NOR2_X1 U87792 ( .A1(n98499), .A2(n104694), .ZN(n81276) );
  AOI21_X1 U87793 ( .B1(n98087), .B2(n94771), .A(n98500), .ZN(n81275) );
  NOR2_X1 U87794 ( .A1(n81273), .A2(n105095), .ZN(n98500) );
  AOI21_X1 U87795 ( .B1(n105205), .B2(n94848), .A(n94663), .ZN(n94771) );
  NAND2_X1 U87796 ( .A1(n98090), .A2(n105199), .ZN(n98087) );
  NAND2_X1 U87797 ( .A1(n94772), .A2(n104871), .ZN(n81273) );
  NOR2_X1 U87798 ( .A1(n98501), .A2(n107128), .ZN(n94772) );
  OAI21_X1 U87799 ( .B1(n106147), .B2(n105258), .A(n98503), .ZN(
        \DLX_Datapath/RegisterFile/N22890 ) );
  AOI22_X1 U87800 ( .A1(n104885), .A2(n107913), .B1(n105256), .B2(n94559), 
        .ZN(n98503) );
  OAI21_X1 U87801 ( .B1(n81651), .B2(n105258), .A(n98506), .ZN(
        \DLX_Datapath/RegisterFile/N22889 ) );
  AOI22_X1 U87802 ( .A1(n104885), .A2(n108009), .B1(n105256), .B2(n94562), 
        .ZN(n98506) );
  OAI21_X1 U87803 ( .B1(n81378), .B2(n105258), .A(n98507), .ZN(
        \DLX_Datapath/RegisterFile/N22888 ) );
  AOI22_X1 U87804 ( .A1(n104886), .A2(n107280), .B1(n105255), .B2(n94564), 
        .ZN(n98507) );
  OAI21_X1 U87805 ( .B1(n106211), .B2(n105258), .A(n98508), .ZN(
        \DLX_Datapath/RegisterFile/N22887 ) );
  AOI22_X1 U87806 ( .A1(n104885), .A2(n107818), .B1(n98505), .B2(n94566), .ZN(
        n98508) );
  OAI21_X1 U87807 ( .B1(n106206), .B2(n105258), .A(n98509), .ZN(
        \DLX_Datapath/RegisterFile/N22886 ) );
  AOI22_X1 U87808 ( .A1(n98504), .A2(n110714), .B1(n105256), .B2(n94568), .ZN(
        n98509) );
  OAI21_X1 U87809 ( .B1(n106101), .B2(n105258), .A(n98510), .ZN(
        \DLX_Datapath/RegisterFile/N22885 ) );
  AOI22_X1 U87810 ( .A1(n104886), .A2(n108117), .B1(n98505), .B2(n94570), .ZN(
        n98510) );
  OAI21_X1 U87811 ( .B1(n106257), .B2(n105258), .A(n98511), .ZN(
        \DLX_Datapath/RegisterFile/N22884 ) );
  AOI22_X1 U87812 ( .A1(n98504), .A2(n110816), .B1(n105256), .B2(n94572), .ZN(
        n98511) );
  OAI21_X1 U87813 ( .B1(n105990), .B2(n105258), .A(n98512), .ZN(
        \DLX_Datapath/RegisterFile/N22883 ) );
  AOI22_X1 U87814 ( .A1(n104885), .A2(n110916), .B1(n105255), .B2(n94574), 
        .ZN(n98512) );
  OAI21_X1 U87815 ( .B1(n80190), .B2(n105258), .A(n98513), .ZN(
        \DLX_Datapath/RegisterFile/N22882 ) );
  AOI22_X1 U87816 ( .A1(n104885), .A2(n110511), .B1(n105255), .B2(n94576), 
        .ZN(n98513) );
  OAI21_X1 U87817 ( .B1(n106193), .B2(n105257), .A(n98514), .ZN(
        \DLX_Datapath/RegisterFile/N22881 ) );
  AOI22_X1 U87818 ( .A1(n104886), .A2(n110294), .B1(n105255), .B2(n94578), 
        .ZN(n98514) );
  OAI21_X1 U87819 ( .B1(n106131), .B2(n105257), .A(n98515), .ZN(
        \DLX_Datapath/RegisterFile/N22880 ) );
  AOI22_X1 U87820 ( .A1(n104885), .A2(n110614), .B1(n105255), .B2(n94580), 
        .ZN(n98515) );
  OAI21_X1 U87821 ( .B1(n106188), .B2(n105257), .A(n98516), .ZN(
        \DLX_Datapath/RegisterFile/N22879 ) );
  AOI22_X1 U87822 ( .A1(n104886), .A2(n110403), .B1(n105255), .B2(n94582), 
        .ZN(n98516) );
  OAI21_X1 U87823 ( .B1(n81345), .B2(n105257), .A(n98517), .ZN(
        \DLX_Datapath/RegisterFile/N22878 ) );
  AOI22_X1 U87824 ( .A1(n104886), .A2(n110081), .B1(n105255), .B2(n94584), 
        .ZN(n98517) );
  OAI21_X1 U87825 ( .B1(n106106), .B2(n105257), .A(n98518), .ZN(
        \DLX_Datapath/RegisterFile/N22877 ) );
  AOI22_X1 U87826 ( .A1(n104885), .A2(n110188), .B1(n105255), .B2(n94586), 
        .ZN(n98518) );
  OAI21_X1 U87827 ( .B1(n106221), .B2(n105257), .A(n98519), .ZN(
        \DLX_Datapath/RegisterFile/N22876 ) );
  AOI22_X1 U87828 ( .A1(n104885), .A2(n109973), .B1(n105255), .B2(n94588), 
        .ZN(n98519) );
  OAI21_X1 U87829 ( .B1(n106111), .B2(n105257), .A(n98520), .ZN(
        \DLX_Datapath/RegisterFile/N22875 ) );
  AOI22_X1 U87830 ( .A1(n104885), .A2(n109856), .B1(n105255), .B2(n94590), 
        .ZN(n98520) );
  OAI21_X1 U87831 ( .B1(n106233), .B2(n105257), .A(n98521), .ZN(
        \DLX_Datapath/RegisterFile/N22874 ) );
  AOI22_X1 U87832 ( .A1(n104886), .A2(n108230), .B1(n105255), .B2(n94592), 
        .ZN(n98521) );
  OAI21_X1 U87833 ( .B1(n106173), .B2(n105257), .A(n98522), .ZN(
        \DLX_Datapath/RegisterFile/N22873 ) );
  AOI22_X1 U87834 ( .A1(n104885), .A2(n108353), .B1(n105255), .B2(n94594), 
        .ZN(n98522) );
  OAI21_X1 U87835 ( .B1(n106238), .B2(n105257), .A(n98523), .ZN(
        \DLX_Datapath/RegisterFile/N22872 ) );
  AOI22_X1 U87836 ( .A1(n98504), .A2(n108464), .B1(n105255), .B2(n94596), .ZN(
        n98523) );
  OAI21_X1 U87837 ( .B1(n81451), .B2(n105257), .A(n98524), .ZN(
        \DLX_Datapath/RegisterFile/N22871 ) );
  AOI22_X1 U87838 ( .A1(n104885), .A2(n107702), .B1(n105255), .B2(n94598), 
        .ZN(n98524) );
  OAI21_X1 U87839 ( .B1(n106200), .B2(n105257), .A(n98525), .ZN(
        \DLX_Datapath/RegisterFile/N22870 ) );
  AOI22_X1 U87840 ( .A1(n104886), .A2(n109617), .B1(n98505), .B2(n94600), .ZN(
        n98525) );
  OAI21_X1 U87841 ( .B1(n106245), .B2(n105258), .A(n98526), .ZN(
        \DLX_Datapath/RegisterFile/N22869 ) );
  AOI22_X1 U87842 ( .A1(n104886), .A2(n108579), .B1(n105256), .B2(n94602), 
        .ZN(n98526) );
  OAI21_X1 U87843 ( .B1(n106160), .B2(n105257), .A(n98527), .ZN(
        \DLX_Datapath/RegisterFile/N22868 ) );
  AOI22_X1 U87844 ( .A1(n104886), .A2(n109724), .B1(n98505), .B2(n94604), .ZN(
        n98527) );
  OAI21_X1 U87845 ( .B1(n106116), .B2(n105258), .A(n98528), .ZN(
        \DLX_Datapath/RegisterFile/N22867 ) );
  AOI22_X1 U87846 ( .A1(n104886), .A2(n109509), .B1(n98505), .B2(n94606), .ZN(
        n98528) );
  OAI21_X1 U87847 ( .B1(n106007), .B2(n105258), .A(n98529), .ZN(
        \DLX_Datapath/RegisterFile/N22866 ) );
  AOI22_X1 U87848 ( .A1(n98504), .A2(n109046), .B1(n105256), .B2(n94608), .ZN(
        n98529) );
  OAI21_X1 U87849 ( .B1(n106262), .B2(n105257), .A(n98530), .ZN(
        \DLX_Datapath/RegisterFile/N22865 ) );
  AOI22_X1 U87850 ( .A1(n98504), .A2(n109394), .B1(n105256), .B2(n94610), .ZN(
        n98530) );
  OAI21_X1 U87851 ( .B1(n106046), .B2(n105258), .A(n98531), .ZN(
        \DLX_Datapath/RegisterFile/N22864 ) );
  AOI22_X1 U87852 ( .A1(n104885), .A2(n109276), .B1(n98505), .B2(n94612), .ZN(
        n98531) );
  OAI21_X1 U87853 ( .B1(n106051), .B2(n105257), .A(n98532), .ZN(
        \DLX_Datapath/RegisterFile/N22863 ) );
  AOI22_X1 U87854 ( .A1(n104886), .A2(n109167), .B1(n105256), .B2(n94614), 
        .ZN(n98532) );
  OAI21_X1 U87855 ( .B1(n106096), .B2(n105258), .A(n98533), .ZN(
        \DLX_Datapath/RegisterFile/N22862 ) );
  AOI22_X1 U87856 ( .A1(n104885), .A2(n108703), .B1(n98505), .B2(n94616), .ZN(
        n98533) );
  OAI21_X1 U87857 ( .B1(n106056), .B2(n105257), .A(n98534), .ZN(
        \DLX_Datapath/RegisterFile/N22861 ) );
  AOI22_X1 U87858 ( .A1(n98504), .A2(n108930), .B1(n105256), .B2(n94618), .ZN(
        n98534) );
  OAI21_X1 U87859 ( .B1(n105215), .B2(n105258), .A(n98535), .ZN(
        \DLX_Datapath/RegisterFile/N22860 ) );
  AOI22_X1 U87860 ( .A1(n98504), .A2(n108818), .B1(n105256), .B2(n94620), .ZN(
        n98535) );
  OAI21_X1 U87861 ( .B1(n81262), .B2(n105258), .A(n98536), .ZN(
        \DLX_Datapath/RegisterFile/N22859 ) );
  AOI22_X1 U87862 ( .A1(n104885), .A2(n107358), .B1(n105256), .B2(n94622), 
        .ZN(n98536) );
  NOR2_X1 U87863 ( .A1(n98499), .A2(n98537), .ZN(n98505) );
  NOR2_X1 U87864 ( .A1(n98538), .A2(n98537), .ZN(n98504) );
  NOR2_X1 U87865 ( .A1(n98502), .A2(n105094), .ZN(n98537) );
  NAND2_X1 U87866 ( .A1(n105124), .A2(n94810), .ZN(n98502) );
  NOR2_X1 U87867 ( .A1(n98539), .A2(n107128), .ZN(n94810) );
  OAI21_X1 U87868 ( .B1(n106148), .B2(n105254), .A(n98541), .ZN(
        \DLX_Datapath/RegisterFile/N22858 ) );
  AOI22_X1 U87869 ( .A1(n98542), .A2(n107914), .B1(n105251), .B2(n81521), .ZN(
        n98541) );
  OAI21_X1 U87870 ( .B1(n105971), .B2(n105254), .A(n98544), .ZN(
        \DLX_Datapath/RegisterFile/N22857 ) );
  AOI22_X1 U87871 ( .A1(n104883), .A2(n108010), .B1(n105252), .B2(n81653), 
        .ZN(n98544) );
  OAI21_X1 U87872 ( .B1(n81378), .B2(n105254), .A(n98545), .ZN(
        \DLX_Datapath/RegisterFile/N22856 ) );
  AOI22_X1 U87873 ( .A1(n98542), .A2(n107281), .B1(n105252), .B2(n81380), .ZN(
        n98545) );
  OAI21_X1 U87874 ( .B1(n106211), .B2(n105254), .A(n98546), .ZN(
        \DLX_Datapath/RegisterFile/N22855 ) );
  AOI22_X1 U87875 ( .A1(n104883), .A2(n107819), .B1(n105252), .B2(n81377), 
        .ZN(n98546) );
  OAI21_X1 U87876 ( .B1(n106206), .B2(n105254), .A(n98547), .ZN(
        \DLX_Datapath/RegisterFile/N22854 ) );
  AOI22_X1 U87877 ( .A1(n104884), .A2(n110715), .B1(n105251), .B2(n81428), 
        .ZN(n98547) );
  OAI21_X1 U87878 ( .B1(n81408), .B2(n105254), .A(n98548), .ZN(
        \DLX_Datapath/RegisterFile/N22853 ) );
  AOI22_X1 U87879 ( .A1(n104884), .A2(n108118), .B1(n105251), .B2(n81410), 
        .ZN(n98548) );
  OAI21_X1 U87880 ( .B1(n106257), .B2(n105254), .A(n98549), .ZN(
        \DLX_Datapath/RegisterFile/N22852 ) );
  AOI22_X1 U87881 ( .A1(n98542), .A2(n110817), .B1(n105251), .B2(n81700), .ZN(
        n98549) );
  OAI21_X1 U87882 ( .B1(n105990), .B2(n105254), .A(n98550), .ZN(
        \DLX_Datapath/RegisterFile/N22851 ) );
  AOI22_X1 U87883 ( .A1(n104883), .A2(n110917), .B1(n105252), .B2(n81632), 
        .ZN(n98550) );
  OAI21_X1 U87884 ( .B1(n80190), .B2(n105254), .A(n98551), .ZN(
        \DLX_Datapath/RegisterFile/N22850 ) );
  AOI22_X1 U87885 ( .A1(n104883), .A2(n110512), .B1(n105252), .B2(n81414), 
        .ZN(n98551) );
  OAI21_X1 U87886 ( .B1(n106193), .B2(n105253), .A(n98552), .ZN(
        \DLX_Datapath/RegisterFile/N22849 ) );
  AOI22_X1 U87887 ( .A1(n104883), .A2(n110295), .B1(n98543), .B2(n81317), .ZN(
        n98552) );
  OAI21_X1 U87888 ( .B1(n81383), .B2(n105253), .A(n98553), .ZN(
        \DLX_Datapath/RegisterFile/N22848 ) );
  AOI22_X1 U87889 ( .A1(n98542), .A2(n110615), .B1(n105252), .B2(n81386), .ZN(
        n98553) );
  OAI21_X1 U87890 ( .B1(n106188), .B2(n105253), .A(n98554), .ZN(
        \DLX_Datapath/RegisterFile/N22847 ) );
  AOI22_X1 U87891 ( .A1(n104884), .A2(n110404), .B1(n98543), .B2(n81320), .ZN(
        n98554) );
  OAI21_X1 U87892 ( .B1(n106164), .B2(n105253), .A(n98555), .ZN(
        \DLX_Datapath/RegisterFile/N22846 ) );
  AOI22_X1 U87893 ( .A1(n104884), .A2(n110082), .B1(n98543), .B2(n81604), .ZN(
        n98555) );
  OAI21_X1 U87894 ( .B1(n81403), .B2(n105253), .A(n98556), .ZN(
        \DLX_Datapath/RegisterFile/N22845 ) );
  AOI22_X1 U87895 ( .A1(n104883), .A2(n110189), .B1(n105252), .B2(n81405), 
        .ZN(n98556) );
  OAI21_X1 U87896 ( .B1(n106221), .B2(n105253), .A(n98557), .ZN(
        \DLX_Datapath/RegisterFile/N22844 ) );
  AOI22_X1 U87897 ( .A1(n104883), .A2(n109974), .B1(n105251), .B2(n81402), 
        .ZN(n98557) );
  OAI21_X1 U87898 ( .B1(n81398), .B2(n105253), .A(n98558), .ZN(
        \DLX_Datapath/RegisterFile/N22843 ) );
  AOI22_X1 U87899 ( .A1(n104884), .A2(n109857), .B1(n105252), .B2(n81400), 
        .ZN(n98558) );
  OAI21_X1 U87900 ( .B1(n106233), .B2(n105253), .A(n98559), .ZN(
        \DLX_Datapath/RegisterFile/N22842 ) );
  AOI22_X1 U87901 ( .A1(n104884), .A2(n108231), .B1(n98543), .B2(n81332), .ZN(
        n98559) );
  OAI21_X1 U87902 ( .B1(n106173), .B2(n105253), .A(n98560), .ZN(
        \DLX_Datapath/RegisterFile/N22841 ) );
  AOI22_X1 U87903 ( .A1(n98542), .A2(n108354), .B1(n105251), .B2(n81373), .ZN(
        n98560) );
  OAI21_X1 U87904 ( .B1(n106238), .B2(n105253), .A(n98561), .ZN(
        \DLX_Datapath/RegisterFile/N22840 ) );
  AOI22_X1 U87905 ( .A1(n104883), .A2(n108465), .B1(n105252), .B2(n81322), 
        .ZN(n98561) );
  OAI21_X1 U87906 ( .B1(n81451), .B2(n105253), .A(n98562), .ZN(
        \DLX_Datapath/RegisterFile/N22839 ) );
  AOI22_X1 U87907 ( .A1(n104883), .A2(n107703), .B1(n105251), .B2(n81506), 
        .ZN(n98562) );
  OAI21_X1 U87908 ( .B1(n106200), .B2(n105253), .A(n98563), .ZN(
        \DLX_Datapath/RegisterFile/N22838 ) );
  AOI22_X1 U87909 ( .A1(n104884), .A2(n109618), .B1(n105251), .B2(n81313), 
        .ZN(n98563) );
  OAI21_X1 U87910 ( .B1(n106243), .B2(n105254), .A(n98564), .ZN(
        \DLX_Datapath/RegisterFile/N22837 ) );
  AOI22_X1 U87911 ( .A1(n104884), .A2(n108580), .B1(n98543), .B2(n81330), .ZN(
        n98564) );
  OAI21_X1 U87912 ( .B1(n81349), .B2(n105253), .A(n98565), .ZN(
        \DLX_Datapath/RegisterFile/N22836 ) );
  AOI22_X1 U87913 ( .A1(n104883), .A2(n109725), .B1(n105252), .B2(n81425), 
        .ZN(n98565) );
  OAI21_X1 U87914 ( .B1(n81394), .B2(n105253), .A(n98566), .ZN(
        \DLX_Datapath/RegisterFile/N22835 ) );
  AOI22_X1 U87915 ( .A1(n98542), .A2(n109510), .B1(n98543), .B2(n81396), .ZN(
        n98566) );
  OAI21_X1 U87916 ( .B1(n106007), .B2(n105254), .A(n98567), .ZN(
        \DLX_Datapath/RegisterFile/N22834 ) );
  AOI22_X1 U87917 ( .A1(n104884), .A2(n109047), .B1(n98543), .B2(n81590), .ZN(
        n98567) );
  OAI21_X1 U87918 ( .B1(n106262), .B2(n105254), .A(n98568), .ZN(
        \DLX_Datapath/RegisterFile/N22833 ) );
  AOI22_X1 U87919 ( .A1(n104883), .A2(n109395), .B1(n105251), .B2(n81423), 
        .ZN(n98568) );
  OAI21_X1 U87920 ( .B1(n106046), .B2(n105253), .A(n98569), .ZN(
        \DLX_Datapath/RegisterFile/N22832 ) );
  AOI22_X1 U87921 ( .A1(n104883), .A2(n109277), .B1(n105252), .B2(n81511), 
        .ZN(n98569) );
  OAI21_X1 U87922 ( .B1(n106051), .B2(n105254), .A(n98570), .ZN(
        \DLX_Datapath/RegisterFile/N22831 ) );
  AOI22_X1 U87923 ( .A1(n98542), .A2(n109168), .B1(n105251), .B2(n81503), .ZN(
        n98570) );
  OAI21_X1 U87924 ( .B1(n81415), .B2(n105254), .A(n98571), .ZN(
        \DLX_Datapath/RegisterFile/N22830 ) );
  AOI22_X1 U87925 ( .A1(n104884), .A2(n108704), .B1(n105251), .B2(n81417), 
        .ZN(n98571) );
  OAI21_X1 U87926 ( .B1(n106056), .B2(n105253), .A(n98572), .ZN(
        \DLX_Datapath/RegisterFile/N22829 ) );
  AOI22_X1 U87927 ( .A1(n104884), .A2(n108931), .B1(n98543), .B2(n81500), .ZN(
        n98572) );
  OAI21_X1 U87928 ( .B1(n105215), .B2(n105254), .A(n98573), .ZN(
        \DLX_Datapath/RegisterFile/N22828 ) );
  AOI22_X1 U87929 ( .A1(n104883), .A2(n108819), .B1(n98543), .B2(n81335), .ZN(
        n98573) );
  OAI21_X1 U87930 ( .B1(n81262), .B2(n105254), .A(n98574), .ZN(
        \DLX_Datapath/RegisterFile/N22827 ) );
  AOI22_X1 U87931 ( .A1(n104883), .A2(n107359), .B1(n98543), .B2(n81327), .ZN(
        n98574) );
  NOR2_X1 U87932 ( .A1(n98499), .A2(n98575), .ZN(n98543) );
  NOR2_X1 U87933 ( .A1(n98538), .A2(n98575), .ZN(n98542) );
  NOR2_X1 U87934 ( .A1(n98540), .A2(n105095), .ZN(n98575) );
  NAND2_X1 U87935 ( .A1(n104871), .A2(n94853), .ZN(n98540) );
  NOR2_X1 U87936 ( .A1(n94470), .A2(n107128), .ZN(n94853) );
  OAI21_X1 U87937 ( .B1(n106146), .B2(n105250), .A(n98577), .ZN(
        \DLX_Datapath/RegisterFile/N22826 ) );
  AOI22_X1 U87938 ( .A1(n104826), .A2(n94667), .B1(n105247), .B2(n70386), .ZN(
        n98577) );
  OAI21_X1 U87939 ( .B1(n81651), .B2(n105250), .A(n98580), .ZN(
        \DLX_Datapath/RegisterFile/N22825 ) );
  AOI22_X1 U87940 ( .A1(n104825), .A2(n94670), .B1(n105248), .B2(n108011), 
        .ZN(n98580) );
  OAI21_X1 U87941 ( .B1(n81378), .B2(n105250), .A(n98581), .ZN(
        \DLX_Datapath/RegisterFile/N22824 ) );
  AOI22_X1 U87942 ( .A1(n104825), .A2(n94672), .B1(n105248), .B2(n69581), .ZN(
        n98581) );
  OAI21_X1 U87943 ( .B1(n106211), .B2(n105250), .A(n98582), .ZN(
        \DLX_Datapath/RegisterFile/N22823 ) );
  AOI22_X1 U87944 ( .A1(n104826), .A2(n94674), .B1(n105247), .B2(n70242), .ZN(
        n98582) );
  OAI21_X1 U87945 ( .B1(n106206), .B2(n105250), .A(n98583), .ZN(
        \DLX_Datapath/RegisterFile/N22822 ) );
  AOI22_X1 U87946 ( .A1(n104825), .A2(n94676), .B1(n105248), .B2(n74088), .ZN(
        n98583) );
  OAI21_X1 U87947 ( .B1(n106100), .B2(n105250), .A(n98584), .ZN(
        \DLX_Datapath/RegisterFile/N22821 ) );
  AOI22_X1 U87948 ( .A1(n104825), .A2(n94678), .B1(n105247), .B2(n70675), .ZN(
        n98584) );
  OAI21_X1 U87949 ( .B1(n106257), .B2(n105250), .A(n98585), .ZN(
        \DLX_Datapath/RegisterFile/N22820 ) );
  AOI22_X1 U87950 ( .A1(n98578), .A2(n94680), .B1(n105247), .B2(n74229), .ZN(
        n98585) );
  OAI21_X1 U87951 ( .B1(n105990), .B2(n105250), .A(n98586), .ZN(
        \DLX_Datapath/RegisterFile/N22819 ) );
  AOI22_X1 U87952 ( .A1(n104825), .A2(n94682), .B1(n105248), .B2(n110918), 
        .ZN(n98586) );
  OAI21_X1 U87953 ( .B1(n80190), .B2(n105250), .A(n98587), .ZN(
        \DLX_Datapath/RegisterFile/N22818 ) );
  AOI22_X1 U87954 ( .A1(n104825), .A2(n94684), .B1(n105247), .B2(n73805), .ZN(
        n98587) );
  OAI21_X1 U87955 ( .B1(n106193), .B2(n105249), .A(n98588), .ZN(
        \DLX_Datapath/RegisterFile/N22817 ) );
  AOI22_X1 U87956 ( .A1(n104825), .A2(n94686), .B1(n105247), .B2(n110296), 
        .ZN(n98588) );
  OAI21_X1 U87957 ( .B1(n81383), .B2(n105249), .A(n98589), .ZN(
        \DLX_Datapath/RegisterFile/N22816 ) );
  AOI22_X1 U87958 ( .A1(n104826), .A2(n94688), .B1(n105248), .B2(n110616), 
        .ZN(n98589) );
  OAI21_X1 U87959 ( .B1(n106188), .B2(n105249), .A(n98590), .ZN(
        \DLX_Datapath/RegisterFile/N22815 ) );
  AOI22_X1 U87960 ( .A1(n98578), .A2(n94690), .B1(n98579), .B2(n110405), .ZN(
        n98590) );
  OAI21_X1 U87961 ( .B1(n106165), .B2(n105249), .A(n98591), .ZN(
        \DLX_Datapath/RegisterFile/N22814 ) );
  AOI22_X1 U87962 ( .A1(n98578), .A2(n94692), .B1(n98579), .B2(n110083), .ZN(
        n98591) );
  OAI21_X1 U87963 ( .B1(n106103), .B2(n105249), .A(n98592), .ZN(
        \DLX_Datapath/RegisterFile/N22813 ) );
  AOI22_X1 U87964 ( .A1(n104825), .A2(n94694), .B1(n98579), .B2(n110190), .ZN(
        n98592) );
  OAI21_X1 U87965 ( .B1(n106221), .B2(n105249), .A(n98593), .ZN(
        \DLX_Datapath/RegisterFile/N22812 ) );
  AOI22_X1 U87966 ( .A1(n104825), .A2(n94696), .B1(n105247), .B2(n109975), 
        .ZN(n98593) );
  OAI21_X1 U87967 ( .B1(n106108), .B2(n105249), .A(n98594), .ZN(
        \DLX_Datapath/RegisterFile/N22811 ) );
  AOI22_X1 U87968 ( .A1(n104826), .A2(n94698), .B1(n98579), .B2(n109858), .ZN(
        n98594) );
  OAI21_X1 U87969 ( .B1(n106233), .B2(n105249), .A(n98595), .ZN(
        \DLX_Datapath/RegisterFile/N22810 ) );
  AOI22_X1 U87970 ( .A1(n98578), .A2(n94700), .B1(n98579), .B2(n108232), .ZN(
        n98595) );
  OAI21_X1 U87971 ( .B1(n106172), .B2(n105249), .A(n98596), .ZN(
        \DLX_Datapath/RegisterFile/N22809 ) );
  AOI22_X1 U87972 ( .A1(n104826), .A2(n94702), .B1(n98579), .B2(n108355), .ZN(
        n98596) );
  OAI21_X1 U87973 ( .B1(n106238), .B2(n105249), .A(n98597), .ZN(
        \DLX_Datapath/RegisterFile/N22808 ) );
  AOI22_X1 U87974 ( .A1(n104825), .A2(n94704), .B1(n98579), .B2(n108466), .ZN(
        n98597) );
  OAI21_X1 U87975 ( .B1(n81451), .B2(n105249), .A(n98598), .ZN(
        \DLX_Datapath/RegisterFile/N22807 ) );
  AOI22_X1 U87976 ( .A1(n104826), .A2(n94706), .B1(n105247), .B2(n107704), 
        .ZN(n98598) );
  OAI21_X1 U87977 ( .B1(n106200), .B2(n105249), .A(n98599), .ZN(
        \DLX_Datapath/RegisterFile/N22806 ) );
  AOI22_X1 U87978 ( .A1(n98578), .A2(n94708), .B1(n105247), .B2(n109619), .ZN(
        n98599) );
  OAI21_X1 U87979 ( .B1(n106244), .B2(n105250), .A(n98600), .ZN(
        \DLX_Datapath/RegisterFile/N22805 ) );
  AOI22_X1 U87980 ( .A1(n104825), .A2(n94710), .B1(n105248), .B2(n108581), 
        .ZN(n98600) );
  OAI21_X1 U87981 ( .B1(n106160), .B2(n105249), .A(n98601), .ZN(
        \DLX_Datapath/RegisterFile/N22804 ) );
  AOI22_X1 U87982 ( .A1(n98578), .A2(n94712), .B1(n105247), .B2(n109726), .ZN(
        n98601) );
  OAI21_X1 U87983 ( .B1(n81394), .B2(n105249), .A(n98602), .ZN(
        \DLX_Datapath/RegisterFile/N22803 ) );
  AOI22_X1 U87984 ( .A1(n104826), .A2(n94714), .B1(n105248), .B2(n109511), 
        .ZN(n98602) );
  OAI21_X1 U87985 ( .B1(n81588), .B2(n105250), .A(n98603), .ZN(
        \DLX_Datapath/RegisterFile/N22802 ) );
  AOI22_X1 U87986 ( .A1(n104826), .A2(n81259), .B1(n105247), .B2(n109048), 
        .ZN(n98603) );
  OAI21_X1 U87987 ( .B1(n106262), .B2(n105250), .A(n98604), .ZN(
        \DLX_Datapath/RegisterFile/N22801 ) );
  AOI22_X1 U87988 ( .A1(n104826), .A2(n94717), .B1(n105248), .B2(n109396), 
        .ZN(n98604) );
  OAI21_X1 U87989 ( .B1(n106046), .B2(n105249), .A(n98605), .ZN(
        \DLX_Datapath/RegisterFile/N22800 ) );
  AOI22_X1 U87990 ( .A1(n104825), .A2(n94719), .B1(n105247), .B2(n109278), 
        .ZN(n98605) );
  OAI21_X1 U87991 ( .B1(n106051), .B2(n105250), .A(n98606), .ZN(
        \DLX_Datapath/RegisterFile/N22799 ) );
  AOI22_X1 U87992 ( .A1(n104825), .A2(n94721), .B1(n105248), .B2(n109169), 
        .ZN(n98606) );
  OAI21_X1 U87993 ( .B1(n106094), .B2(n105250), .A(n98607), .ZN(
        \DLX_Datapath/RegisterFile/N22798 ) );
  AOI22_X1 U87994 ( .A1(n104825), .A2(n94723), .B1(n105247), .B2(n108705), 
        .ZN(n98607) );
  OAI21_X1 U87995 ( .B1(n106056), .B2(n105249), .A(n98608), .ZN(
        \DLX_Datapath/RegisterFile/N22797 ) );
  AOI22_X1 U87996 ( .A1(n104826), .A2(n94725), .B1(n105247), .B2(n108932), 
        .ZN(n98608) );
  OAI21_X1 U87997 ( .B1(n105215), .B2(n105250), .A(n98609), .ZN(
        \DLX_Datapath/RegisterFile/N22796 ) );
  AOI22_X1 U87998 ( .A1(n98578), .A2(n94727), .B1(n105248), .B2(n108820), .ZN(
        n98609) );
  OAI21_X1 U87999 ( .B1(n81262), .B2(n105250), .A(n98610), .ZN(
        \DLX_Datapath/RegisterFile/N22795 ) );
  AOI22_X1 U88000 ( .A1(n104826), .A2(n94729), .B1(n105248), .B2(n107360), 
        .ZN(n98610) );
  NOR2_X1 U88001 ( .A1(n98538), .A2(n98611), .ZN(n98579) );
  AOI21_X1 U88002 ( .B1(n105205), .B2(n98499), .A(n94663), .ZN(n98538) );
  NOR2_X1 U88003 ( .A1(n98499), .A2(n98611), .ZN(n98578) );
  NOR2_X1 U88004 ( .A1(n98576), .A2(n105093), .ZN(n98611) );
  OR2_X1 U88005 ( .A1(n94848), .A2(n98090), .ZN(n98499) );
  NAND2_X1 U88006 ( .A1(n98612), .A2(n94851), .ZN(n98090) );
  XOR2_X1 U88007 ( .A(n106764), .B(n98613), .Z(n94851) );
  NOR2_X1 U88008 ( .A1(n107028), .A2(n96488), .ZN(n98612) );
  XNOR2_X1 U88009 ( .A(n98614), .B(n59515), .ZN(n96488) );
  XNOR2_X1 U88010 ( .A(n111027), .B(
        \dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .ZN(n94852) );
  NAND2_X1 U88011 ( .A1(n62212), .A2(n104582), .ZN(n94848) );
  NAND2_X1 U88012 ( .A1(n94892), .A2(n105124), .ZN(n98576) );
  NAND2_X1 U88014 ( .A1(n94895), .A2(n107126), .ZN(n96529) );
  NOR2_X1 U88015 ( .A1(n98615), .A2(n107128), .ZN(n94892) );
  OAI21_X1 U88016 ( .B1(n106147), .B2(n105246), .A(n98617), .ZN(
        \DLX_Datapath/RegisterFile/N22794 ) );
  AOI22_X1 U88017 ( .A1(n105244), .A2(n81360), .B1(n98619), .B2(n107915), .ZN(
        n98617) );
  OAI21_X1 U88018 ( .B1(n81651), .B2(n105246), .A(n98620), .ZN(
        \DLX_Datapath/RegisterFile/N22793 ) );
  AOI22_X1 U88019 ( .A1(n105244), .A2(n94511), .B1(n98619), .B2(n108012), .ZN(
        n98620) );
  OAI21_X1 U88020 ( .B1(n81378), .B2(n105246), .A(n98621), .ZN(
        \DLX_Datapath/RegisterFile/N22792 ) );
  AOI22_X1 U88021 ( .A1(n105244), .A2(n81539), .B1(n98619), .B2(n107282), .ZN(
        n98621) );
  OAI21_X1 U88022 ( .B1(n106211), .B2(n105246), .A(n98622), .ZN(
        \DLX_Datapath/RegisterFile/N22791 ) );
  AOI22_X1 U88023 ( .A1(n105244), .A2(n81301), .B1(n98619), .B2(n107820), .ZN(
        n98622) );
  OAI21_X1 U88024 ( .B1(n106206), .B2(n105246), .A(n98623), .ZN(
        \DLX_Datapath/RegisterFile/N22790 ) );
  AOI22_X1 U88025 ( .A1(n105244), .A2(n81308), .B1(n98619), .B2(n110716), .ZN(
        n98623) );
  OAI21_X1 U88026 ( .B1(n106101), .B2(n105246), .A(n98624), .ZN(
        \DLX_Datapath/RegisterFile/N22789 ) );
  AOI22_X1 U88027 ( .A1(n105244), .A2(n94516), .B1(n98619), .B2(n108119), .ZN(
        n98624) );
  OAI21_X1 U88028 ( .B1(n106254), .B2(n105246), .A(n98625), .ZN(
        \DLX_Datapath/RegisterFile/N22788 ) );
  AOI22_X1 U88029 ( .A1(n105244), .A2(n81272), .B1(n98619), .B2(n110818), .ZN(
        n98625) );
  OAI21_X1 U88030 ( .B1(n105990), .B2(n105246), .A(n98626), .ZN(
        \DLX_Datapath/RegisterFile/N22787 ) );
  AOI22_X1 U88031 ( .A1(n105244), .A2(n94519), .B1(n98619), .B2(n110919), .ZN(
        n98626) );
  OAI21_X1 U88032 ( .B1(n80190), .B2(n105246), .A(n98627), .ZN(
        \DLX_Datapath/RegisterFile/N22786 ) );
  AOI22_X1 U88033 ( .A1(n105243), .A2(n80192), .B1(n105242), .B2(n110513), 
        .ZN(n98627) );
  AND2_X2 U88034 ( .A1(stackBus_In[119]), .A2(n105204), .ZN(n80192) );
  OAI21_X1 U88035 ( .B1(n106193), .B2(n105245), .A(n98628), .ZN(
        \DLX_Datapath/RegisterFile/N22785 ) );
  AOI22_X1 U88036 ( .A1(n105243), .A2(n81474), .B1(n105242), .B2(n110297), 
        .ZN(n98628) );
  OAI21_X1 U88037 ( .B1(n81383), .B2(n105245), .A(n98629), .ZN(
        \DLX_Datapath/RegisterFile/N22784 ) );
  AOI22_X1 U88038 ( .A1(n105243), .A2(n94523), .B1(n105242), .B2(n110617), 
        .ZN(n98629) );
  OAI21_X1 U88039 ( .B1(n106188), .B2(n105245), .A(n98630), .ZN(
        \DLX_Datapath/RegisterFile/N22783 ) );
  AOI22_X1 U88040 ( .A1(n105243), .A2(n106060), .B1(n105242), .B2(n110406), 
        .ZN(n98630) );
  OAI21_X1 U88041 ( .B1(n106163), .B2(n105245), .A(n98631), .ZN(
        \DLX_Datapath/RegisterFile/N22782 ) );
  AOI22_X1 U88042 ( .A1(n98618), .A2(n81347), .B1(n105242), .B2(n110084), .ZN(
        n98631) );
  OAI21_X1 U88043 ( .B1(n106105), .B2(n105245), .A(n98632), .ZN(
        \DLX_Datapath/RegisterFile/N22781 ) );
  AOI22_X1 U88044 ( .A1(n105243), .A2(n94527), .B1(n105242), .B2(n110191), 
        .ZN(n98632) );
  OAI21_X1 U88045 ( .B1(n106221), .B2(n105245), .A(n98633), .ZN(
        \DLX_Datapath/RegisterFile/N22780 ) );
  AOI22_X1 U88046 ( .A1(n105243), .A2(n81297), .B1(n105242), .B2(n109976), 
        .ZN(n98633) );
  OAI21_X1 U88047 ( .B1(n106108), .B2(n105245), .A(n98634), .ZN(
        \DLX_Datapath/RegisterFile/N22779 ) );
  AOI22_X1 U88048 ( .A1(n105243), .A2(n94530), .B1(n105242), .B2(n109859), 
        .ZN(n98634) );
  OAI21_X1 U88049 ( .B1(n106233), .B2(n105245), .A(n98635), .ZN(
        \DLX_Datapath/RegisterFile/N22778 ) );
  AOI22_X1 U88050 ( .A1(n98618), .A2(n81286), .B1(n105242), .B2(n108233), .ZN(
        n98635) );
  OAI21_X1 U88051 ( .B1(n106171), .B2(n105245), .A(n98636), .ZN(
        \DLX_Datapath/RegisterFile/N22777 ) );
  AOI22_X1 U88052 ( .A1(n98618), .A2(n106167), .B1(n105242), .B2(n108356), 
        .ZN(n98636) );
  OAI21_X1 U88053 ( .B1(n106238), .B2(n105245), .A(n98637), .ZN(
        \DLX_Datapath/RegisterFile/N22776 ) );
  AOI22_X1 U88054 ( .A1(n98618), .A2(n81283), .B1(n105242), .B2(n108467), .ZN(
        n98637) );
  OAI21_X1 U88055 ( .B1(n81451), .B2(n105245), .A(n98638), .ZN(
        \DLX_Datapath/RegisterFile/N22775 ) );
  AOI22_X1 U88056 ( .A1(n105243), .A2(n81453), .B1(n105242), .B2(n107705), 
        .ZN(n98638) );
  OAI21_X1 U88057 ( .B1(n106200), .B2(n105245), .A(n98639), .ZN(
        \DLX_Datapath/RegisterFile/N22774 ) );
  AOI22_X1 U88058 ( .A1(n105243), .A2(n105626), .B1(n105241), .B2(n109620), 
        .ZN(n98639) );
  OAI21_X1 U88059 ( .B1(n106243), .B2(n105246), .A(n98640), .ZN(
        \DLX_Datapath/RegisterFile/N22773 ) );
  AOI22_X1 U88060 ( .A1(n105243), .A2(n106240), .B1(n105241), .B2(n108582), 
        .ZN(n98640) );
  OAI21_X1 U88061 ( .B1(n106158), .B2(n105245), .A(n98641), .ZN(
        \DLX_Datapath/RegisterFile/N22772 ) );
  AOI22_X1 U88062 ( .A1(n105243), .A2(n81351), .B1(n105241), .B2(n109727), 
        .ZN(n98641) );
  OAI21_X1 U88063 ( .B1(n81394), .B2(n105245), .A(n98642), .ZN(
        \DLX_Datapath/RegisterFile/N22771 ) );
  AOI22_X1 U88064 ( .A1(n105243), .A2(n106019), .B1(n105241), .B2(n109512), 
        .ZN(n98642) );
  OAI21_X1 U88065 ( .B1(n106007), .B2(n105246), .A(n98643), .ZN(
        \DLX_Datapath/RegisterFile/N22770 ) );
  AOI22_X1 U88066 ( .A1(n105243), .A2(n94541), .B1(n105241), .B2(n109049), 
        .ZN(n98643) );
  OAI21_X1 U88067 ( .B1(n106259), .B2(n105246), .A(n98644), .ZN(
        \DLX_Datapath/RegisterFile/N22769 ) );
  AOI22_X1 U88068 ( .A1(n105243), .A2(n81269), .B1(n105241), .B2(n109397), 
        .ZN(n98644) );
  OAI21_X1 U88069 ( .B1(n106046), .B2(n105246), .A(n98645), .ZN(
        \DLX_Datapath/RegisterFile/N22768 ) );
  AOI22_X1 U88070 ( .A1(n105243), .A2(n105623), .B1(n105241), .B2(n109279), 
        .ZN(n98645) );
  OAI21_X1 U88071 ( .B1(n106051), .B2(n105245), .A(n98646), .ZN(
        \DLX_Datapath/RegisterFile/N22767 ) );
  AOI22_X1 U88072 ( .A1(n105243), .A2(n105622), .B1(n105241), .B2(n109170), 
        .ZN(n98646) );
  OAI21_X1 U88073 ( .B1(n106093), .B2(n105246), .A(n98647), .ZN(
        \DLX_Datapath/RegisterFile/N22766 ) );
  AOI22_X1 U88074 ( .A1(n105243), .A2(n105621), .B1(n105241), .B2(n108706), 
        .ZN(n98647) );
  OAI21_X1 U88075 ( .B1(n106055), .B2(n105246), .A(n98648), .ZN(
        \DLX_Datapath/RegisterFile/N22765 ) );
  AOI22_X1 U88076 ( .A1(n105243), .A2(n105911), .B1(n105241), .B2(n108933), 
        .ZN(n98648) );
  OAI21_X1 U88077 ( .B1(n105215), .B2(n105246), .A(n98649), .ZN(
        \DLX_Datapath/RegisterFile/N22764 ) );
  AOI22_X1 U88078 ( .A1(n105243), .A2(n80188), .B1(n105241), .B2(n108821), 
        .ZN(n98649) );
  AND2_X2 U88079 ( .A1(stackBus_In[97]), .A2(n105204), .ZN(n80188) );
  OAI21_X1 U88080 ( .B1(n106269), .B2(n105245), .A(n98650), .ZN(
        \DLX_Datapath/RegisterFile/N22763 ) );
  AOI22_X1 U88081 ( .A1(n105243), .A2(n81265), .B1(n105241), .B2(n107361), 
        .ZN(n98650) );
  AOI21_X1 U88082 ( .B1(n98651), .B2(n105602), .A(n98652), .ZN(n98619) );
  OAI21_X1 U88083 ( .B1(n94999), .B2(n96489), .A(n105204), .ZN(n98651) );
  NOR2_X1 U88084 ( .A1(n98653), .A2(n94999), .ZN(n98618) );
  OR2_X1 U88085 ( .A1(n98652), .A2(n96489), .ZN(n98653) );
  NOR2_X1 U88086 ( .A1(n98616), .A2(n105094), .ZN(n98652) );
  NAND2_X1 U88087 ( .A1(n94934), .A2(n98654), .ZN(n98616) );
  NOR2_X1 U88088 ( .A1(n98369), .A2(n104762), .ZN(n94934) );
  OR2_X1 U88089 ( .A1(n98655), .A2(n107123), .ZN(n98369) );
  OAI21_X1 U88090 ( .B1(n81358), .B2(n105240), .A(n98657), .ZN(
        \DLX_Datapath/RegisterFile/N22762 ) );
  AOI22_X1 U88091 ( .A1(n98658), .A2(n94559), .B1(n98659), .B2(n70388), .ZN(
        n98657) );
  OAI21_X1 U88092 ( .B1(n105971), .B2(n98656), .A(n98660), .ZN(
        \DLX_Datapath/RegisterFile/N22761 ) );
  AOI22_X1 U88093 ( .A1(n98658), .A2(n94562), .B1(n105239), .B2(n70530), .ZN(
        n98660) );
  OAI21_X1 U88094 ( .B1(n81378), .B2(n105240), .A(n98661), .ZN(
        \DLX_Datapath/RegisterFile/N22760 ) );
  AOI22_X1 U88095 ( .A1(n98658), .A2(n94564), .B1(n105238), .B2(n69583), .ZN(
        n98661) );
  OAI21_X1 U88096 ( .B1(n106211), .B2(n105240), .A(n98662), .ZN(
        \DLX_Datapath/RegisterFile/N22759 ) );
  AOI22_X1 U88097 ( .A1(n98658), .A2(n94566), .B1(n98659), .B2(n70244), .ZN(
        n98662) );
  OAI21_X1 U88098 ( .B1(n106206), .B2(n105240), .A(n98663), .ZN(
        \DLX_Datapath/RegisterFile/N22758 ) );
  AOI22_X1 U88099 ( .A1(n98658), .A2(n94568), .B1(n105239), .B2(n74090), .ZN(
        n98663) );
  OAI21_X1 U88100 ( .B1(n106101), .B2(n98656), .A(n98664), .ZN(
        \DLX_Datapath/RegisterFile/N22757 ) );
  AOI22_X1 U88101 ( .A1(n98658), .A2(n94570), .B1(n105238), .B2(n70677), .ZN(
        n98664) );
  OAI21_X1 U88102 ( .B1(n106257), .B2(n98656), .A(n98665), .ZN(
        \DLX_Datapath/RegisterFile/N22756 ) );
  AOI22_X1 U88103 ( .A1(n98658), .A2(n94572), .B1(n98659), .B2(n74231), .ZN(
        n98665) );
  OAI21_X1 U88104 ( .B1(n105990), .B2(n105240), .A(n98666), .ZN(
        \DLX_Datapath/RegisterFile/N22755 ) );
  AOI22_X1 U88105 ( .A1(n98658), .A2(n94574), .B1(n105238), .B2(n74371), .ZN(
        n98666) );
  OAI21_X1 U88106 ( .B1(n80190), .B2(n105240), .A(n98667), .ZN(
        \DLX_Datapath/RegisterFile/N22754 ) );
  AOI22_X1 U88107 ( .A1(n98658), .A2(n94576), .B1(n105239), .B2(n73807), .ZN(
        n98667) );
  OAI21_X1 U88108 ( .B1(n106193), .B2(n105240), .A(n98668), .ZN(
        \DLX_Datapath/RegisterFile/N22753 ) );
  AOI22_X1 U88109 ( .A1(n98658), .A2(n94578), .B1(n105238), .B2(n73511), .ZN(
        n98668) );
  OAI21_X1 U88110 ( .B1(n106131), .B2(n98656), .A(n98669), .ZN(
        \DLX_Datapath/RegisterFile/N22752 ) );
  AOI22_X1 U88111 ( .A1(n98658), .A2(n94580), .B1(n98659), .B2(n110618), .ZN(
        n98669) );
  OAI21_X1 U88112 ( .B1(n106188), .B2(n105240), .A(n98670), .ZN(
        \DLX_Datapath/RegisterFile/N22751 ) );
  AOI22_X1 U88113 ( .A1(n98658), .A2(n94582), .B1(n105239), .B2(n73660), .ZN(
        n98670) );
  OAI21_X1 U88114 ( .B1(n81345), .B2(n105240), .A(n98671), .ZN(
        \DLX_Datapath/RegisterFile/N22750 ) );
  AOI22_X1 U88115 ( .A1(n98658), .A2(n94584), .B1(n98659), .B2(n73222), .ZN(
        n98671) );
  OAI21_X1 U88116 ( .B1(n106106), .B2(n105240), .A(n98672), .ZN(
        \DLX_Datapath/RegisterFile/N22749 ) );
  AOI22_X1 U88117 ( .A1(n98658), .A2(n94586), .B1(n105239), .B2(n73364), .ZN(
        n98672) );
  OAI21_X1 U88118 ( .B1(n106221), .B2(n105240), .A(n98673), .ZN(
        \DLX_Datapath/RegisterFile/N22748 ) );
  AOI22_X1 U88119 ( .A1(n98658), .A2(n94588), .B1(n105238), .B2(n73080), .ZN(
        n98673) );
  OAI21_X1 U88120 ( .B1(n106111), .B2(n105240), .A(n98674), .ZN(
        \DLX_Datapath/RegisterFile/N22747 ) );
  AOI22_X1 U88121 ( .A1(n98658), .A2(n94590), .B1(n98659), .B2(n72930), .ZN(
        n98674) );
  OAI21_X1 U88122 ( .B1(n106233), .B2(n105240), .A(n98675), .ZN(
        \DLX_Datapath/RegisterFile/N22746 ) );
  AOI22_X1 U88123 ( .A1(n98658), .A2(n94592), .B1(n105239), .B2(n70826), .ZN(
        n98675) );
  OAI21_X1 U88124 ( .B1(n81340), .B2(n105240), .A(n98676), .ZN(
        \DLX_Datapath/RegisterFile/N22745 ) );
  AOI22_X1 U88125 ( .A1(n98658), .A2(n94594), .B1(n105238), .B2(n70985), .ZN(
        n98676) );
  OAI21_X1 U88126 ( .B1(n106238), .B2(n105240), .A(n98677), .ZN(
        \DLX_Datapath/RegisterFile/N22744 ) );
  AOI22_X1 U88127 ( .A1(n98658), .A2(n94596), .B1(n98659), .B2(n71130), .ZN(
        n98677) );
  OAI21_X1 U88128 ( .B1(n81451), .B2(n105240), .A(n98678), .ZN(
        \DLX_Datapath/RegisterFile/N22743 ) );
  AOI22_X1 U88129 ( .A1(n98658), .A2(n94598), .B1(n105239), .B2(n70091), .ZN(
        n98678) );
  OAI21_X1 U88130 ( .B1(n106200), .B2(n105240), .A(n98679), .ZN(
        \DLX_Datapath/RegisterFile/N22742 ) );
  AOI22_X1 U88131 ( .A1(n98658), .A2(n94600), .B1(n105238), .B2(n72620), .ZN(
        n98679) );
  OAI21_X1 U88132 ( .B1(n106245), .B2(n105240), .A(n98680), .ZN(
        \DLX_Datapath/RegisterFile/N22741 ) );
  AOI22_X1 U88133 ( .A1(n98658), .A2(n94602), .B1(n98659), .B2(n71279), .ZN(
        n98680) );
  OAI21_X1 U88134 ( .B1(n81349), .B2(n105240), .A(n98681), .ZN(
        \DLX_Datapath/RegisterFile/N22740 ) );
  AOI22_X1 U88135 ( .A1(n98658), .A2(n94604), .B1(n105239), .B2(n72762), .ZN(
        n98681) );
  OAI21_X1 U88136 ( .B1(n106116), .B2(n105240), .A(n98682), .ZN(
        \DLX_Datapath/RegisterFile/N22739 ) );
  AOI22_X1 U88137 ( .A1(n98658), .A2(n94606), .B1(n105238), .B2(n72472), .ZN(
        n98682) );
  OAI21_X1 U88138 ( .B1(n106011), .B2(n98656), .A(n98683), .ZN(
        \DLX_Datapath/RegisterFile/N22738 ) );
  AOI22_X1 U88139 ( .A1(n98658), .A2(n94608), .B1(n105239), .B2(n71872), .ZN(
        n98683) );
  OAI21_X1 U88140 ( .B1(n106262), .B2(n105240), .A(n98684), .ZN(
        \DLX_Datapath/RegisterFile/N22737 ) );
  AOI22_X1 U88141 ( .A1(n98658), .A2(n94610), .B1(n105238), .B2(n72321), .ZN(
        n98684) );
  OAI21_X1 U88142 ( .B1(n106046), .B2(n105240), .A(n98685), .ZN(
        \DLX_Datapath/RegisterFile/N22736 ) );
  AOI22_X1 U88143 ( .A1(n98658), .A2(n94612), .B1(n98659), .B2(n72170), .ZN(
        n98685) );
  OAI21_X1 U88144 ( .B1(n106051), .B2(n105240), .A(n98686), .ZN(
        \DLX_Datapath/RegisterFile/N22735 ) );
  AOI22_X1 U88145 ( .A1(n98658), .A2(n94614), .B1(n105239), .B2(n72026), .ZN(
        n98686) );
  OAI21_X1 U88146 ( .B1(n106096), .B2(n105240), .A(n98687), .ZN(
        \DLX_Datapath/RegisterFile/N22734 ) );
  AOI22_X1 U88147 ( .A1(n98658), .A2(n94616), .B1(n105238), .B2(n71428), .ZN(
        n98687) );
  OAI21_X1 U88148 ( .B1(n106056), .B2(n98656), .A(n98688), .ZN(
        \DLX_Datapath/RegisterFile/N22733 ) );
  AOI22_X1 U88149 ( .A1(n98658), .A2(n94618), .B1(n98659), .B2(n71723), .ZN(
        n98688) );
  OAI21_X1 U88150 ( .B1(n105215), .B2(n105240), .A(n98689), .ZN(
        \DLX_Datapath/RegisterFile/N22732 ) );
  AOI22_X1 U88151 ( .A1(n98658), .A2(n94620), .B1(n105238), .B2(n71579), .ZN(
        n98689) );
  OAI21_X1 U88152 ( .B1(n106269), .B2(n105240), .A(n98690), .ZN(
        \DLX_Datapath/RegisterFile/N22731 ) );
  AOI22_X1 U88153 ( .A1(n98658), .A2(n94622), .B1(n105239), .B2(n69688), .ZN(
        n98690) );
  AND2_X2 U88154 ( .A1(n98691), .A2(n98692), .ZN(n98659) );
  AND2_X2 U88155 ( .A1(n98693), .A2(n98691), .ZN(n98658) );
  OR2_X1 U88156 ( .A1(n98656), .A2(n105089), .ZN(n98691) );
  NAND2_X1 U88157 ( .A1(n94296), .A2(n98654), .ZN(n98656) );
  NOR2_X1 U88158 ( .A1(n98407), .A2(n104762), .ZN(n94296) );
  OR2_X1 U88159 ( .A1(n98694), .A2(n90120), .ZN(n98407) );
  NAND2_X1 U88160 ( .A1(n90119), .A2(n90127), .ZN(n98694) );
  OAI21_X1 U88161 ( .B1(n81358), .B2(n105237), .A(n98696), .ZN(
        \DLX_Datapath/RegisterFile/N22730 ) );
  AOI22_X1 U88162 ( .A1(n98697), .A2(n107916), .B1(n98698), .B2(n81521), .ZN(
        n98696) );
  OAI21_X1 U88163 ( .B1(n105970), .B2(n105237), .A(n98699), .ZN(
        \DLX_Datapath/RegisterFile/N22729 ) );
  AOI22_X1 U88164 ( .A1(n98697), .A2(n108013), .B1(n98698), .B2(n81653), .ZN(
        n98699) );
  OAI21_X1 U88165 ( .B1(n81378), .B2(n105237), .A(n98700), .ZN(
        \DLX_Datapath/RegisterFile/N22728 ) );
  AOI22_X1 U88166 ( .A1(n98697), .A2(n107283), .B1(n98698), .B2(n81380), .ZN(
        n98700) );
  OAI21_X1 U88167 ( .B1(n106211), .B2(n105237), .A(n98701), .ZN(
        \DLX_Datapath/RegisterFile/N22727 ) );
  AOI22_X1 U88168 ( .A1(n98697), .A2(n107821), .B1(n98698), .B2(n81377), .ZN(
        n98701) );
  OAI21_X1 U88169 ( .B1(n106206), .B2(n105237), .A(n98702), .ZN(
        \DLX_Datapath/RegisterFile/N22726 ) );
  AOI22_X1 U88170 ( .A1(n98697), .A2(n110717), .B1(n98698), .B2(n81428), .ZN(
        n98702) );
  OAI21_X1 U88171 ( .B1(n81408), .B2(n105237), .A(n98703), .ZN(
        \DLX_Datapath/RegisterFile/N22725 ) );
  AOI22_X1 U88172 ( .A1(n98697), .A2(n108120), .B1(n98698), .B2(n81410), .ZN(
        n98703) );
  OAI21_X1 U88173 ( .B1(n106257), .B2(n105237), .A(n98704), .ZN(
        \DLX_Datapath/RegisterFile/N22724 ) );
  AOI22_X1 U88174 ( .A1(n98697), .A2(n110819), .B1(n98698), .B2(n81700), .ZN(
        n98704) );
  OAI21_X1 U88175 ( .B1(n105990), .B2(n105237), .A(n98705), .ZN(
        \DLX_Datapath/RegisterFile/N22723 ) );
  AOI22_X1 U88176 ( .A1(n98697), .A2(n110920), .B1(n98698), .B2(n81632), .ZN(
        n98705) );
  OAI21_X1 U88177 ( .B1(n80190), .B2(n105237), .A(n98706), .ZN(
        \DLX_Datapath/RegisterFile/N22722 ) );
  AOI22_X1 U88178 ( .A1(n98697), .A2(n110514), .B1(n98698), .B2(n81414), .ZN(
        n98706) );
  OAI21_X1 U88179 ( .B1(n106193), .B2(n105237), .A(n98707), .ZN(
        \DLX_Datapath/RegisterFile/N22721 ) );
  AOI22_X1 U88180 ( .A1(n98697), .A2(n110298), .B1(n98698), .B2(n81317), .ZN(
        n98707) );
  OAI21_X1 U88181 ( .B1(n81383), .B2(n105237), .A(n98708), .ZN(
        \DLX_Datapath/RegisterFile/N22720 ) );
  AOI22_X1 U88182 ( .A1(n98697), .A2(n110619), .B1(n98698), .B2(n81386), .ZN(
        n98708) );
  OAI21_X1 U88183 ( .B1(n106188), .B2(n105237), .A(n98709), .ZN(
        \DLX_Datapath/RegisterFile/N22719 ) );
  AOI22_X1 U88184 ( .A1(n98697), .A2(n110407), .B1(n98698), .B2(n81320), .ZN(
        n98709) );
  OAI21_X1 U88185 ( .B1(n81345), .B2(n105237), .A(n98710), .ZN(
        \DLX_Datapath/RegisterFile/N22718 ) );
  AOI22_X1 U88186 ( .A1(n98697), .A2(n110085), .B1(n98698), .B2(n81604), .ZN(
        n98710) );
  OAI21_X1 U88187 ( .B1(n81403), .B2(n105237), .A(n98711), .ZN(
        \DLX_Datapath/RegisterFile/N22717 ) );
  AOI22_X1 U88188 ( .A1(n98697), .A2(n110192), .B1(n98698), .B2(n81405), .ZN(
        n98711) );
  OAI21_X1 U88189 ( .B1(n106221), .B2(n105237), .A(n98712), .ZN(
        \DLX_Datapath/RegisterFile/N22716 ) );
  AOI22_X1 U88190 ( .A1(n98697), .A2(n109977), .B1(n98698), .B2(n81402), .ZN(
        n98712) );
  OAI21_X1 U88191 ( .B1(n81398), .B2(n105237), .A(n98713), .ZN(
        \DLX_Datapath/RegisterFile/N22715 ) );
  AOI22_X1 U88192 ( .A1(n98697), .A2(n109860), .B1(n98698), .B2(n81400), .ZN(
        n98713) );
  OAI21_X1 U88193 ( .B1(n106230), .B2(n105237), .A(n98714), .ZN(
        \DLX_Datapath/RegisterFile/N22714 ) );
  AOI22_X1 U88194 ( .A1(n98697), .A2(n108234), .B1(n98698), .B2(n81332), .ZN(
        n98714) );
  OAI21_X1 U88195 ( .B1(n81340), .B2(n105237), .A(n98715), .ZN(
        \DLX_Datapath/RegisterFile/N22713 ) );
  AOI22_X1 U88196 ( .A1(n98697), .A2(n108357), .B1(n98698), .B2(n81373), .ZN(
        n98715) );
  OAI21_X1 U88197 ( .B1(n106235), .B2(n105237), .A(n98716), .ZN(
        \DLX_Datapath/RegisterFile/N22712 ) );
  AOI22_X1 U88198 ( .A1(n98697), .A2(n108468), .B1(n98698), .B2(n81322), .ZN(
        n98716) );
  OAI21_X1 U88199 ( .B1(n81451), .B2(n105237), .A(n98717), .ZN(
        \DLX_Datapath/RegisterFile/N22711 ) );
  AOI22_X1 U88200 ( .A1(n98697), .A2(n107706), .B1(n98698), .B2(n81506), .ZN(
        n98717) );
  OAI21_X1 U88201 ( .B1(n106200), .B2(n105237), .A(n98718), .ZN(
        \DLX_Datapath/RegisterFile/N22710 ) );
  AOI22_X1 U88202 ( .A1(n98697), .A2(n109621), .B1(n98698), .B2(n81313), .ZN(
        n98718) );
  OAI21_X1 U88203 ( .B1(n106243), .B2(n105237), .A(n98719), .ZN(
        \DLX_Datapath/RegisterFile/N22709 ) );
  AOI22_X1 U88204 ( .A1(n98697), .A2(n108583), .B1(n98698), .B2(n81330), .ZN(
        n98719) );
  OAI21_X1 U88205 ( .B1(n81349), .B2(n105237), .A(n98720), .ZN(
        \DLX_Datapath/RegisterFile/N22708 ) );
  AOI22_X1 U88206 ( .A1(n98697), .A2(n109728), .B1(n98698), .B2(n81425), .ZN(
        n98720) );
  OAI21_X1 U88207 ( .B1(n81394), .B2(n105237), .A(n98721), .ZN(
        \DLX_Datapath/RegisterFile/N22707 ) );
  AOI22_X1 U88208 ( .A1(n98697), .A2(n109513), .B1(n98698), .B2(n81396), .ZN(
        n98721) );
  OAI21_X1 U88209 ( .B1(n106010), .B2(n98695), .A(n98722), .ZN(
        \DLX_Datapath/RegisterFile/N22706 ) );
  AOI22_X1 U88210 ( .A1(n98698), .A2(n81590), .B1(n98697), .B2(n109050), .ZN(
        n98722) );
  AND2_X2 U88211 ( .A1(stackBus_In[39]), .A2(n105203), .ZN(n81590) );
  OAI21_X1 U88212 ( .B1(n106262), .B2(n98695), .A(n98723), .ZN(
        \DLX_Datapath/RegisterFile/N22705 ) );
  AOI22_X1 U88213 ( .A1(n98697), .A2(n109398), .B1(n98698), .B2(n81423), .ZN(
        n98723) );
  OAI21_X1 U88214 ( .B1(n106046), .B2(n98695), .A(n98724), .ZN(
        \DLX_Datapath/RegisterFile/N22704 ) );
  AOI22_X1 U88215 ( .A1(n98697), .A2(n72171), .B1(n98698), .B2(n81511), .ZN(
        n98724) );
  OAI21_X1 U88216 ( .B1(n106051), .B2(n98695), .A(n98725), .ZN(
        \DLX_Datapath/RegisterFile/N22703 ) );
  AOI22_X1 U88217 ( .A1(n98697), .A2(n109171), .B1(n98698), .B2(n81503), .ZN(
        n98725) );
  OAI21_X1 U88218 ( .B1(n81415), .B2(n105237), .A(n98726), .ZN(
        \DLX_Datapath/RegisterFile/N22702 ) );
  AOI22_X1 U88219 ( .A1(n98697), .A2(n71429), .B1(n98698), .B2(n81417), .ZN(
        n98726) );
  OAI21_X1 U88220 ( .B1(n106056), .B2(n98695), .A(n98727), .ZN(
        \DLX_Datapath/RegisterFile/N22701 ) );
  AOI22_X1 U88221 ( .A1(n98698), .A2(n81500), .B1(n98697), .B2(n108934), .ZN(
        n98727) );
  AND2_X2 U88222 ( .A1(stackBus_In[34]), .A2(n105204), .ZN(n81500) );
  OAI21_X1 U88223 ( .B1(n105215), .B2(n105237), .A(n98728), .ZN(
        \DLX_Datapath/RegisterFile/N22700 ) );
  AOI22_X1 U88224 ( .A1(n98697), .A2(n108822), .B1(n98698), .B2(n81335), .ZN(
        n98728) );
  OAI21_X1 U88225 ( .B1(n106269), .B2(n98695), .A(n98729), .ZN(
        \DLX_Datapath/RegisterFile/N22699 ) );
  AOI22_X1 U88226 ( .A1(n98697), .A2(n69689), .B1(n98698), .B2(n81327), .ZN(
        n98729) );
  AND2_X2 U88227 ( .A1(n98693), .A2(n98730), .ZN(n98698) );
  AND2_X2 U88228 ( .A1(n98692), .A2(n98730), .ZN(n98697) );
  OR2_X1 U88229 ( .A1(n98695), .A2(n105089), .ZN(n98730) );
  NAND2_X1 U88230 ( .A1(n94331), .A2(n98654), .ZN(n98695) );
  NOR2_X1 U88231 ( .A1(n98435), .A2(n104762), .ZN(n94331) );
  OR2_X1 U88232 ( .A1(n98731), .A2(n90119), .ZN(n98435) );
  NAND2_X1 U88233 ( .A1(n90120), .A2(n90127), .ZN(n98731) );
  OAI21_X1 U88234 ( .B1(n81358), .B2(n105236), .A(n98733), .ZN(
        \DLX_Datapath/RegisterFile/N22698 ) );
  AOI22_X1 U88235 ( .A1(n98734), .A2(n94667), .B1(n98735), .B2(n107917), .ZN(
        n98733) );
  OAI21_X1 U88236 ( .B1(n105968), .B2(n98732), .A(n98736), .ZN(
        \DLX_Datapath/RegisterFile/N22697 ) );
  AOI22_X1 U88237 ( .A1(n98734), .A2(n94670), .B1(n98735), .B2(n108014), .ZN(
        n98736) );
  OAI21_X1 U88238 ( .B1(n81378), .B2(n105236), .A(n98737), .ZN(
        \DLX_Datapath/RegisterFile/N22696 ) );
  AOI22_X1 U88239 ( .A1(n98734), .A2(n94672), .B1(n98735), .B2(n107284), .ZN(
        n98737) );
  OAI21_X1 U88240 ( .B1(n106208), .B2(n105236), .A(n98738), .ZN(
        \DLX_Datapath/RegisterFile/N22695 ) );
  AOI22_X1 U88241 ( .A1(n98734), .A2(n94674), .B1(n98735), .B2(n107822), .ZN(
        n98738) );
  OAI21_X1 U88242 ( .B1(n106203), .B2(n105236), .A(n98739), .ZN(
        \DLX_Datapath/RegisterFile/N22694 ) );
  AOI22_X1 U88243 ( .A1(n98734), .A2(n94676), .B1(n98735), .B2(n110718), .ZN(
        n98739) );
  OAI21_X1 U88244 ( .B1(n81408), .B2(n105236), .A(n98740), .ZN(
        \DLX_Datapath/RegisterFile/N22693 ) );
  AOI22_X1 U88245 ( .A1(n98734), .A2(n94678), .B1(n98735), .B2(n108121), .ZN(
        n98740) );
  OAI21_X1 U88246 ( .B1(n106256), .B2(n105236), .A(n98741), .ZN(
        \DLX_Datapath/RegisterFile/N22692 ) );
  AOI22_X1 U88247 ( .A1(n98734), .A2(n94680), .B1(n98735), .B2(n110820), .ZN(
        n98741) );
  OAI21_X1 U88248 ( .B1(n105990), .B2(n105236), .A(n98742), .ZN(
        \DLX_Datapath/RegisterFile/N22691 ) );
  AOI22_X1 U88249 ( .A1(n98734), .A2(n94682), .B1(n98735), .B2(n110921), .ZN(
        n98742) );
  OAI21_X1 U88250 ( .B1(n80190), .B2(n105236), .A(n98743), .ZN(
        \DLX_Datapath/RegisterFile/N22690 ) );
  AOI22_X1 U88251 ( .A1(n98734), .A2(n94684), .B1(n98735), .B2(n110515), .ZN(
        n98743) );
  OAI21_X1 U88252 ( .B1(n106193), .B2(n98732), .A(n98744), .ZN(
        \DLX_Datapath/RegisterFile/N22689 ) );
  AOI22_X1 U88253 ( .A1(n98734), .A2(n94686), .B1(n98735), .B2(n110299), .ZN(
        n98744) );
  OAI21_X1 U88254 ( .B1(n81383), .B2(n105236), .A(n98745), .ZN(
        \DLX_Datapath/RegisterFile/N22688 ) );
  AOI22_X1 U88255 ( .A1(n98734), .A2(n94688), .B1(n98735), .B2(n110620), .ZN(
        n98745) );
  OAI21_X1 U88256 ( .B1(n106188), .B2(n98732), .A(n98746), .ZN(
        \DLX_Datapath/RegisterFile/N22687 ) );
  AOI22_X1 U88257 ( .A1(n98734), .A2(n94690), .B1(n98735), .B2(n110408), .ZN(
        n98746) );
  OAI21_X1 U88258 ( .B1(n81345), .B2(n105236), .A(n98747), .ZN(
        \DLX_Datapath/RegisterFile/N22686 ) );
  AOI22_X1 U88259 ( .A1(n98734), .A2(n94692), .B1(n98735), .B2(n110086), .ZN(
        n98747) );
  OAI21_X1 U88260 ( .B1(n81403), .B2(n105236), .A(n98748), .ZN(
        \DLX_Datapath/RegisterFile/N22685 ) );
  AOI22_X1 U88261 ( .A1(n98734), .A2(n94694), .B1(n98735), .B2(n110193), .ZN(
        n98748) );
  OAI21_X1 U88262 ( .B1(n106218), .B2(n105236), .A(n98749), .ZN(
        \DLX_Datapath/RegisterFile/N22684 ) );
  AOI22_X1 U88263 ( .A1(n98734), .A2(n94696), .B1(n98735), .B2(n109978), .ZN(
        n98749) );
  OAI21_X1 U88264 ( .B1(n81398), .B2(n105236), .A(n98750), .ZN(
        \DLX_Datapath/RegisterFile/N22683 ) );
  AOI22_X1 U88265 ( .A1(n98734), .A2(n94698), .B1(n98735), .B2(n109861), .ZN(
        n98750) );
  OAI21_X1 U88266 ( .B1(n106231), .B2(n105236), .A(n98751), .ZN(
        \DLX_Datapath/RegisterFile/N22682 ) );
  AOI22_X1 U88267 ( .A1(n98734), .A2(n94700), .B1(n98735), .B2(n108235), .ZN(
        n98751) );
  OAI21_X1 U88268 ( .B1(n81340), .B2(n105236), .A(n98752), .ZN(
        \DLX_Datapath/RegisterFile/N22681 ) );
  AOI22_X1 U88269 ( .A1(n98734), .A2(n94702), .B1(n98735), .B2(n108358), .ZN(
        n98752) );
  OAI21_X1 U88270 ( .B1(n106237), .B2(n105236), .A(n98753), .ZN(
        \DLX_Datapath/RegisterFile/N22680 ) );
  AOI22_X1 U88271 ( .A1(n98734), .A2(n94704), .B1(n98735), .B2(n108469), .ZN(
        n98753) );
  OAI21_X1 U88272 ( .B1(n81451), .B2(n105236), .A(n98754), .ZN(
        \DLX_Datapath/RegisterFile/N22679 ) );
  AOI22_X1 U88273 ( .A1(n98734), .A2(n94706), .B1(n98735), .B2(n107707), .ZN(
        n98754) );
  OAI21_X1 U88274 ( .B1(n106200), .B2(n105236), .A(n98755), .ZN(
        \DLX_Datapath/RegisterFile/N22678 ) );
  AOI22_X1 U88275 ( .A1(n98734), .A2(n94708), .B1(n98735), .B2(n109622), .ZN(
        n98755) );
  OAI21_X1 U88276 ( .B1(n106244), .B2(n105236), .A(n98756), .ZN(
        \DLX_Datapath/RegisterFile/N22677 ) );
  AOI22_X1 U88277 ( .A1(n98734), .A2(n94710), .B1(n98735), .B2(n108584), .ZN(
        n98756) );
  OAI21_X1 U88278 ( .B1(n81349), .B2(n105236), .A(n98757), .ZN(
        \DLX_Datapath/RegisterFile/N22676 ) );
  AOI22_X1 U88279 ( .A1(n98734), .A2(n94712), .B1(n98735), .B2(n109729), .ZN(
        n98757) );
  OAI21_X1 U88280 ( .B1(n81394), .B2(n105236), .A(n98758), .ZN(
        \DLX_Datapath/RegisterFile/N22675 ) );
  AOI22_X1 U88281 ( .A1(n98734), .A2(n94714), .B1(n98735), .B2(n109514), .ZN(
        n98758) );
  OAI21_X1 U88282 ( .B1(n81588), .B2(n105236), .A(n98759), .ZN(
        \DLX_Datapath/RegisterFile/N22674 ) );
  AOI22_X1 U88283 ( .A1(n98734), .A2(n81259), .B1(n98735), .B2(n109051), .ZN(
        n98759) );
  AND2_X2 U88284 ( .A1(stackBus_In[7]), .A2(n105204), .ZN(n81259) );
  OAI21_X1 U88285 ( .B1(n106261), .B2(n98732), .A(n98760), .ZN(
        \DLX_Datapath/RegisterFile/N22673 ) );
  AOI22_X1 U88286 ( .A1(n98734), .A2(n94717), .B1(n98735), .B2(n109399), .ZN(
        n98760) );
  OAI21_X1 U88287 ( .B1(n106046), .B2(n98732), .A(n98761), .ZN(
        \DLX_Datapath/RegisterFile/N22672 ) );
  AOI22_X1 U88288 ( .A1(n98734), .A2(n94719), .B1(n98735), .B2(n109280), .ZN(
        n98761) );
  OAI21_X1 U88289 ( .B1(n106051), .B2(n98732), .A(n98762), .ZN(
        \DLX_Datapath/RegisterFile/N22671 ) );
  AOI22_X1 U88290 ( .A1(n98734), .A2(n94721), .B1(n98735), .B2(n109172), .ZN(
        n98762) );
  OAI21_X1 U88291 ( .B1(n81415), .B2(n105236), .A(n98763), .ZN(
        \DLX_Datapath/RegisterFile/N22670 ) );
  AOI22_X1 U88292 ( .A1(n98734), .A2(n94723), .B1(n98735), .B2(n108707), .ZN(
        n98763) );
  OAI21_X1 U88293 ( .B1(n106056), .B2(n105236), .A(n98764), .ZN(
        \DLX_Datapath/RegisterFile/N22669 ) );
  AOI22_X1 U88294 ( .A1(n98734), .A2(n94725), .B1(n98735), .B2(n108935), .ZN(
        n98764) );
  OAI21_X1 U88295 ( .B1(n105215), .B2(n105236), .A(n98765), .ZN(
        \DLX_Datapath/RegisterFile/N22668 ) );
  AOI22_X1 U88296 ( .A1(n98734), .A2(n94727), .B1(n98735), .B2(n108823), .ZN(
        n98765) );
  OAI21_X1 U88297 ( .B1(n106266), .B2(n105236), .A(n98766), .ZN(
        \DLX_Datapath/RegisterFile/N22667 ) );
  AOI22_X1 U88298 ( .A1(n98734), .A2(n94729), .B1(n98735), .B2(n107362), .ZN(
        n98766) );
  AND2_X2 U88299 ( .A1(n98692), .A2(n98767), .ZN(n98735) );
  OAI21_X1 U88300 ( .B1(n98693), .B2(n94366), .A(n105602), .ZN(n98692) );
  AND2_X2 U88301 ( .A1(n98693), .A2(n98767), .ZN(n98734) );
  OR2_X1 U88302 ( .A1(n98732), .A2(n105092), .ZN(n98767) );
  NOR2_X1 U88303 ( .A1(n94999), .A2(n96489), .ZN(n98693) );
  NAND2_X1 U88304 ( .A1(n62190), .A2(n111027), .ZN(n94999) );
  NAND2_X1 U88305 ( .A1(n94367), .A2(n98654), .ZN(n98732) );
  NOR2_X1 U88306 ( .A1(n98472), .A2(n104762), .ZN(n94367) );
  OR2_X1 U88307 ( .A1(n98768), .A2(n90120), .ZN(n98472) );
  NAND2_X1 U88308 ( .A1(n90127), .A2(n107122), .ZN(n98768) );
  OAI21_X1 U88309 ( .B1(n106341), .B2(n81358), .A(n98769), .ZN(
        \DLX_Datapath/RegisterFile/N22666 ) );
  AOI22_X1 U88310 ( .A1(n81360), .A2(n106338), .B1(n106337), .B2(n107918), 
        .ZN(n98769) );
  AND2_X2 U88311 ( .A1(stackBus_In[127]), .A2(n105204), .ZN(n81360) );
  OAI21_X1 U88312 ( .B1(n106341), .B2(n81651), .A(n98770), .ZN(
        \DLX_Datapath/RegisterFile/N22665 ) );
  AOI22_X1 U88313 ( .A1(n94511), .A2(n106338), .B1(n106337), .B2(n108015), 
        .ZN(n98770) );
  AND2_X2 U88314 ( .A1(stackBus_In[126]), .A2(n105204), .ZN(n94511) );
  OAI21_X1 U88315 ( .B1(n106341), .B2(n106136), .A(n98771), .ZN(
        \DLX_Datapath/RegisterFile/N22664 ) );
  AOI22_X1 U88316 ( .A1(n81539), .A2(n106338), .B1(n106337), .B2(n107285), 
        .ZN(n98771) );
  AND2_X2 U88317 ( .A1(stackBus_In[125]), .A2(n105204), .ZN(n81539) );
  OAI21_X1 U88318 ( .B1(n106341), .B2(n106210), .A(n98772), .ZN(
        \DLX_Datapath/RegisterFile/N22663 ) );
  AOI22_X1 U88319 ( .A1(n81301), .A2(n106338), .B1(n106337), .B2(n107823), 
        .ZN(n98772) );
  AND2_X2 U88320 ( .A1(stackBus_In[124]), .A2(n105203), .ZN(n81301) );
  OAI21_X1 U88321 ( .B1(n106341), .B2(n81306), .A(n98773), .ZN(
        \DLX_Datapath/RegisterFile/N22662 ) );
  AOI22_X1 U88322 ( .A1(n81308), .A2(n106338), .B1(n106337), .B2(n110719), 
        .ZN(n98773) );
  AND2_X2 U88323 ( .A1(stackBus_In[123]), .A2(n105204), .ZN(n81308) );
  OAI21_X1 U88324 ( .B1(n106341), .B2(n81408), .A(n98774), .ZN(
        \DLX_Datapath/RegisterFile/N22661 ) );
  AOI22_X1 U88325 ( .A1(n94516), .A2(n106338), .B1(n106337), .B2(n108122), 
        .ZN(n98774) );
  AND2_X2 U88326 ( .A1(stackBus_In[122]), .A2(n105203), .ZN(n94516) );
  OAI21_X1 U88327 ( .B1(n106341), .B2(n106255), .A(n98775), .ZN(
        \DLX_Datapath/RegisterFile/N22660 ) );
  AOI22_X1 U88328 ( .A1(n81272), .A2(n106339), .B1(n106336), .B2(n110821), 
        .ZN(n98775) );
  AND2_X2 U88329 ( .A1(stackBus_In[121]), .A2(n105203), .ZN(n81272) );
  OAI21_X1 U88330 ( .B1(n106341), .B2(n105992), .A(n98776), .ZN(
        \DLX_Datapath/RegisterFile/N22659 ) );
  AOI22_X1 U88331 ( .A1(n94519), .A2(n106339), .B1(n106336), .B2(n110922), 
        .ZN(n98776) );
  AND2_X2 U88332 ( .A1(stackBus_In[120]), .A2(n105203), .ZN(n94519) );
  OAI21_X1 U88333 ( .B1(n106341), .B2(n106190), .A(n98777), .ZN(
        \DLX_Datapath/RegisterFile/N22657 ) );
  AOI22_X1 U88334 ( .A1(n81474), .A2(n106340), .B1(n106336), .B2(n110300), 
        .ZN(n98777) );
  AND2_X2 U88335 ( .A1(stackBus_In[118]), .A2(n105203), .ZN(n81474) );
  OAI21_X1 U88336 ( .B1(n106341), .B2(n106131), .A(n98778), .ZN(
        \DLX_Datapath/RegisterFile/N22656 ) );
  AOI22_X1 U88337 ( .A1(n94523), .A2(n106339), .B1(n106336), .B2(n110621), 
        .ZN(n98778) );
  AND2_X2 U88338 ( .A1(stackBus_In[117]), .A2(n105203), .ZN(n94523) );
  OAI21_X1 U88339 ( .B1(n106341), .B2(n81318), .A(n98779), .ZN(
        \DLX_Datapath/RegisterFile/N22655 ) );
  AOI22_X1 U88340 ( .A1(n106061), .A2(n106339), .B1(n106336), .B2(n110409), 
        .ZN(n98779) );
  AND2_X2 U88341 ( .A1(stackBus_In[116]), .A2(n105203), .ZN(n81472) );
  OAI21_X1 U88342 ( .B1(n80185), .B2(n106162), .A(n98780), .ZN(
        \DLX_Datapath/RegisterFile/N22654 ) );
  AOI22_X1 U88343 ( .A1(n81347), .A2(n106340), .B1(n106336), .B2(n110087), 
        .ZN(n98780) );
  AND2_X2 U88344 ( .A1(stackBus_In[115]), .A2(n105203), .ZN(n81347) );
  OAI21_X1 U88345 ( .B1(n80185), .B2(n106106), .A(n98781), .ZN(
        \DLX_Datapath/RegisterFile/N22653 ) );
  AOI22_X1 U88346 ( .A1(n94527), .A2(n106338), .B1(n106336), .B2(n110194), 
        .ZN(n98781) );
  AND2_X2 U88347 ( .A1(stackBus_In[114]), .A2(n105203), .ZN(n94527) );
  OAI21_X1 U88348 ( .B1(n80185), .B2(n106219), .A(n98782), .ZN(
        \DLX_Datapath/RegisterFile/N22652 ) );
  AOI22_X1 U88349 ( .A1(n81297), .A2(n106339), .B1(n106336), .B2(n109979), 
        .ZN(n98782) );
  AND2_X2 U88350 ( .A1(stackBus_In[113]), .A2(n105202), .ZN(n81297) );
  OAI21_X1 U88351 ( .B1(n106341), .B2(n81398), .A(n98783), .ZN(
        \DLX_Datapath/RegisterFile/N22651 ) );
  AOI22_X1 U88352 ( .A1(n94530), .A2(n106338), .B1(n106336), .B2(n109862), 
        .ZN(n98783) );
  AND2_X2 U88353 ( .A1(stackBus_In[112]), .A2(n105203), .ZN(n94530) );
  OAI21_X1 U88354 ( .B1(n80185), .B2(n106233), .A(n98784), .ZN(
        \DLX_Datapath/RegisterFile/N22650 ) );
  AOI22_X1 U88355 ( .A1(n81286), .A2(n106340), .B1(n106336), .B2(n108236), 
        .ZN(n98784) );
  AND2_X2 U88356 ( .A1(stackBus_In[111]), .A2(n105202), .ZN(n81286) );
  OAI21_X1 U88357 ( .B1(n80185), .B2(n106171), .A(n98785), .ZN(
        \DLX_Datapath/RegisterFile/N22649 ) );
  AOI22_X1 U88358 ( .A1(n106168), .A2(n106338), .B1(n106336), .B2(n108359), 
        .ZN(n98785) );
  AND2_X2 U88359 ( .A1(stackBus_In[110]), .A2(n105203), .ZN(n81342) );
  OAI21_X1 U88360 ( .B1(n106341), .B2(n81281), .A(n98786), .ZN(
        \DLX_Datapath/RegisterFile/N22648 ) );
  AOI22_X1 U88361 ( .A1(n81283), .A2(n106339), .B1(n106336), .B2(n108470), 
        .ZN(n98786) );
  AND2_X2 U88362 ( .A1(stackBus_In[109]), .A2(n105202), .ZN(n81283) );
  OAI21_X1 U88363 ( .B1(n80185), .B2(n106070), .A(n98787), .ZN(
        \DLX_Datapath/RegisterFile/N22647 ) );
  AOI22_X1 U88364 ( .A1(n81453), .A2(n106340), .B1(n106335), .B2(n107708), 
        .ZN(n98787) );
  AND2_X2 U88365 ( .A1(stackBus_In[108]), .A2(n105202), .ZN(n81453) );
  OAI21_X1 U88366 ( .B1(n106341), .B2(n106197), .A(n98788), .ZN(
        \DLX_Datapath/RegisterFile/N22646 ) );
  AOI22_X1 U88367 ( .A1(n105626), .A2(n106340), .B1(n106335), .B2(n109623), 
        .ZN(n98788) );
  AND2_X2 U88368 ( .A1(stackBus_In[107]), .A2(n105202), .ZN(n94536) );
  OAI21_X1 U88369 ( .B1(n106341), .B2(n106245), .A(n98789), .ZN(
        \DLX_Datapath/RegisterFile/N22645 ) );
  AOI22_X1 U88370 ( .A1(n106241), .A2(n106340), .B1(n106335), .B2(n108585), 
        .ZN(n98789) );
  AND2_X2 U88371 ( .A1(stackBus_In[106]), .A2(n105202), .ZN(n81280) );
  OAI21_X1 U88372 ( .B1(n106341), .B2(n106158), .A(n98790), .ZN(
        \DLX_Datapath/RegisterFile/N22644 ) );
  AOI22_X1 U88373 ( .A1(n81351), .A2(n106339), .B1(n106335), .B2(n109730), 
        .ZN(n98790) );
  AND2_X2 U88374 ( .A1(stackBus_In[105]), .A2(n105201), .ZN(n81351) );
  OAI21_X1 U88375 ( .B1(n80185), .B2(n106113), .A(n98791), .ZN(
        \DLX_Datapath/RegisterFile/N22643 ) );
  AOI22_X1 U88376 ( .A1(n106019), .A2(n106340), .B1(n106335), .B2(n109515), 
        .ZN(n98791) );
  AND2_X2 U88377 ( .A1(stackBus_In[104]), .A2(n105202), .ZN(n81567) );
  OAI21_X1 U88378 ( .B1(n106341), .B2(n106007), .A(n98792), .ZN(
        \DLX_Datapath/RegisterFile/N22642 ) );
  AOI22_X1 U88379 ( .A1(n94541), .A2(n106339), .B1(n106335), .B2(n109052), 
        .ZN(n98792) );
  AND2_X2 U88380 ( .A1(stackBus_In[103]), .A2(n105202), .ZN(n94541) );
  OAI21_X1 U88381 ( .B1(n106341), .B2(n81267), .A(n98793), .ZN(
        \DLX_Datapath/RegisterFile/N22641 ) );
  AOI22_X1 U88382 ( .A1(n81269), .A2(n106340), .B1(n106335), .B2(n109400), 
        .ZN(n98793) );
  AND2_X2 U88383 ( .A1(stackBus_In[102]), .A2(n105202), .ZN(n81269) );
  OAI21_X1 U88384 ( .B1(n106341), .B2(n81509), .A(n98794), .ZN(
        \DLX_Datapath/RegisterFile/N22640 ) );
  AOI22_X1 U88385 ( .A1(n105623), .A2(n106340), .B1(n106335), .B2(n109281), 
        .ZN(n98794) );
  AND2_X2 U88386 ( .A1(stackBus_In[101]), .A2(n105202), .ZN(n94544) );
  OAI21_X1 U88387 ( .B1(n106341), .B2(n81501), .A(n98795), .ZN(
        \DLX_Datapath/RegisterFile/N22639 ) );
  AOI22_X1 U88388 ( .A1(n105622), .A2(n106340), .B1(n106335), .B2(n109173), 
        .ZN(n98795) );
  AND2_X2 U88389 ( .A1(stackBus_In[100]), .A2(n105202), .ZN(n94546) );
  OAI21_X1 U88390 ( .B1(n106341), .B2(n81415), .A(n98796), .ZN(
        \DLX_Datapath/RegisterFile/N22638 ) );
  AOI22_X1 U88391 ( .A1(n105621), .A2(n106339), .B1(n106335), .B2(n108708), 
        .ZN(n98796) );
  AND2_X2 U88392 ( .A1(stackBus_In[99]), .A2(n105201), .ZN(n94548) );
  OAI21_X1 U88393 ( .B1(n106341), .B2(n81498), .A(n98797), .ZN(
        \DLX_Datapath/RegisterFile/N22637 ) );
  AOI22_X1 U88394 ( .A1(n105911), .A2(n106339), .B1(n106335), .B2(n108936), 
        .ZN(n98797) );
  AND2_X2 U88395 ( .A1(stackBus_In[98]), .A2(n105202), .ZN(n81783) );
  OAI21_X1 U88396 ( .B1(n106341), .B2(n81262), .A(n98798), .ZN(
        \DLX_Datapath/RegisterFile/N22635 ) );
  AOI22_X1 U88397 ( .A1(n81265), .A2(n106339), .B1(n106335), .B2(n107363), 
        .ZN(n98798) );
  AOI21_X1 U88398 ( .B1(n98799), .B2(n105602), .A(n98800), .ZN(n80189) );
  OAI21_X1 U88399 ( .B1(n95131), .B2(n96489), .A(n107022), .ZN(n98799) );
  OR2_X1 U88401 ( .A1(n98800), .A2(n96489), .ZN(n98801) );
  NOR2_X1 U88402 ( .A1(n105089), .A2(n80185), .ZN(n98800) );
  AND2_X2 U88403 ( .A1(stackBus_In[96]), .A2(n105201), .ZN(n81265) );
  NAND2_X1 U88404 ( .A1(n98654), .A2(n94399), .ZN(n80185) );
  NOR2_X1 U88405 ( .A1(n98501), .A2(n104762), .ZN(n94399) );
  OR2_X1 U88406 ( .A1(n98655), .A2(n90127), .ZN(n98501) );
  NAND2_X1 U88407 ( .A1(n90120), .A2(n90119), .ZN(n98655) );
  OAI21_X1 U88408 ( .B1(n81358), .B2(n104492), .A(n98803), .ZN(
        \DLX_Datapath/RegisterFile/N22634 ) );
  AOI22_X1 U88409 ( .A1(n105233), .A2(n94559), .B1(n105194), .B2(n107919), 
        .ZN(n98803) );
  AND2_X2 U88410 ( .A1(stackBus_In[95]), .A2(n105201), .ZN(n94559) );
  OAI21_X1 U88411 ( .B1(n105969), .B2(n98802), .A(n98805), .ZN(
        \DLX_Datapath/RegisterFile/N22633 ) );
  AOI22_X1 U88412 ( .A1(n98804), .A2(n94562), .B1(n105194), .B2(n108016), .ZN(
        n98805) );
  AND2_X2 U88413 ( .A1(stackBus_In[94]), .A2(n105201), .ZN(n94562) );
  OAI21_X1 U88414 ( .B1(n81378), .B2(n104492), .A(n98806), .ZN(
        \DLX_Datapath/RegisterFile/N22632 ) );
  AOI22_X1 U88415 ( .A1(n98804), .A2(n94564), .B1(n105194), .B2(n107286), .ZN(
        n98806) );
  AND2_X2 U88416 ( .A1(stackBus_In[93]), .A2(n105201), .ZN(n94564) );
  OAI21_X1 U88417 ( .B1(n106211), .B2(n104492), .A(n98807), .ZN(
        \DLX_Datapath/RegisterFile/N22631 ) );
  AOI22_X1 U88418 ( .A1(n98804), .A2(n94566), .B1(n105194), .B2(n107824), .ZN(
        n98807) );
  AND2_X2 U88419 ( .A1(stackBus_In[92]), .A2(n105201), .ZN(n94566) );
  OAI21_X1 U88420 ( .B1(n106206), .B2(n104492), .A(n98808), .ZN(
        \DLX_Datapath/RegisterFile/N22630 ) );
  AOI22_X1 U88421 ( .A1(n98804), .A2(n94568), .B1(n105194), .B2(n110720), .ZN(
        n98808) );
  AND2_X2 U88422 ( .A1(stackBus_In[91]), .A2(n105201), .ZN(n94568) );
  OAI21_X1 U88423 ( .B1(n81408), .B2(n98802), .A(n98809), .ZN(
        \DLX_Datapath/RegisterFile/N22629 ) );
  AOI22_X1 U88424 ( .A1(n98804), .A2(n94570), .B1(n105194), .B2(n108123), .ZN(
        n98809) );
  AND2_X2 U88425 ( .A1(stackBus_In[90]), .A2(n105201), .ZN(n94570) );
  OAI21_X1 U88426 ( .B1(n106257), .B2(n104492), .A(n98810), .ZN(
        \DLX_Datapath/RegisterFile/N22628 ) );
  AOI22_X1 U88427 ( .A1(n98804), .A2(n94572), .B1(n105194), .B2(n110822), .ZN(
        n98810) );
  AND2_X2 U88428 ( .A1(stackBus_In[89]), .A2(n105201), .ZN(n94572) );
  OAI21_X1 U88429 ( .B1(n105990), .B2(n104492), .A(n98811), .ZN(
        \DLX_Datapath/RegisterFile/N22627 ) );
  AOI22_X1 U88430 ( .A1(n98804), .A2(n94574), .B1(n105193), .B2(n110923), .ZN(
        n98811) );
  AND2_X2 U88431 ( .A1(stackBus_In[88]), .A2(n105201), .ZN(n94574) );
  OAI21_X1 U88432 ( .B1(n80190), .B2(n104492), .A(n98812), .ZN(
        \DLX_Datapath/RegisterFile/N22626 ) );
  AOI22_X1 U88433 ( .A1(n105234), .A2(n94576), .B1(n105193), .B2(n110517), 
        .ZN(n98812) );
  AND2_X2 U88434 ( .A1(stackBus_In[87]), .A2(n105201), .ZN(n94576) );
  OAI21_X1 U88435 ( .B1(n106193), .B2(n104492), .A(n98813), .ZN(
        \DLX_Datapath/RegisterFile/N22625 ) );
  AOI22_X1 U88436 ( .A1(n105234), .A2(n94578), .B1(n105193), .B2(n110301), 
        .ZN(n98813) );
  AND2_X2 U88437 ( .A1(stackBus_In[86]), .A2(n105200), .ZN(n94578) );
  OAI21_X1 U88438 ( .B1(n81383), .B2(n104492), .A(n98814), .ZN(
        \DLX_Datapath/RegisterFile/N22624 ) );
  AOI22_X1 U88439 ( .A1(n105234), .A2(n94580), .B1(n105193), .B2(n110622), 
        .ZN(n98814) );
  AND2_X2 U88440 ( .A1(stackBus_In[85]), .A2(n105200), .ZN(n94580) );
  OAI21_X1 U88441 ( .B1(n106188), .B2(n104492), .A(n98815), .ZN(
        \DLX_Datapath/RegisterFile/N22623 ) );
  AOI22_X1 U88442 ( .A1(n105234), .A2(n94582), .B1(n105193), .B2(n110410), 
        .ZN(n98815) );
  AND2_X2 U88443 ( .A1(stackBus_In[84]), .A2(n105200), .ZN(n94582) );
  OAI21_X1 U88444 ( .B1(n81345), .B2(n104492), .A(n98816), .ZN(
        \DLX_Datapath/RegisterFile/N22622 ) );
  AOI22_X1 U88445 ( .A1(n105234), .A2(n94584), .B1(n105193), .B2(n110088), 
        .ZN(n98816) );
  AND2_X2 U88446 ( .A1(stackBus_In[83]), .A2(n105200), .ZN(n94584) );
  OAI21_X1 U88447 ( .B1(n81403), .B2(n104492), .A(n98817), .ZN(
        \DLX_Datapath/RegisterFile/N22621 ) );
  AOI22_X1 U88448 ( .A1(n105234), .A2(n94586), .B1(n105193), .B2(n110195), 
        .ZN(n98817) );
  AND2_X2 U88449 ( .A1(stackBus_In[82]), .A2(n105200), .ZN(n94586) );
  OAI21_X1 U88450 ( .B1(n106221), .B2(n104492), .A(n98818), .ZN(
        \DLX_Datapath/RegisterFile/N22620 ) );
  AOI22_X1 U88451 ( .A1(n105234), .A2(n94588), .B1(n105193), .B2(n109980), 
        .ZN(n98818) );
  AND2_X2 U88452 ( .A1(stackBus_In[81]), .A2(n105200), .ZN(n94588) );
  OAI21_X1 U88453 ( .B1(n81398), .B2(n104492), .A(n98819), .ZN(
        \DLX_Datapath/RegisterFile/N22619 ) );
  AOI22_X1 U88454 ( .A1(n105234), .A2(n94590), .B1(n105193), .B2(n109863), 
        .ZN(n98819) );
  AND2_X2 U88455 ( .A1(stackBus_In[80]), .A2(n105200), .ZN(n94590) );
  OAI21_X1 U88456 ( .B1(n106233), .B2(n98802), .A(n98820), .ZN(
        \DLX_Datapath/RegisterFile/N22618 ) );
  AOI22_X1 U88457 ( .A1(n105234), .A2(n94592), .B1(n105193), .B2(n108237), 
        .ZN(n98820) );
  AND2_X2 U88458 ( .A1(stackBus_In[79]), .A2(n105200), .ZN(n94592) );
  OAI21_X1 U88459 ( .B1(n81340), .B2(n104492), .A(n98821), .ZN(
        \DLX_Datapath/RegisterFile/N22617 ) );
  AOI22_X1 U88460 ( .A1(n105234), .A2(n94594), .B1(n105193), .B2(n108360), 
        .ZN(n98821) );
  AND2_X2 U88461 ( .A1(stackBus_In[78]), .A2(n105200), .ZN(n94594) );
  OAI21_X1 U88462 ( .B1(n106236), .B2(n104492), .A(n98822), .ZN(
        \DLX_Datapath/RegisterFile/N22616 ) );
  AOI22_X1 U88463 ( .A1(n105234), .A2(n94596), .B1(n105193), .B2(n108471), 
        .ZN(n98822) );
  AND2_X2 U88464 ( .A1(stackBus_In[77]), .A2(n105200), .ZN(n94596) );
  OAI21_X1 U88465 ( .B1(n81451), .B2(n104492), .A(n98823), .ZN(
        \DLX_Datapath/RegisterFile/N22615 ) );
  AOI22_X1 U88466 ( .A1(n105233), .A2(n94598), .B1(n105192), .B2(n107709), 
        .ZN(n98823) );
  AND2_X2 U88467 ( .A1(stackBus_In[76]), .A2(n105200), .ZN(n94598) );
  OAI21_X1 U88468 ( .B1(n106200), .B2(n104492), .A(n98824), .ZN(
        \DLX_Datapath/RegisterFile/N22614 ) );
  AOI22_X1 U88469 ( .A1(n105233), .A2(n94600), .B1(n105192), .B2(n109624), 
        .ZN(n98824) );
  AND2_X2 U88470 ( .A1(stackBus_In[75]), .A2(n105200), .ZN(n94600) );
  OAI21_X1 U88471 ( .B1(n106246), .B2(n104492), .A(n98825), .ZN(
        \DLX_Datapath/RegisterFile/N22613 ) );
  AOI22_X1 U88472 ( .A1(n105233), .A2(n94602), .B1(n105192), .B2(n108586), 
        .ZN(n98825) );
  AND2_X2 U88473 ( .A1(stackBus_In[74]), .A2(n105200), .ZN(n94602) );
  OAI21_X1 U88474 ( .B1(n81349), .B2(n104492), .A(n98826), .ZN(
        \DLX_Datapath/RegisterFile/N22612 ) );
  AOI22_X1 U88475 ( .A1(n105233), .A2(n94604), .B1(n105192), .B2(n109731), 
        .ZN(n98826) );
  AND2_X2 U88476 ( .A1(stackBus_In[73]), .A2(n105201), .ZN(n94604) );
  OAI21_X1 U88477 ( .B1(n81394), .B2(n98802), .A(n98827), .ZN(
        \DLX_Datapath/RegisterFile/N22611 ) );
  AOI22_X1 U88478 ( .A1(n105233), .A2(n94606), .B1(n105192), .B2(n109516), 
        .ZN(n98827) );
  AND2_X2 U88479 ( .A1(stackBus_In[72]), .A2(n105203), .ZN(n94606) );
  OAI21_X1 U88480 ( .B1(n101624), .B2(n98828), .A(n98829), .ZN(
        \DLX_Datapath/RegisterFile/N22610 ) );
  AOI22_X1 U88481 ( .A1(n105235), .A2(n106012), .B1(n98804), .B2(n94608), .ZN(
        n98829) );
  AND2_X2 U88482 ( .A1(stackBus_In[71]), .A2(n105201), .ZN(n94608) );
  NAND2_X1 U88483 ( .A1(n105502), .A2(n89271), .ZN(n81588) );
  OAI21_X1 U88484 ( .B1(n111064), .B2(n108975), .A(n98830), .ZN(n89271) );
  AOI22_X1 U88485 ( .A1(n98831), .A2(n69730), .B1(n98832), .B2(n111088), .ZN(
        n98830) );
  OAI21_X1 U88486 ( .B1(n106260), .B2(n104492), .A(n98833), .ZN(
        \DLX_Datapath/RegisterFile/N22609 ) );
  AOI22_X1 U88487 ( .A1(n105233), .A2(n94610), .B1(n105192), .B2(n109401), 
        .ZN(n98833) );
  AND2_X2 U88488 ( .A1(stackBus_In[70]), .A2(n105202), .ZN(n94610) );
  OAI21_X1 U88489 ( .B1(n106045), .B2(n104492), .A(n98834), .ZN(
        \DLX_Datapath/RegisterFile/N22608 ) );
  AOI22_X1 U88490 ( .A1(n105233), .A2(n94612), .B1(n105192), .B2(n109282), 
        .ZN(n98834) );
  AND2_X2 U88491 ( .A1(stackBus_In[69]), .A2(n105200), .ZN(n94612) );
  OAI21_X1 U88492 ( .B1(n106050), .B2(n104492), .A(n98835), .ZN(
        \DLX_Datapath/RegisterFile/N22607 ) );
  AOI22_X1 U88493 ( .A1(n105233), .A2(n94614), .B1(n105192), .B2(n109174), 
        .ZN(n98835) );
  AND2_X2 U88494 ( .A1(stackBus_In[68]), .A2(n105203), .ZN(n94614) );
  OAI21_X1 U88495 ( .B1(n81415), .B2(n104492), .A(n98836), .ZN(
        \DLX_Datapath/RegisterFile/N22606 ) );
  AOI22_X1 U88496 ( .A1(n105233), .A2(n94616), .B1(n105192), .B2(n108709), 
        .ZN(n98836) );
  AND2_X2 U88497 ( .A1(stackBus_In[67]), .A2(n107022), .ZN(n94616) );
  OAI21_X1 U88498 ( .B1(n106056), .B2(n104492), .A(n98837), .ZN(
        \DLX_Datapath/RegisterFile/N22605 ) );
  AOI22_X1 U88499 ( .A1(n105233), .A2(n94618), .B1(n105192), .B2(n108937), 
        .ZN(n98837) );
  AND2_X2 U88500 ( .A1(stackBus_In[66]), .A2(n105202), .ZN(n94618) );
  OAI21_X1 U88501 ( .B1(n105215), .B2(n104492), .A(n98838), .ZN(
        \DLX_Datapath/RegisterFile/N22604 ) );
  AOI22_X1 U88502 ( .A1(n105233), .A2(n94620), .B1(n105192), .B2(n108825), 
        .ZN(n98838) );
  AND2_X2 U88503 ( .A1(stackBus_In[65]), .A2(n107022), .ZN(n94620) );
  OAI21_X1 U88504 ( .B1(n106268), .B2(n98802), .A(n98839), .ZN(
        \DLX_Datapath/RegisterFile/N22603 ) );
  AOI22_X1 U88505 ( .A1(n105234), .A2(n94622), .B1(n105192), .B2(n107364), 
        .ZN(n98839) );
  NAND2_X1 U88506 ( .A1(n98840), .A2(n98841), .ZN(n98828) );
  AND2_X2 U88507 ( .A1(stackBus_In[64]), .A2(n105205), .ZN(n94622) );
  AND2_X2 U88508 ( .A1(n98842), .A2(n98841), .ZN(n98804) );
  NAND2_X1 U88509 ( .A1(n105235), .A2(n105502), .ZN(n98841) );
  NAND2_X1 U88510 ( .A1(n94434), .A2(n98654), .ZN(n98802) );
  NOR2_X1 U88511 ( .A1(n98539), .A2(n104762), .ZN(n94434) );
  OR2_X1 U88512 ( .A1(n98843), .A2(n90120), .ZN(n98539) );
  NAND2_X1 U88513 ( .A1(n90119), .A2(n107123), .ZN(n98843) );
  OAI21_X1 U88514 ( .B1(n106146), .B2(n105901), .A(n98844), .ZN(
        \DLX_Datapath/RegisterFile/N22602 ) );
  AOI22_X1 U88515 ( .A1(n81797), .A2(n81521), .B1(n106759), .B2(n107920), .ZN(
        n98844) );
  AND2_X2 U88516 ( .A1(stackBus_In[63]), .A2(n105200), .ZN(n81521) );
  OAI21_X1 U88517 ( .B1(n105968), .B2(n105902), .A(n98845), .ZN(
        \DLX_Datapath/RegisterFile/N22601 ) );
  AOI22_X1 U88518 ( .A1(n81797), .A2(n81653), .B1(n70535), .B2(n106759), .ZN(
        n98845) );
  AND2_X2 U88519 ( .A1(stackBus_In[62]), .A2(n105200), .ZN(n81653) );
  OAI21_X1 U88520 ( .B1(n81378), .B2(n105901), .A(n98846), .ZN(
        \DLX_Datapath/RegisterFile/N22600 ) );
  AOI22_X1 U88521 ( .A1(n81797), .A2(n81380), .B1(n69588), .B2(n105191), .ZN(
        n98846) );
  AND2_X2 U88522 ( .A1(stackBus_In[61]), .A2(n105201), .ZN(n81380) );
  OAI21_X1 U88523 ( .B1(n81299), .B2(n105902), .A(n98847), .ZN(
        \DLX_Datapath/RegisterFile/N22599 ) );
  AOI22_X1 U88524 ( .A1(n81797), .A2(n81377), .B1(n70249), .B2(n105191), .ZN(
        n98847) );
  AND2_X2 U88525 ( .A1(stackBus_In[60]), .A2(n105202), .ZN(n81377) );
  OAI21_X1 U88526 ( .B1(n81306), .B2(n105901), .A(n98848), .ZN(
        \DLX_Datapath/RegisterFile/N22598 ) );
  AOI22_X1 U88527 ( .A1(n81797), .A2(n81428), .B1(n74095), .B2(n105191), .ZN(
        n98848) );
  AND2_X2 U88528 ( .A1(stackBus_In[59]), .A2(n105203), .ZN(n81428) );
  OAI21_X1 U88529 ( .B1(n81408), .B2(n105902), .A(n98849), .ZN(
        \DLX_Datapath/RegisterFile/N22597 ) );
  AOI22_X1 U88530 ( .A1(n81797), .A2(n81410), .B1(n106759), .B2(n108124), .ZN(
        n98849) );
  AND2_X2 U88531 ( .A1(stackBus_In[58]), .A2(n105203), .ZN(n81410) );
  OAI21_X1 U88532 ( .B1(n106254), .B2(n105902), .A(n98850), .ZN(
        \DLX_Datapath/RegisterFile/N22596 ) );
  AOI22_X1 U88533 ( .A1(n81797), .A2(n81700), .B1(n106759), .B2(n110823), .ZN(
        n98850) );
  AND2_X2 U88534 ( .A1(stackBus_In[57]), .A2(n105201), .ZN(n81700) );
  OAI21_X1 U88535 ( .B1(n105990), .B2(n105902), .A(n98851), .ZN(
        \DLX_Datapath/RegisterFile/N22595 ) );
  AOI22_X1 U88536 ( .A1(n81797), .A2(n81632), .B1(n106759), .B2(n110924), .ZN(
        n98851) );
  AND2_X2 U88537 ( .A1(stackBus_In[56]), .A2(n105201), .ZN(n81632) );
  OAI21_X1 U88538 ( .B1(n80190), .B2(n105902), .A(n98852), .ZN(
        \DLX_Datapath/RegisterFile/N22594 ) );
  AOI22_X1 U88539 ( .A1(n81797), .A2(n81414), .B1(n73812), .B2(n105191), .ZN(
        n98852) );
  AND2_X2 U88540 ( .A1(stackBus_In[55]), .A2(n105203), .ZN(n81414) );
  OAI21_X1 U88541 ( .B1(n81315), .B2(n105902), .A(n98853), .ZN(
        \DLX_Datapath/RegisterFile/N22593 ) );
  AOI22_X1 U88542 ( .A1(n81797), .A2(n81317), .B1(n106759), .B2(n110302), .ZN(
        n98853) );
  AND2_X2 U88543 ( .A1(stackBus_In[54]), .A2(n105200), .ZN(n81317) );
  OAI21_X1 U88544 ( .B1(n106129), .B2(n105902), .A(n98854), .ZN(
        \DLX_Datapath/RegisterFile/N22592 ) );
  AOI22_X1 U88545 ( .A1(n81797), .A2(n81386), .B1(n73953), .B2(n106759), .ZN(
        n98854) );
  AND2_X2 U88546 ( .A1(stackBus_In[53]), .A2(n105202), .ZN(n81386) );
  OAI21_X1 U88547 ( .B1(n81318), .B2(n105902), .A(n98855), .ZN(
        \DLX_Datapath/RegisterFile/N22591 ) );
  AOI22_X1 U88548 ( .A1(n81797), .A2(n81320), .B1(n105190), .B2(n110411), .ZN(
        n98855) );
  AND2_X2 U88549 ( .A1(stackBus_In[52]), .A2(n105201), .ZN(n81320) );
  OAI21_X1 U88550 ( .B1(n106165), .B2(n105902), .A(n98856), .ZN(
        \DLX_Datapath/RegisterFile/N22590 ) );
  AOI22_X1 U88551 ( .A1(n81797), .A2(n81604), .B1(n105190), .B2(n110089), .ZN(
        n98856) );
  AND2_X2 U88552 ( .A1(stackBus_In[51]), .A2(n105202), .ZN(n81604) );
  OAI21_X1 U88553 ( .B1(n106103), .B2(n105902), .A(n98857), .ZN(
        \DLX_Datapath/RegisterFile/N22589 ) );
  AOI22_X1 U88554 ( .A1(n81797), .A2(n81405), .B1(n105190), .B2(n110196), .ZN(
        n98857) );
  AND2_X2 U88555 ( .A1(stackBus_In[50]), .A2(n105201), .ZN(n81405) );
  OAI21_X1 U88556 ( .B1(n81294), .B2(n105902), .A(n98858), .ZN(
        \DLX_Datapath/RegisterFile/N22588 ) );
  AOI22_X1 U88557 ( .A1(n81797), .A2(n81402), .B1(n105190), .B2(n109981), .ZN(
        n98858) );
  AND2_X2 U88558 ( .A1(stackBus_In[49]), .A2(n105203), .ZN(n81402) );
  OAI21_X1 U88559 ( .B1(n106111), .B2(n105902), .A(n98859), .ZN(
        \DLX_Datapath/RegisterFile/N22587 ) );
  AOI22_X1 U88560 ( .A1(n81797), .A2(n81400), .B1(n105190), .B2(n109864), .ZN(
        n98859) );
  AND2_X2 U88561 ( .A1(stackBus_In[48]), .A2(n105202), .ZN(n81400) );
  OAI21_X1 U88562 ( .B1(n81284), .B2(n105902), .A(n98860), .ZN(
        \DLX_Datapath/RegisterFile/N22586 ) );
  AOI22_X1 U88563 ( .A1(n81797), .A2(n81332), .B1(n105190), .B2(n108238), .ZN(
        n98860) );
  AND2_X2 U88564 ( .A1(stackBus_In[47]), .A2(n105201), .ZN(n81332) );
  OAI21_X1 U88565 ( .B1(n81340), .B2(n105902), .A(n98861), .ZN(
        \DLX_Datapath/RegisterFile/N22585 ) );
  AOI22_X1 U88566 ( .A1(n81797), .A2(n81373), .B1(n105190), .B2(n108361), .ZN(
        n98861) );
  AND2_X2 U88567 ( .A1(stackBus_In[46]), .A2(n105201), .ZN(n81373) );
  OAI21_X1 U88568 ( .B1(n106235), .B2(n105901), .A(n98862), .ZN(
        \DLX_Datapath/RegisterFile/N22584 ) );
  AOI22_X1 U88569 ( .A1(n81797), .A2(n81322), .B1(n105190), .B2(n108472), .ZN(
        n98862) );
  AND2_X2 U88570 ( .A1(stackBus_In[45]), .A2(n105203), .ZN(n81322) );
  OAI21_X1 U88571 ( .B1(n81451), .B2(n105901), .A(n98863), .ZN(
        \DLX_Datapath/RegisterFile/N22583 ) );
  AOI22_X1 U88572 ( .A1(n81797), .A2(n81506), .B1(n105190), .B2(n107710), .ZN(
        n98863) );
  AND2_X2 U88573 ( .A1(stackBus_In[44]), .A2(n105200), .ZN(n81506) );
  OAI21_X1 U88574 ( .B1(n81310), .B2(n105901), .A(n98864), .ZN(
        \DLX_Datapath/RegisterFile/N22582 ) );
  AOI22_X1 U88575 ( .A1(n81797), .A2(n81313), .B1(n105190), .B2(n109625), .ZN(
        n98864) );
  AND2_X2 U88576 ( .A1(stackBus_In[43]), .A2(n105200), .ZN(n81313) );
  OAI21_X1 U88577 ( .B1(n81278), .B2(n105901), .A(n98865), .ZN(
        \DLX_Datapath/RegisterFile/N22581 ) );
  AOI22_X1 U88578 ( .A1(n81797), .A2(n81330), .B1(n105190), .B2(n108587), .ZN(
        n98865) );
  AND2_X2 U88579 ( .A1(stackBus_In[42]), .A2(n105199), .ZN(n81330) );
  OAI21_X1 U88580 ( .B1(n106160), .B2(n105901), .A(n98866), .ZN(
        \DLX_Datapath/RegisterFile/N22580 ) );
  AOI22_X1 U88581 ( .A1(n81797), .A2(n81425), .B1(n105191), .B2(n109732), .ZN(
        n98866) );
  AND2_X2 U88582 ( .A1(stackBus_In[41]), .A2(n105201), .ZN(n81425) );
  OAI21_X1 U88583 ( .B1(n106115), .B2(n105901), .A(n98867), .ZN(
        \DLX_Datapath/RegisterFile/N22579 ) );
  AOI22_X1 U88584 ( .A1(n81797), .A2(n81396), .B1(n105191), .B2(n109517), .ZN(
        n98867) );
  AND2_X2 U88585 ( .A1(stackBus_In[40]), .A2(n105202), .ZN(n81396) );
  OAI21_X1 U88586 ( .B1(n81267), .B2(n105901), .A(n98868), .ZN(
        \DLX_Datapath/RegisterFile/N22577 ) );
  AOI22_X1 U88587 ( .A1(n81797), .A2(n81423), .B1(n105191), .B2(n109402), .ZN(
        n98868) );
  AND2_X2 U88588 ( .A1(stackBus_In[38]), .A2(n105205), .ZN(n81423) );
  OAI21_X1 U88589 ( .B1(n106043), .B2(n105901), .A(n98869), .ZN(
        \DLX_Datapath/RegisterFile/N22576 ) );
  AOI22_X1 U88590 ( .A1(n81797), .A2(n81511), .B1(n105191), .B2(n109283), .ZN(
        n98869) );
  AND2_X2 U88591 ( .A1(stackBus_In[37]), .A2(n105202), .ZN(n81511) );
  OAI21_X1 U88592 ( .B1(n106049), .B2(n105901), .A(n98870), .ZN(
        \DLX_Datapath/RegisterFile/N22575 ) );
  AOI22_X1 U88593 ( .A1(n81797), .A2(n81503), .B1(n105191), .B2(n109175), .ZN(
        n98870) );
  AND2_X2 U88594 ( .A1(stackBus_In[36]), .A2(n105202), .ZN(n81503) );
  OAI21_X1 U88595 ( .B1(n106096), .B2(n105901), .A(n98871), .ZN(
        \DLX_Datapath/RegisterFile/N22574 ) );
  AOI22_X1 U88596 ( .A1(n81797), .A2(n81417), .B1(n105191), .B2(n108710), .ZN(
        n98871) );
  AND2_X2 U88597 ( .A1(stackBus_In[35]), .A2(n105203), .ZN(n81417) );
  OAI21_X1 U88598 ( .B1(n105215), .B2(n105901), .A(n98872), .ZN(
        \DLX_Datapath/RegisterFile/N22572 ) );
  AOI22_X1 U88599 ( .A1(n81797), .A2(n81335), .B1(n105191), .B2(n108826), .ZN(
        n98872) );
  AND2_X2 U88600 ( .A1(stackBus_In[33]), .A2(n105199), .ZN(n81335) );
  OAI21_X1 U88601 ( .B1(n106266), .B2(n105901), .A(n98873), .ZN(
        \DLX_Datapath/RegisterFile/N22571 ) );
  AOI22_X1 U88602 ( .A1(n81797), .A2(n81327), .B1(n106759), .B2(n107365), .ZN(
        n98873) );
  NAND2_X1 U88603 ( .A1(n98840), .A2(n98874), .ZN(n81798) );
  AND2_X2 U88604 ( .A1(stackBus_In[32]), .A2(n105200), .ZN(n81327) );
  AND2_X2 U88605 ( .A1(n98842), .A2(n98874), .ZN(n81797) );
  NAND2_X1 U88606 ( .A1(n105903), .A2(n105501), .ZN(n98874) );
  NAND2_X1 U88607 ( .A1(n98654), .A2(n95132), .ZN(n81795) );
  NOR2_X1 U88608 ( .A1(n94470), .A2(n104762), .ZN(n95132) );
  NAND2_X1 U88609 ( .A1(n98875), .A2(n107122), .ZN(n94470) );
  NOR2_X1 U88610 ( .A1(n107114), .A2(n90127), .ZN(n98875) );
  OAI21_X1 U88611 ( .B1(n107921), .B2(n81256), .A(n98876), .ZN(
        \DLX_Datapath/RegisterFile/N22570 ) );
  AOI22_X1 U88612 ( .A1(n94667), .A2(n81258), .B1(n106150), .B2(n106273), .ZN(
        n98876) );
  NAND2_X1 U88613 ( .A1(n105501), .A2(n86303), .ZN(n81358) );
  OAI21_X1 U88614 ( .B1(n111064), .B2(n107749), .A(n98877), .ZN(n86303) );
  AOI22_X1 U88615 ( .A1(n98831), .A2(n69708), .B1(n98832), .B2(n111069), .ZN(
        n98877) );
  AND2_X2 U88616 ( .A1(stackBus_In[31]), .A2(n105202), .ZN(n94667) );
  OAI21_X1 U88617 ( .B1(n108017), .B2(n81256), .A(n98878), .ZN(
        \DLX_Datapath/RegisterFile/N22569 ) );
  AOI22_X1 U88618 ( .A1(n94670), .A2(n81258), .B1(n105972), .B2(n81260), .ZN(
        n98878) );
  NAND2_X1 U88619 ( .A1(n105501), .A2(n86558), .ZN(n81651) );
  OAI21_X1 U88620 ( .B1(n111064), .B2(n107750), .A(n98879), .ZN(n86558) );
  AOI22_X1 U88621 ( .A1(n98831), .A2(n69709), .B1(n98832), .B2(n111090), .ZN(
        n98879) );
  AND2_X2 U88622 ( .A1(stackBus_In[30]), .A2(n105201), .ZN(n94670) );
  OAI21_X1 U88623 ( .B1(n107287), .B2(n81256), .A(n98880), .ZN(
        \DLX_Datapath/RegisterFile/N22568 ) );
  AOI22_X1 U88624 ( .A1(n94672), .A2(n81258), .B1(n106139), .B2(n106273), .ZN(
        n98880) );
  NAND2_X1 U88625 ( .A1(n105501), .A2(n86676), .ZN(n81378) );
  OAI21_X1 U88626 ( .B1(n111064), .B2(n106837), .A(n98881), .ZN(n86676) );
  AOI22_X1 U88627 ( .A1(n98831), .A2(n69710), .B1(n98832), .B2(n111070), .ZN(
        n98881) );
  AND2_X2 U88628 ( .A1(stackBus_In[29]), .A2(n105200), .ZN(n94672) );
  OAI21_X1 U88629 ( .B1(n107825), .B2(n81256), .A(n98882), .ZN(
        \DLX_Datapath/RegisterFile/N22567 ) );
  AOI22_X1 U88630 ( .A1(n94674), .A2(n81258), .B1(n106212), .B2(n81260), .ZN(
        n98882) );
  NAND2_X1 U88631 ( .A1(n105500), .A2(n86794), .ZN(n81299) );
  OAI21_X1 U88632 ( .B1(n111064), .B2(n107751), .A(n98883), .ZN(n86794) );
  AOI22_X1 U88633 ( .A1(n98831), .A2(n69711), .B1(n98832), .B2(n111091), .ZN(
        n98883) );
  AND2_X2 U88634 ( .A1(stackBus_In[28]), .A2(n105202), .ZN(n94674) );
  OAI21_X1 U88635 ( .B1(n110721), .B2(n81256), .A(n98884), .ZN(
        \DLX_Datapath/RegisterFile/N22566 ) );
  AOI22_X1 U88636 ( .A1(n94676), .A2(n81258), .B1(n106207), .B2(n106273), .ZN(
        n98884) );
  NAND2_X1 U88637 ( .A1(n105502), .A2(n86912), .ZN(n81306) );
  OAI21_X1 U88638 ( .B1(n111064), .B2(n110654), .A(n98885), .ZN(n86912) );
  AOI22_X1 U88639 ( .A1(n98831), .A2(n69712), .B1(n98832), .B2(n111092), .ZN(
        n98885) );
  AND2_X2 U88640 ( .A1(stackBus_In[27]), .A2(n105199), .ZN(n94676) );
  OAI21_X1 U88641 ( .B1(n108125), .B2(n81256), .A(n98886), .ZN(
        \DLX_Datapath/RegisterFile/N22565 ) );
  AOI22_X1 U88642 ( .A1(n94678), .A2(n81258), .B1(n106102), .B2(n81260), .ZN(
        n98886) );
  NAND2_X1 U88643 ( .A1(n105500), .A2(n87030), .ZN(n81408) );
  OAI21_X1 U88644 ( .B1(n111064), .B2(n108053), .A(n98887), .ZN(n87030) );
  AOI22_X1 U88645 ( .A1(n98831), .A2(n69713), .B1(n98832), .B2(n111093), .ZN(
        n98887) );
  AND2_X2 U88646 ( .A1(stackBus_In[26]), .A2(n105203), .ZN(n94678) );
  OAI21_X1 U88647 ( .B1(n110824), .B2(n81256), .A(n98888), .ZN(
        \DLX_Datapath/RegisterFile/N22564 ) );
  AOI22_X1 U88648 ( .A1(n94680), .A2(n81258), .B1(n106258), .B2(n106273), .ZN(
        n98888) );
  NAND2_X1 U88649 ( .A1(n105500), .A2(n87148), .ZN(n81270) );
  OAI21_X1 U88650 ( .B1(n111064), .B2(n110751), .A(n98889), .ZN(n87148) );
  AOI22_X1 U88651 ( .A1(n98831), .A2(n69714), .B1(n98832), .B2(n111094), .ZN(
        n98889) );
  AND2_X2 U88652 ( .A1(stackBus_In[25]), .A2(n105205), .ZN(n94680) );
  OAI21_X1 U88653 ( .B1(n110925), .B2(n106274), .A(n98890), .ZN(
        \DLX_Datapath/RegisterFile/N22563 ) );
  AOI22_X1 U88654 ( .A1(n94682), .A2(n81258), .B1(n105993), .B2(n106273), .ZN(
        n98890) );
  NAND2_X1 U88655 ( .A1(n105501), .A2(n87266), .ZN(n81629) );
  OAI21_X1 U88656 ( .B1(n111064), .B2(n110852), .A(n98891), .ZN(n87266) );
  AOI22_X1 U88657 ( .A1(n105232), .A2(n69715), .B1(n98832), .B2(n111095), .ZN(
        n98891) );
  AND2_X2 U88658 ( .A1(stackBus_In[24]), .A2(n105199), .ZN(n94682) );
  OAI21_X1 U88659 ( .B1(n110518), .B2(n106274), .A(n98892), .ZN(
        \DLX_Datapath/RegisterFile/N22562 ) );
  AOI22_X1 U88660 ( .A1(n94684), .A2(n81258), .B1(n81260), .B2(n106334), .ZN(
        n98892) );
  NAND2_X1 U88661 ( .A1(n105502), .A2(n87384), .ZN(n80190) );
  OAI21_X1 U88662 ( .B1(n111064), .B2(n110447), .A(n98893), .ZN(n87384) );
  AOI22_X1 U88663 ( .A1(n98831), .A2(n69716), .B1(n98832), .B2(n111071), .ZN(
        n98893) );
  AND2_X2 U88664 ( .A1(stackBus_In[23]), .A2(n107022), .ZN(n94684) );
  OAI21_X1 U88665 ( .B1(n110303), .B2(n106274), .A(n98894), .ZN(
        \DLX_Datapath/RegisterFile/N22561 ) );
  AOI22_X1 U88666 ( .A1(n94686), .A2(n81258), .B1(n106194), .B2(n106273), .ZN(
        n98894) );
  NAND2_X1 U88667 ( .A1(n105500), .A2(n87502), .ZN(n81315) );
  OAI21_X1 U88668 ( .B1(n111064), .B2(n110230), .A(n98895), .ZN(n87502) );
  AOI22_X1 U88669 ( .A1(n105232), .A2(n69717), .B1(n98832), .B2(n111066), .ZN(
        n98895) );
  AND2_X2 U88670 ( .A1(stackBus_In[22]), .A2(n107022), .ZN(n94686) );
  OAI21_X1 U88671 ( .B1(n110623), .B2(n106274), .A(n98896), .ZN(
        \DLX_Datapath/RegisterFile/N22560 ) );
  AOI22_X1 U88672 ( .A1(n94688), .A2(n81258), .B1(n106132), .B2(n106273), .ZN(
        n98896) );
  NAND2_X1 U88673 ( .A1(n105500), .A2(n87620), .ZN(n81383) );
  OAI21_X1 U88674 ( .B1(n111064), .B2(n110547), .A(n98897), .ZN(n87620) );
  AOI22_X1 U88675 ( .A1(n105232), .A2(n69718), .B1(n98832), .B2(n111067), .ZN(
        n98897) );
  AND2_X2 U88676 ( .A1(stackBus_In[21]), .A2(n105203), .ZN(n94688) );
  OAI21_X1 U88677 ( .B1(n110412), .B2(n106274), .A(n98898), .ZN(
        \DLX_Datapath/RegisterFile/N22559 ) );
  AOI22_X1 U88678 ( .A1(n94690), .A2(n81258), .B1(n106189), .B2(n106273), .ZN(
        n98898) );
  NAND2_X1 U88679 ( .A1(n105500), .A2(n87738), .ZN(n81318) );
  OAI21_X1 U88680 ( .B1(n111064), .B2(n110338), .A(n98899), .ZN(n87738) );
  AOI22_X1 U88681 ( .A1(n98831), .A2(n69719), .B1(n98832), .B2(n111068), .ZN(
        n98899) );
  AND2_X2 U88682 ( .A1(stackBus_In[20]), .A2(n105205), .ZN(n94690) );
  OAI21_X1 U88683 ( .B1(n110090), .B2(n106274), .A(n98900), .ZN(
        \DLX_Datapath/RegisterFile/N22558 ) );
  AOI22_X1 U88684 ( .A1(n94692), .A2(n81258), .B1(n106166), .B2(n106273), .ZN(
        n98900) );
  NAND2_X1 U88685 ( .A1(n105500), .A2(n87856), .ZN(n81345) );
  OAI21_X1 U88686 ( .B1(n111064), .B2(n110012), .A(n98901), .ZN(n87856) );
  AOI22_X1 U88687 ( .A1(n105232), .A2(n69720), .B1(n98832), .B2(n111072), .ZN(
        n98901) );
  AND2_X2 U88688 ( .A1(stackBus_In[19]), .A2(n105205), .ZN(n94692) );
  OAI21_X1 U88689 ( .B1(n110197), .B2(n106274), .A(n98902), .ZN(
        \DLX_Datapath/RegisterFile/N22557 ) );
  AOI22_X1 U88690 ( .A1(n94694), .A2(n81258), .B1(n106107), .B2(n106273), .ZN(
        n98902) );
  NAND2_X1 U88691 ( .A1(n105500), .A2(n87974), .ZN(n81403) );
  OAI21_X1 U88692 ( .B1(n111064), .B2(n110120), .A(n98903), .ZN(n87974) );
  AOI22_X1 U88693 ( .A1(n105232), .A2(n69721), .B1(n98832), .B2(n111073), .ZN(
        n98903) );
  AND2_X2 U88694 ( .A1(stackBus_In[18]), .A2(n105199), .ZN(n94694) );
  OAI21_X1 U88695 ( .B1(n109982), .B2(n106274), .A(n98904), .ZN(
        \DLX_Datapath/RegisterFile/N22556 ) );
  AOI22_X1 U88696 ( .A1(n94696), .A2(n81258), .B1(n106222), .B2(n106273), .ZN(
        n98904) );
  NAND2_X1 U88697 ( .A1(n105500), .A2(n88092), .ZN(n81294) );
  OAI21_X1 U88698 ( .B1(n111064), .B2(n109903), .A(n98905), .ZN(n88092) );
  AOI22_X1 U88699 ( .A1(n105232), .A2(n69722), .B1(n98832), .B2(n111078), .ZN(
        n98905) );
  AND2_X2 U88700 ( .A1(stackBus_In[17]), .A2(n105205), .ZN(n94696) );
  OAI21_X1 U88701 ( .B1(n109865), .B2(n106274), .A(n98906), .ZN(
        \DLX_Datapath/RegisterFile/N22555 ) );
  AOI22_X1 U88702 ( .A1(n94698), .A2(n81258), .B1(n106112), .B2(n106273), .ZN(
        n98906) );
  NAND2_X1 U88703 ( .A1(n105501), .A2(n88210), .ZN(n81398) );
  OAI21_X1 U88704 ( .B1(n111064), .B2(n109785), .A(n98907), .ZN(n88210) );
  AOI22_X1 U88705 ( .A1(n105232), .A2(n69723), .B1(n98832), .B2(n111074), .ZN(
        n98907) );
  AND2_X2 U88706 ( .A1(stackBus_In[16]), .A2(n105205), .ZN(n94698) );
  OAI21_X1 U88707 ( .B1(n108239), .B2(n106274), .A(n98908), .ZN(
        \DLX_Datapath/RegisterFile/N22554 ) );
  AOI22_X1 U88708 ( .A1(n94700), .A2(n81258), .B1(n106234), .B2(n106273), .ZN(
        n98908) );
  NAND2_X1 U88709 ( .A1(n105502), .A2(n88328), .ZN(n81284) );
  OAI21_X1 U88710 ( .B1(n111064), .B2(n111116), .A(n98909), .ZN(n88328) );
  AOI22_X1 U88711 ( .A1(n105232), .A2(n69724), .B1(n98832), .B2(n111096), .ZN(
        n98909) );
  AND2_X2 U88712 ( .A1(stackBus_In[15]), .A2(n107022), .ZN(n94700) );
  OAI21_X1 U88713 ( .B1(n108362), .B2(n106274), .A(n98910), .ZN(
        \DLX_Datapath/RegisterFile/N22553 ) );
  AOI22_X1 U88714 ( .A1(n94702), .A2(n81258), .B1(n106174), .B2(n106273), .ZN(
        n98910) );
  NAND2_X1 U88715 ( .A1(n105500), .A2(n88446), .ZN(n81340) );
  OAI21_X1 U88716 ( .B1(n111064), .B2(n111117), .A(n98911), .ZN(n88446) );
  AOI22_X1 U88717 ( .A1(n98831), .A2(n69725), .B1(n98832), .B2(n111079), .ZN(
        n98911) );
  AND2_X2 U88718 ( .A1(stackBus_In[14]), .A2(n105199), .ZN(n94702) );
  OAI21_X1 U88719 ( .B1(n108473), .B2(n106274), .A(n98912), .ZN(
        \DLX_Datapath/RegisterFile/N22552 ) );
  AOI22_X1 U88720 ( .A1(n94704), .A2(n81258), .B1(n106239), .B2(n81260), .ZN(
        n98912) );
  NAND2_X1 U88721 ( .A1(n105502), .A2(n88564), .ZN(n81281) );
  OAI21_X1 U88722 ( .B1(n111064), .B2(n108282), .A(n98913), .ZN(n88564) );
  AOI22_X1 U88723 ( .A1(n105232), .A2(n69726), .B1(n98832), .B2(n111080), .ZN(
        n98913) );
  AND2_X2 U88724 ( .A1(stackBus_In[13]), .A2(n105205), .ZN(n94704) );
  OAI21_X1 U88725 ( .B1(n104523), .B2(n81256), .A(n98914), .ZN(
        \DLX_Datapath/RegisterFile/N22551 ) );
  AOI22_X1 U88726 ( .A1(n94706), .A2(n81258), .B1(n106073), .B2(n106273), .ZN(
        n98914) );
  NAND2_X1 U88727 ( .A1(n105502), .A2(n88682), .ZN(n81451) );
  OAI21_X1 U88728 ( .B1(n111064), .B2(n107631), .A(n98915), .ZN(n88682) );
  AOI22_X1 U88729 ( .A1(n105232), .A2(n69727), .B1(n98832), .B2(n111097), .ZN(
        n98915) );
  AND2_X2 U88730 ( .A1(stackBus_In[12]), .A2(n105200), .ZN(n94706) );
  OAI21_X1 U88731 ( .B1(n104522), .B2(n81256), .A(n98916), .ZN(
        \DLX_Datapath/RegisterFile/N22550 ) );
  AOI22_X1 U88732 ( .A1(n94708), .A2(n81258), .B1(n106201), .B2(n106273), .ZN(
        n98916) );
  NAND2_X1 U88733 ( .A1(n105500), .A2(n88800), .ZN(n81310) );
  OAI21_X1 U88734 ( .B1(n111064), .B2(n111110), .A(n98917), .ZN(n88800) );
  AOI22_X1 U88735 ( .A1(n105232), .A2(n69728), .B1(n98832), .B2(n111081), .ZN(
        n98917) );
  AND2_X2 U88736 ( .A1(stackBus_In[11]), .A2(n105200), .ZN(n94708) );
  OAI21_X1 U88737 ( .B1(n104521), .B2(n81256), .A(n98918), .ZN(
        \DLX_Datapath/RegisterFile/N22549 ) );
  AOI22_X1 U88738 ( .A1(n94710), .A2(n81258), .B1(n106247), .B2(n106273), .ZN(
        n98918) );
  NAND2_X1 U88739 ( .A1(n105501), .A2(n88918), .ZN(n81278) );
  OAI21_X1 U88740 ( .B1(n111064), .B2(n108510), .A(n98919), .ZN(n88918) );
  AOI22_X1 U88741 ( .A1(n105232), .A2(n69729), .B1(n98832), .B2(n111082), .ZN(
        n98919) );
  AND2_X2 U88742 ( .A1(stackBus_In[10]), .A2(n105203), .ZN(n94710) );
  OAI21_X1 U88743 ( .B1(n104520), .B2(n81256), .A(n98920), .ZN(
        \DLX_Datapath/RegisterFile/N22548 ) );
  AOI22_X1 U88744 ( .A1(n94712), .A2(n81258), .B1(n106161), .B2(n106273), .ZN(
        n98920) );
  NAND2_X1 U88745 ( .A1(n105501), .A2(n81794), .ZN(n81349) );
  OAI21_X1 U88746 ( .B1(n111064), .B2(n111111), .A(n98921), .ZN(n81794) );
  AOI22_X1 U88747 ( .A1(n105232), .A2(n69706), .B1(n98832), .B2(n111075), .ZN(
        n98921) );
  AND2_X2 U88748 ( .A1(stackBus_In[9]), .A2(n105203), .ZN(n94712) );
  OAI21_X1 U88749 ( .B1(n104519), .B2(n81256), .A(n98922), .ZN(
        \DLX_Datapath/RegisterFile/N22547 ) );
  AOI22_X1 U88750 ( .A1(n94714), .A2(n81258), .B1(n106117), .B2(n106273), .ZN(
        n98922) );
  NAND2_X1 U88751 ( .A1(n105501), .A2(n89153), .ZN(n81394) );
  OAI21_X1 U88752 ( .B1(n111064), .B2(n111112), .A(n98923), .ZN(n89153) );
  AOI22_X1 U88753 ( .A1(n105232), .A2(n69707), .B1(n98832), .B2(n111076), .ZN(
        n98923) );
  AND2_X2 U88754 ( .A1(stackBus_In[8]), .A2(n105201), .ZN(n94714) );
  OAI21_X1 U88755 ( .B1(n104518), .B2(n81256), .A(n98924), .ZN(
        \DLX_Datapath/RegisterFile/N22545 ) );
  AOI22_X1 U88756 ( .A1(n94717), .A2(n81258), .B1(n106263), .B2(n106273), .ZN(
        n98924) );
  NAND2_X1 U88757 ( .A1(n105502), .A2(n81792), .ZN(n81267) );
  OAI21_X1 U88758 ( .B1(n111064), .B2(n111113), .A(n98925), .ZN(n81792) );
  AOI22_X1 U88759 ( .A1(n105232), .A2(n69699), .B1(n98832), .B2(n111083), .ZN(
        n98925) );
  AND2_X2 U88760 ( .A1(stackBus_In[6]), .A2(n105201), .ZN(n94717) );
  OAI21_X1 U88761 ( .B1(n104517), .B2(n81256), .A(n98926), .ZN(
        \DLX_Datapath/RegisterFile/N22544 ) );
  AOI22_X1 U88762 ( .A1(n94719), .A2(n81258), .B1(n106047), .B2(n106273), .ZN(
        n98926) );
  NAND2_X1 U88763 ( .A1(n105502), .A2(n89506), .ZN(n81509) );
  OAI21_X1 U88764 ( .B1(n111064), .B2(n111114), .A(n98927), .ZN(n89506) );
  AOI22_X1 U88765 ( .A1(n105232), .A2(n69700), .B1(n98832), .B2(n111077), .ZN(
        n98927) );
  AND2_X2 U88766 ( .A1(stackBus_In[5]), .A2(n105199), .ZN(n94719) );
  OAI21_X1 U88767 ( .B1(n104516), .B2(n81256), .A(n98928), .ZN(
        \DLX_Datapath/RegisterFile/N22543 ) );
  AOI22_X1 U88768 ( .A1(n94721), .A2(n81258), .B1(n106052), .B2(n106273), .ZN(
        n98928) );
  NAND2_X1 U88769 ( .A1(n105500), .A2(n89624), .ZN(n81501) );
  OAI21_X1 U88770 ( .B1(n111064), .B2(n111115), .A(n98929), .ZN(n89624) );
  AOI22_X1 U88771 ( .A1(n105232), .A2(n69701), .B1(n98832), .B2(n111089), .ZN(
        n98929) );
  AND2_X2 U88772 ( .A1(stackBus_In[4]), .A2(n105203), .ZN(n94721) );
  OAI21_X1 U88773 ( .B1(n104515), .B2(n81256), .A(n98930), .ZN(
        \DLX_Datapath/RegisterFile/N22542 ) );
  AOI22_X1 U88774 ( .A1(n94723), .A2(n81258), .B1(n106097), .B2(n106273), .ZN(
        n98930) );
  NAND2_X1 U88775 ( .A1(n105501), .A2(n89742), .ZN(n81415) );
  OAI21_X1 U88776 ( .B1(n111064), .B2(n111107), .A(n98931), .ZN(n89742) );
  AOI22_X1 U88777 ( .A1(n105232), .A2(n69702), .B1(n98832), .B2(n111084), .ZN(
        n98931) );
  AND2_X2 U88778 ( .A1(stackBus_In[3]), .A2(n105202), .ZN(n94723) );
  OAI21_X1 U88779 ( .B1(n104514), .B2(n81256), .A(n98932), .ZN(
        \DLX_Datapath/RegisterFile/N22541 ) );
  AOI22_X1 U88780 ( .A1(n94725), .A2(n81258), .B1(n106057), .B2(n106273), .ZN(
        n98932) );
  NAND2_X1 U88781 ( .A1(n105502), .A2(n81790), .ZN(n81498) );
  OAI21_X1 U88782 ( .B1(n111064), .B2(n111108), .A(n98933), .ZN(n81790) );
  AOI22_X1 U88783 ( .A1(n105232), .A2(n69703), .B1(n98832), .B2(n111085), .ZN(
        n98933) );
  AND2_X2 U88784 ( .A1(stackBus_In[2]), .A2(n105202), .ZN(n94725) );
  OAI21_X1 U88785 ( .B1(n104513), .B2(n81256), .A(n98934), .ZN(
        \DLX_Datapath/RegisterFile/N22540 ) );
  AOI22_X1 U88786 ( .A1(n94727), .A2(n81258), .B1(n106273), .B2(n96125), .ZN(
        n98934) );
  NOR2_X1 U88787 ( .A1(n105089), .A2(n111058), .ZN(n96125) );
  OAI21_X1 U88788 ( .B1(n111064), .B2(n111109), .A(n98935), .ZN(n89977) );
  AOI22_X1 U88789 ( .A1(n105232), .A2(n69704), .B1(n98832), .B2(n111086), .ZN(
        n98935) );
  AND2_X2 U88790 ( .A1(stackBus_In[1]), .A2(n105200), .ZN(n94727) );
  OAI21_X1 U88791 ( .B1(n104512), .B2(n81256), .A(n98936), .ZN(
        \DLX_Datapath/RegisterFile/N22539 ) );
  AOI22_X1 U88792 ( .A1(n94729), .A2(n81258), .B1(n106270), .B2(n106273), .ZN(
        n98936) );
  NAND2_X1 U88793 ( .A1(n105502), .A2(n90096), .ZN(n81262) );
  OAI21_X1 U88794 ( .B1(n111064), .B2(n111106), .A(n98937), .ZN(n90096) );
  AOI22_X1 U88795 ( .A1(n69705), .A2(n105232), .B1(n98832), .B2(n111087), .ZN(
        n98937) );
  AND2_X2 U88796 ( .A1(n100629), .A2(n111064), .ZN(n98832) );
  NOR2_X1 U88797 ( .A1(n64655), .A2(n100629), .ZN(n98831) );
  AND2_X2 U88798 ( .A1(n98842), .A2(n98938), .ZN(n81258) );
  AND2_X2 U88799 ( .A1(stackBus_In[0]), .A2(n105200), .ZN(n94729) );
  NAND2_X1 U88800 ( .A1(n98840), .A2(n98938), .ZN(n81256) );
  NAND2_X1 U88801 ( .A1(n81260), .A2(n105501), .ZN(n98938) );
  NAND2_X1 U88802 ( .A1(n69424), .A2(n94093), .ZN(n95451) );
  AND2_X2 U88803 ( .A1(n94505), .A2(n98654), .ZN(n81260) );
  XOR2_X1 U88807 ( .A(n90133), .B(n107128), .Z(n95412) );
  XNOR2_X1 U88808 ( .A(n104491), .B(n96531), .ZN(n96530) );
  XNOR2_X1 U88809 ( .A(
        \add_0_root_sub_0_root_DLX_Datapath/RegisterFile/add_172/carry[6] ), 
        .B(\DLX_Datapath/RegisterFile/old_CWP2[2] ), .ZN(n96531) );
  NAND2_X1 U88810 ( .A1(\DLX_Datapath/RegisterFile/N9337 ), .A2(n98940), .ZN(
        n98941) );
  NOR2_X1 U88811 ( .A1(n90137), .A2(n90133), .ZN(n98940) );
  XNOR2_X1 U88812 ( .A(n81876), .B(n100801), .ZN(n90133) );
  AOI21_X1 U88813 ( .B1(n90137), .B2(n107131), .A(n104922), .ZN(n81876) );
  OAI21_X1 U88815 ( .B1(n98942), .B2(n107143), .A(n98943), .ZN(n94081) );
  NAND2_X1 U88816 ( .A1(n104730), .A2(n54623), .ZN(n98943) );
  NOR2_X1 U88817 ( .A1(n98615), .A2(n104762), .ZN(n94505) );
  OR2_X1 U88820 ( .A1(n98946), .A2(n90120), .ZN(n98615) );
  OAI21_X1 U88821 ( .B1(n105028), .B2(n107133), .A(n98947), .ZN(n90120) );
  NAND2_X1 U88822 ( .A1(n54614), .A2(n104730), .ZN(n98947) );
  NAND2_X1 U88823 ( .A1(n107123), .A2(n107122), .ZN(n98946) );
  OAI21_X1 U88824 ( .B1(n105028), .B2(n107135), .A(n98948), .ZN(n90119) );
  NAND2_X1 U88825 ( .A1(n54616), .A2(n104730), .ZN(n98948) );
  OAI21_X1 U88826 ( .B1(n105028), .B2(n107138), .A(n98949), .ZN(n90127) );
  NAND2_X1 U88827 ( .A1(n54618), .A2(n104730), .ZN(n98949) );
  OAI21_X1 U88830 ( .B1(n98842), .B2(n94366), .A(n105602), .ZN(n98840) );
  NAND2_X1 U88831 ( .A1(n86222), .A2(n80203), .ZN(n94663) );
  NOR2_X1 U88832 ( .A1(n95131), .A2(n96489), .ZN(n98842) );
  OR2_X1 U88833 ( .A1(n98614), .A2(n59515), .ZN(n96489) );
  NAND2_X1 U88834 ( .A1(n98613), .A2(n106764), .ZN(n98614) );
  NOR2_X1 U88835 ( .A1(n62212), .A2(
        \dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .ZN(n98613) );
  NAND2_X1 U88836 ( .A1(n104582), .A2(n111027), .ZN(n95131) );
  NOR2_X1 U88837 ( .A1(n107149), .A2(net73629), .ZN(\DLX_Datapath/N358 ) );
  NAND2_X1 U88838 ( .A1(n104753), .A2(n106847), .ZN(\DLX_Datapath/N357 ) );
  NOR2_X1 U88839 ( .A1(n104498), .A2(net113155), .ZN(\DLX_Datapath/N356 ) );
  NAND2_X1 U88840 ( .A1(net113102), .A2(n106936), .ZN(\DLX_Datapath/N355 ) );
  NOR2_X1 U88841 ( .A1(n104496), .A2(net113159), .ZN(\DLX_Datapath/N354 ) );
  NAND2_X1 U88842 ( .A1(n104753), .A2(n106942), .ZN(\DLX_Datapath/N353 ) );
  NOR2_X1 U88843 ( .A1(n59454), .A2(net113157), .ZN(\DLX_Datapath/N352 ) );
  NOR2_X1 U88844 ( .A1(n59453), .A2(net113155), .ZN(\DLX_Datapath/N351 ) );
  NOR2_X1 U88845 ( .A1(n59452), .A2(net113157), .ZN(\DLX_Datapath/N350 ) );
  NOR2_X1 U88846 ( .A1(n59451), .A2(net113156), .ZN(\DLX_Datapath/N349 ) );
  NOR2_X1 U88847 ( .A1(n59445), .A2(net113159), .ZN(\DLX_Datapath/N348 ) );
  NOR2_X1 U88848 ( .A1(n59444), .A2(net113156), .ZN(\DLX_Datapath/N347 ) );
  NOR2_X1 U88849 ( .A1(n59443), .A2(net113156), .ZN(\DLX_Datapath/N346 ) );
  NOR2_X1 U88850 ( .A1(n59442), .A2(net113155), .ZN(\DLX_Datapath/N345 ) );
  NOR2_X1 U88851 ( .A1(n59441), .A2(net113157), .ZN(\DLX_Datapath/N344 ) );
  NOR2_X1 U88852 ( .A1(n59435), .A2(net113156), .ZN(\DLX_Datapath/N343 ) );
  AOI21_X1 U88853 ( .B1(IR_in[17]), .B2(n111134), .A(n111135), .ZN(n82407) );
  NAND2_X1 U88854 ( .A1(IR_in[15]), .A2(n82399), .ZN(n82400) );
  OAI21_X1 U88855 ( .B1(n111148), .B2(n111147), .A(n82334), .ZN(n82399) );
  NOR2_X1 U88856 ( .A1(n80067), .A2(IR_in[30]), .ZN(n82334) );
  NAND2_X1 U88857 ( .A1(n98950), .A2(n111143), .ZN(n80067) );
  NOR2_X1 U88858 ( .A1(IR_in[31]), .A2(IR_in[29]), .ZN(n98950) );
  NAND2_X1 U88859 ( .A1(IR_in[27]), .A2(IR_in[26]), .ZN(n80064) );
  NAND2_X1 U88860 ( .A1(IR_in[27]), .A2(n111149), .ZN(n81975) );
  NAND2_X1 U88861 ( .A1(n98951), .A2(n98952), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [30]) );
  AOI22_X1 U88862 ( .A1(n98953), .A2(n69709), .B1(n98954), .B2(n111090), .ZN(
        n98952) );
  AOI22_X1 U88863 ( .A1(n105229), .A2(DataAddr[30]), .B1(n98956), .B2(n108043), 
        .ZN(n98951) );
  NAND2_X1 U88864 ( .A1(n98957), .A2(n98958), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [29]) );
  AOI22_X1 U88865 ( .A1(n98953), .A2(n69710), .B1(n98954), .B2(n111070), .ZN(
        n98958) );
  AOI22_X1 U88866 ( .A1(n105229), .A2(DataAddr[29]), .B1(n98956), .B2(n107420), 
        .ZN(n98957) );
  NAND4_X2 U88867 ( .A1(n98959), .A2(n98960), .A3(n98961), .A4(n98962), .ZN(
        \DLX_Datapath/ArithLogUnit/N193 ) );
  NOR4_X1 U88868 ( .A1(n98963), .A2(n98964), .A3(n98965), .A4(n98966), .ZN(
        n98962) );
  AOI21_X1 U88869 ( .B1(n98967), .B2(n98968), .A(n106956), .ZN(n98966) );
  AOI21_X1 U88870 ( .B1(n69802), .B2(n98969), .A(n98970), .ZN(n98968) );
  NOR3_X1 U88871 ( .A1(n98971), .A2(n69802), .A3(n98972), .ZN(n98970) );
  OAI21_X1 U88872 ( .B1(n98973), .B2(n110957), .A(n98974), .ZN(n98969) );
  OAI21_X1 U88873 ( .B1(n98975), .B2(n106950), .A(n110957), .ZN(n98974) );
  NOR2_X1 U88874 ( .A1(n98972), .A2(n98976), .ZN(n98975) );
  AOI22_X1 U88875 ( .A1(n98977), .A2(n106951), .B1(n98972), .B2(n106947), .ZN(
        n98967) );
  NOR2_X1 U88876 ( .A1(n98979), .A2(n107573), .ZN(n98965) );
  AOI22_X1 U88877 ( .A1(n79712), .A2(n107571), .B1(
        \DLX_Datapath/ArithLogUnit/A_log [0]), .B2(n79713), .ZN(n98979) );
  AND2_X2 U88878 ( .A1(\DLX_Datapath/ArithLogUnit/sel_log [3]), .A2(n106369), 
        .ZN(n79713) );
  AND2_X2 U88879 ( .A1(\DLX_Datapath/ArithLogUnit/sel_log [1]), .A2(n106369), 
        .ZN(n79712) );
  OAI33_X1 U88880 ( .A1(n107571), .A2(\DLX_Datapath/ArithLogUnit/B_log [0]), 
        .A3(n79714), .B1(n98980), .B2(n98981), .B3(n98977), .ZN(n98964) );
  NOR2_X1 U88881 ( .A1(n69801), .A2(n108747), .ZN(n98981) );
  NAND2_X1 U88882 ( .A1(\DLX_Datapath/ArithLogUnit/sel_log [2]), .A2(n106369), 
        .ZN(n79714) );
  AOI21_X1 U88883 ( .B1(n110957), .B2(n108747), .A(n106955), .ZN(n98963) );
  NOR4_X1 U88884 ( .A1(n98982), .A2(n98983), .A3(n98984), .A4(n98985), .ZN(
        n98972) );
  NAND2_X1 U88885 ( .A1(n98986), .A2(n98987), .ZN(n98985) );
  NOR4_X1 U88886 ( .A1(\DLX_Datapath/ArithLogUnit/Sum_cmp [16]), .A2(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [15]), .A3(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [14]), .A4(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [13]), .ZN(n98987) );
  NOR4_X1 U88887 ( .A1(\DLX_Datapath/ArithLogUnit/Sum_cmp [12]), .A2(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [11]), .A3(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [10]), .A4(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [0]), .ZN(n98986) );
  NAND2_X1 U88888 ( .A1(n98988), .A2(n98989), .ZN(n98984) );
  NOR4_X1 U88889 ( .A1(\DLX_Datapath/ArithLogUnit/Sum_cmp [23]), .A2(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [22]), .A3(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [21]), .A4(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [20]), .ZN(n98989) );
  NOR4_X1 U88890 ( .A1(\DLX_Datapath/ArithLogUnit/Sum_cmp [1]), .A2(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [19]), .A3(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [18]), .A4(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [17]), .ZN(n98988) );
  NAND2_X1 U88891 ( .A1(n98990), .A2(n98991), .ZN(n98983) );
  NOR4_X1 U88892 ( .A1(\DLX_Datapath/ArithLogUnit/Sum_cmp [30]), .A2(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [2]), .A3(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [29]), .A4(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [28]), .ZN(n98991) );
  NOR4_X1 U88893 ( .A1(\DLX_Datapath/ArithLogUnit/Sum_cmp [27]), .A2(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [26]), .A3(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [25]), .A4(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [24]), .ZN(n98990) );
  NAND2_X1 U88894 ( .A1(n98992), .A2(n98993), .ZN(n98982) );
  NOR4_X1 U88895 ( .A1(\DLX_Datapath/ArithLogUnit/Sum_cmp [9]), .A2(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [8]), .A3(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [7]), .A4(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [6]), .ZN(n98993) );
  NOR4_X1 U88896 ( .A1(\DLX_Datapath/ArithLogUnit/Sum_cmp [5]), .A2(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [4]), .A3(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [3]), .A4(
        \DLX_Datapath/ArithLogUnit/Sum_cmp [31]), .ZN(n98992) );
  XNOR2_X1 U88897 ( .A(\DLX_Datapath/ArithLogUnit/useBorrow_cmp ), .B(
        \DLX_Datapath/ArithLogUnit/Cout_cmp ), .ZN(n98977) );
  AOI22_X1 U88898 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N72 ), .A2(n79719), .B1(n104359), .B2(n79744), .ZN(n98961) );
  NAND2_X1 U88899 ( .A1(n98994), .A2(n98995), .ZN(n79744) );
  NOR2_X1 U88900 ( .A1(n105226), .A2(n105096), .ZN(n98994) );
  XOR2_X1 U88901 ( .A(\DLX_Datapath/ArithLogUnit/A_add [0]), .B(n98997), .Z(
        n104359) );
  XOR2_X1 U88902 ( .A(\DLX_Datapath/ArithLogUnit/Cin_add ), .B(
        \DLX_Datapath/ArithLogUnit/B_add [0]), .Z(n98997) );
  AND2_X2 U88903 ( .A1(\DLX_Datapath/ArithLogUnit/sel_shf [1]), .A2(n82617), 
        .ZN(n79719) );
  NAND2_X1 U88904 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N40 ), .A2(n79718), .ZN(n98960) );
  AND2_X2 U88905 ( .A1(n98998), .A2(\DLX_Datapath/ArithLogUnit/sel_shf [0]), 
        .ZN(n79718) );
  NOR2_X1 U88906 ( .A1(\DLX_Datapath/ArithLogUnit/sel_shf [1]), .A2(n106949), 
        .ZN(n98998) );
  AOI22_X1 U88907 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_shift/N8 ), .A2(n106356), .B1(n105123), .B2(\DLX_Datapath/MUX_HDU_ALUInB [0]), .ZN(n98959) );
  NOR4_X1 U88908 ( .A1(n69801), .A2(n69800), .A3(n69330), .A4(n98999), .ZN(
        n79746) );
  NOR2_X1 U88909 ( .A1(n99000), .A2(n106949), .ZN(n79716) );
  OAI21_X1 U88910 ( .B1(n99001), .B2(n98973), .A(n99002), .ZN(n82617) );
  NOR2_X1 U88911 ( .A1(n60443), .A2(n60442), .ZN(n99002) );
  NOR2_X1 U88912 ( .A1(n99001), .A2(n98971), .ZN(n60442) );
  NOR2_X1 U88913 ( .A1(n99001), .A2(n98978), .ZN(n60443) );
  OR2_X1 U88914 ( .A1(\DLX_Datapath/ArithLogUnit/sel_shf [1]), .A2(
        \DLX_Datapath/ArithLogUnit/sel_shf [0]), .ZN(n99000) );
  NOR2_X1 U88915 ( .A1(n99003), .A2(n99004), .ZN(
        \DLX_Datapath/ArithLogUnit/N187 ) );
  XOR2_X1 U88916 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [31]), .B(n106926), .Z(
        n99004) );
  NAND2_X1 U88917 ( .A1(n99005), .A2(n99006), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [31]) );
  AOI22_X1 U88918 ( .A1(n98953), .A2(n69708), .B1(n98954), .B2(n111069), .ZN(
        n99006) );
  AOI22_X1 U88919 ( .A1(n105229), .A2(DataAddr[31]), .B1(n98956), .B2(n107947), 
        .ZN(n99005) );
  AOI21_X1 U88920 ( .B1(n98978), .B2(n98971), .A(n98999), .ZN(
        \DLX_Datapath/ArithLogUnit/N180 ) );
  OAI21_X1 U88921 ( .B1(n98999), .B2(n98971), .A(n106952), .ZN(
        \DLX_Datapath/ArithLogUnit/N178 ) );
  OAI21_X1 U88922 ( .B1(n98978), .B2(n98999), .A(n99007), .ZN(
        \DLX_Datapath/ArithLogUnit/N179 ) );
  NAND2_X1 U88923 ( .A1(n99008), .A2(n69339), .ZN(n99007) );
  NOR2_X1 U88924 ( .A1(n69802), .A2(n98976), .ZN(n99008) );
  OAI21_X1 U88925 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [31]), .B2(n106946), .A(
        n99009), .ZN(\DLX_Datapath/ArithLogUnit/N176 ) );
  AOI22_X1 U88926 ( .A1(n99010), .A2(n105097), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [31]), .ZN(n99009) );
  OAI21_X1 U88927 ( .B1(n107480), .B2(n107491), .A(n99011), .ZN(n99010) );
  OAI21_X1 U88928 ( .B1(n99012), .B2(n81812), .A(n107481), .ZN(n99011) );
  OAI21_X1 U88929 ( .B1(n81817), .B2(n107558), .A(n99013), .ZN(n81812) );
  AOI21_X1 U88930 ( .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[16] ), .B2(
        n81819), .A(n108267), .ZN(n99013) );
  OAI21_X1 U88931 ( .B1(n99015), .B2(n99016), .A(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99014) );
  OAI21_X1 U88932 ( .B1(n99017), .B2(n99018), .A(n99019), .ZN(n99012) );
  NAND2_X1 U88933 ( .A1(n99020), .A2(n99021), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [31]) );
  AOI21_X1 U88934 ( .B1(n69708), .B2(n99022), .A(n99023), .ZN(n99021) );
  OAI21_X1 U88935 ( .B1(n99024), .B2(n104671), .A(n99025), .ZN(n99023) );
  NAND2_X1 U88936 ( .A1(n69795), .A2(n106927), .ZN(n99025) );
  AOI22_X1 U88937 ( .A1(n105224), .A2(n111069), .B1(n99027), .B2(DataAddr[31]), 
        .ZN(n99020) );
  OAI21_X1 U88938 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [30]), .B2(n106946), .A(
        n99028), .ZN(\DLX_Datapath/ArithLogUnit/N175 ) );
  AOI22_X1 U88939 ( .A1(n99029), .A2(n105096), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [30]), .ZN(n99028) );
  OAI21_X1 U88940 ( .B1(n107479), .B2(n81806), .A(n99030), .ZN(n99029) );
  OAI21_X1 U88941 ( .B1(n107481), .B2(n99031), .A(n81808), .ZN(n99030) );
  NAND2_X1 U88942 ( .A1(n99032), .A2(n99033), .ZN(n81808) );
  AOI22_X1 U88943 ( .A1(n105121), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] ), .B2(n105122), .ZN(
        n99033) );
  AOI22_X1 U88944 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] ), .A2(
        n108272), .B1(n99016), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99032) );
  XNOR2_X1 U88945 ( .A(n99034), .B(n99035), .ZN(n81806) );
  XNOR2_X1 U88946 ( .A(n99017), .B(n99036), .ZN(n99035) );
  AOI21_X1 U88947 ( .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[17] ), .B2(
        n99037), .A(n107557), .ZN(n99017) );
  AOI21_X1 U88948 ( .B1(n105119), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[17] ), .A(n99040), .ZN(n99038)
         );
  OAI21_X1 U88949 ( .B1(n99041), .B2(n99018), .A(n99019), .ZN(n99031) );
  NAND2_X1 U88950 ( .A1(n99034), .A2(n99036), .ZN(n99019) );
  NOR2_X1 U88951 ( .A1(n99036), .A2(n99034), .ZN(n99018) );
  NAND2_X1 U88952 ( .A1(n99042), .A2(n99043), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [30]) );
  AOI21_X1 U88953 ( .B1(n69709), .B2(n99022), .A(n99044), .ZN(n99043) );
  OAI21_X1 U88954 ( .B1(n99024), .B2(n104670), .A(n99045), .ZN(n99044) );
  NAND2_X1 U88955 ( .A1(n69796), .A2(n106927), .ZN(n99045) );
  AOI22_X1 U88956 ( .A1(n105224), .A2(n111090), .B1(n99027), .B2(DataAddr[30]), 
        .ZN(n99042) );
  OAI21_X1 U88957 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [29]), .B2(n106946), .A(
        n99046), .ZN(\DLX_Datapath/ArithLogUnit/N174 ) );
  AOI22_X1 U88958 ( .A1(n99047), .A2(n105096), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [29]), .ZN(n99046) );
  OAI21_X1 U88959 ( .B1(n99048), .B2(n99049), .A(n107477), .ZN(n99047) );
  AOI21_X1 U88960 ( .B1(n99049), .B2(n99048), .A(n99051), .ZN(n99050) );
  NAND2_X1 U88961 ( .A1(n99052), .A2(n99053), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [29]) );
  AOI21_X1 U88962 ( .B1(n69710), .B2(n99022), .A(n99054), .ZN(n99053) );
  OAI21_X1 U88963 ( .B1(n99024), .B2(n104669), .A(n99055), .ZN(n99054) );
  NAND2_X1 U88964 ( .A1(n69797), .A2(n106927), .ZN(n99055) );
  AOI22_X1 U88965 ( .A1(n105224), .A2(n111070), .B1(n99027), .B2(DataAddr[29]), 
        .ZN(n99052) );
  OAI21_X1 U88966 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [28]), .B2(n106946), .A(
        n99056), .ZN(\DLX_Datapath/ArithLogUnit/N173 ) );
  AOI22_X1 U88967 ( .A1(n99057), .A2(n105096), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [28]), .ZN(n99056) );
  OAI21_X1 U88968 ( .B1(n107505), .B2(n99058), .A(n99059), .ZN(n99057) );
  OAI21_X1 U88969 ( .B1(n107476), .B2(n99060), .A(n99061), .ZN(n99059) );
  NAND2_X1 U88970 ( .A1(n99062), .A2(n99063), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [28]) );
  AOI21_X1 U88971 ( .B1(n69711), .B2(n99022), .A(n99064), .ZN(n99063) );
  OAI21_X1 U88972 ( .B1(n99024), .B2(n104668), .A(n99065), .ZN(n99064) );
  NAND2_X1 U88973 ( .A1(n69798), .A2(n106927), .ZN(n99065) );
  AOI22_X1 U88974 ( .A1(n105224), .A2(n111091), .B1(n99027), .B2(DataAddr[28]), 
        .ZN(n99062) );
  OAI21_X1 U88975 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [27]), .B2(n106946), .A(
        n99066), .ZN(\DLX_Datapath/ArithLogUnit/N172 ) );
  AOI22_X1 U88976 ( .A1(n99067), .A2(n105097), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [27]), .ZN(n99066) );
  OAI21_X1 U88977 ( .B1(n99068), .B2(n99069), .A(n107470), .ZN(n99067) );
  AOI21_X1 U88978 ( .B1(n99069), .B2(n99068), .A(n99071), .ZN(n99070) );
  NAND2_X1 U88979 ( .A1(n99072), .A2(n99073), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [27]) );
  AOI21_X1 U88980 ( .B1(n69712), .B2(n99022), .A(n99074), .ZN(n99073) );
  OAI21_X1 U88981 ( .B1(n99024), .B2(n104667), .A(n99075), .ZN(n99074) );
  NAND2_X1 U88982 ( .A1(n69799), .A2(n106927), .ZN(n99075) );
  AOI22_X1 U88983 ( .A1(n105224), .A2(n111092), .B1(n99027), .B2(DataAddr[27]), 
        .ZN(n99072) );
  OAI21_X1 U88984 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [26]), .B2(n106946), .A(
        n99076), .ZN(\DLX_Datapath/ArithLogUnit/N171 ) );
  AOI22_X1 U88985 ( .A1(n99077), .A2(n105096), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [26]), .ZN(n99076) );
  OAI21_X1 U88986 ( .B1(n107514), .B2(n99078), .A(n99079), .ZN(n99077) );
  OAI21_X1 U88987 ( .B1(n107465), .B2(n99080), .A(n99081), .ZN(n99079) );
  NAND2_X1 U88988 ( .A1(n99082), .A2(n99083), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [26]) );
  AOI21_X1 U88989 ( .B1(n69713), .B2(n99022), .A(n99084), .ZN(n99083) );
  OAI21_X1 U88990 ( .B1(n99024), .B2(n104666), .A(n99085), .ZN(n99084) );
  NAND2_X1 U88991 ( .A1(n69784), .A2(n106927), .ZN(n99085) );
  AOI22_X1 U88992 ( .A1(n105224), .A2(n111093), .B1(n99027), .B2(DataAddr[26]), 
        .ZN(n99082) );
  OAI21_X1 U88993 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [25]), .B2(n106946), .A(
        n99086), .ZN(\DLX_Datapath/ArithLogUnit/N170 ) );
  AOI22_X1 U88994 ( .A1(n99087), .A2(n105097), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [25]), .ZN(n99086) );
  OAI21_X1 U88995 ( .B1(n99088), .B2(n99089), .A(n107459), .ZN(n99087) );
  AOI21_X1 U88996 ( .B1(n99089), .B2(n99088), .A(n99091), .ZN(n99090) );
  NAND2_X1 U88997 ( .A1(n99092), .A2(n99093), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [25]) );
  AOI21_X1 U88998 ( .B1(n69714), .B2(n99022), .A(n99094), .ZN(n99093) );
  OAI21_X1 U88999 ( .B1(n99024), .B2(n104665), .A(n99095), .ZN(n99094) );
  NAND2_X1 U89000 ( .A1(n69785), .A2(n106927), .ZN(n99095) );
  AOI22_X1 U89001 ( .A1(n105224), .A2(n111094), .B1(n99027), .B2(DataAddr[25]), 
        .ZN(n99092) );
  OAI21_X1 U89002 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [24]), .B2(n106946), .A(
        n99096), .ZN(\DLX_Datapath/ArithLogUnit/N169 ) );
  AOI22_X1 U89003 ( .A1(n99097), .A2(n105097), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [24]), .ZN(n99096) );
  OAI21_X1 U89004 ( .B1(n99098), .B2(n107454), .A(n99099), .ZN(n99097) );
  OAI21_X1 U89005 ( .B1(n99100), .B2(n107458), .A(n99101), .ZN(n99099) );
  NAND2_X1 U89006 ( .A1(n99102), .A2(n99103), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [24]) );
  AOI21_X1 U89007 ( .B1(n69715), .B2(n99022), .A(n99104), .ZN(n99103) );
  OAI21_X1 U89008 ( .B1(n99024), .B2(n104664), .A(n99105), .ZN(n99104) );
  NAND2_X1 U89009 ( .A1(n69786), .A2(n106927), .ZN(n99105) );
  AOI22_X1 U89010 ( .A1(n105224), .A2(n111095), .B1(n99027), .B2(DataAddr[24]), 
        .ZN(n99102) );
  OAI21_X1 U89011 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [23]), .B2(n106946), .A(
        n99106), .ZN(\DLX_Datapath/ArithLogUnit/N168 ) );
  AOI22_X1 U89012 ( .A1(n99107), .A2(n105096), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [23]), .ZN(n99106) );
  OAI21_X1 U89013 ( .B1(n107532), .B2(n107453), .A(n99108), .ZN(n99107) );
  OAI21_X1 U89014 ( .B1(n99109), .B2(n99110), .A(n99111), .ZN(n99108) );
  NAND2_X1 U89015 ( .A1(n99112), .A2(n99113), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [23]) );
  AOI21_X1 U89016 ( .B1(n69716), .B2(n105225), .A(n99114), .ZN(n99113) );
  OAI21_X1 U89017 ( .B1(n99024), .B2(n104663), .A(n99115), .ZN(n99114) );
  NAND2_X1 U89018 ( .A1(n69787), .A2(n106927), .ZN(n99115) );
  AOI22_X1 U89019 ( .A1(n99026), .A2(n111071), .B1(n105223), .B2(DataAddr[23]), 
        .ZN(n99112) );
  OAI21_X1 U89020 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [22]), .B2(n106946), .A(
        n99116), .ZN(\DLX_Datapath/ArithLogUnit/N167 ) );
  AOI22_X1 U89021 ( .A1(n99117), .A2(n105098), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [22]), .ZN(n99116) );
  OAI21_X1 U89022 ( .B1(n107535), .B2(n107446), .A(n99118), .ZN(n99117) );
  OAI21_X1 U89023 ( .B1(n99119), .B2(n99120), .A(n99121), .ZN(n99118) );
  NAND2_X1 U89024 ( .A1(n99122), .A2(n99123), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [22]) );
  AOI21_X1 U89025 ( .B1(n69717), .B2(n105225), .A(n99124), .ZN(n99123) );
  OAI21_X1 U89026 ( .B1(n99024), .B2(n104662), .A(n99125), .ZN(n99124) );
  NAND2_X1 U89027 ( .A1(n69788), .A2(n106927), .ZN(n99125) );
  AOI22_X1 U89028 ( .A1(n99026), .A2(n111066), .B1(n105223), .B2(DataAddr[22]), 
        .ZN(n99122) );
  OAI21_X1 U89029 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [21]), .B2(n106946), .A(
        n99126), .ZN(\DLX_Datapath/ArithLogUnit/N166 ) );
  AOI22_X1 U89030 ( .A1(n99127), .A2(n105098), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [21]), .ZN(n99126) );
  OAI21_X1 U89031 ( .B1(n99128), .B2(n107441), .A(n99129), .ZN(n99127) );
  OAI21_X1 U89032 ( .B1(n99130), .B2(n107437), .A(n99131), .ZN(n99129) );
  NAND2_X1 U89033 ( .A1(n99132), .A2(n99133), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [21]) );
  AOI21_X1 U89034 ( .B1(n69718), .B2(n105225), .A(n99134), .ZN(n99133) );
  OAI21_X1 U89035 ( .B1(n99024), .B2(n104661), .A(n99135), .ZN(n99134) );
  NAND2_X1 U89036 ( .A1(n69789), .A2(n106927), .ZN(n99135) );
  AOI22_X1 U89037 ( .A1(n105224), .A2(n111067), .B1(n105223), .B2(DataAddr[21]), .ZN(n99132) );
  OAI21_X1 U89038 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [20]), .B2(n106946), .A(
        n99136), .ZN(\DLX_Datapath/ArithLogUnit/N165 ) );
  AOI22_X1 U89039 ( .A1(n99137), .A2(n105097), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [20]), .ZN(n99136) );
  OAI21_X1 U89040 ( .B1(n107436), .B2(n99138), .A(n99139), .ZN(n99137) );
  OAI21_X1 U89041 ( .B1(n107434), .B2(n99140), .A(n99141), .ZN(n99139) );
  NAND2_X1 U89042 ( .A1(n99142), .A2(n99143), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [20]) );
  AOI21_X1 U89043 ( .B1(n69719), .B2(n105225), .A(n99144), .ZN(n99143) );
  OAI21_X1 U89044 ( .B1(n99024), .B2(n104660), .A(n99145), .ZN(n99144) );
  NAND2_X1 U89045 ( .A1(n69790), .A2(n106927), .ZN(n99145) );
  AOI22_X1 U89046 ( .A1(n105224), .A2(n111068), .B1(n105223), .B2(DataAddr[20]), .ZN(n99142) );
  OAI21_X1 U89047 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [19]), .B2(n105197), .A(
        n99146), .ZN(\DLX_Datapath/ArithLogUnit/N164 ) );
  AOI22_X1 U89048 ( .A1(n99147), .A2(n105096), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [19]), .ZN(n99146) );
  OAI21_X1 U89049 ( .B1(n99148), .B2(n99149), .A(n107432), .ZN(n99147) );
  AOI21_X1 U89050 ( .B1(n99149), .B2(n99148), .A(n99151), .ZN(n99150) );
  NAND2_X1 U89051 ( .A1(n99152), .A2(n99153), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [19]) );
  AOI21_X1 U89052 ( .B1(n69720), .B2(n105225), .A(n99154), .ZN(n99153) );
  OAI21_X1 U89053 ( .B1(n99024), .B2(n104659), .A(n99155), .ZN(n99154) );
  NAND2_X1 U89054 ( .A1(n69791), .A2(n106927), .ZN(n99155) );
  AOI22_X1 U89055 ( .A1(n105224), .A2(n111072), .B1(n105223), .B2(DataAddr[19]), .ZN(n99152) );
  OAI21_X1 U89056 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [18]), .B2(n106946), .A(
        n99156), .ZN(\DLX_Datapath/ArithLogUnit/N163 ) );
  AOI22_X1 U89057 ( .A1(n99157), .A2(n105097), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [18]), .ZN(n99156) );
  OAI21_X1 U89058 ( .B1(n99158), .B2(n99159), .A(n107431), .ZN(n99157) );
  AOI21_X1 U89059 ( .B1(n99159), .B2(n99158), .A(n99161), .ZN(n99160) );
  NAND2_X1 U89060 ( .A1(n99162), .A2(n99163), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [18]) );
  AOI21_X1 U89061 ( .B1(n69721), .B2(n105225), .A(n99164), .ZN(n99163) );
  OAI21_X1 U89062 ( .B1(n99024), .B2(n104658), .A(n99165), .ZN(n99164) );
  NAND2_X1 U89063 ( .A1(n69792), .A2(n106927), .ZN(n99165) );
  AOI22_X1 U89064 ( .A1(n105224), .A2(n111073), .B1(n105223), .B2(DataAddr[18]), .ZN(n99162) );
  OAI21_X1 U89065 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [17]), .B2(n105197), .A(
        n99166), .ZN(\DLX_Datapath/ArithLogUnit/N162 ) );
  AOI22_X1 U89066 ( .A1(n99167), .A2(n105098), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [17]), .ZN(n99166) );
  OAI21_X1 U89067 ( .B1(n107552), .B2(n107485), .A(n99168), .ZN(n99167) );
  OAI21_X1 U89068 ( .B1(n99169), .B2(n99170), .A(n99171), .ZN(n99168) );
  NAND2_X1 U89069 ( .A1(n99172), .A2(n99173), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [17]) );
  AOI21_X1 U89070 ( .B1(n69722), .B2(n105225), .A(n99174), .ZN(n99173) );
  OAI21_X1 U89071 ( .B1(n99024), .B2(n104657), .A(n99175), .ZN(n99174) );
  NAND2_X1 U89072 ( .A1(n69793), .A2(n106927), .ZN(n99175) );
  AOI22_X1 U89073 ( .A1(n105224), .A2(n111078), .B1(n105223), .B2(DataAddr[17]), .ZN(n99172) );
  OAI21_X1 U89074 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [16]), .B2(n106946), .A(
        n99176), .ZN(\DLX_Datapath/ArithLogUnit/N161 ) );
  AOI22_X1 U89075 ( .A1(n99177), .A2(n105097), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [16]), .ZN(n99176) );
  OAI21_X1 U89076 ( .B1(n107425), .B2(n99178), .A(n99179), .ZN(n99177) );
  OAI21_X1 U89077 ( .B1(n107492), .B2(n99180), .A(n99181), .ZN(n99179) );
  NAND2_X1 U89078 ( .A1(n99182), .A2(n99183), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [16]) );
  AOI21_X1 U89079 ( .B1(n69723), .B2(n105225), .A(n99184), .ZN(n99183) );
  OAI21_X1 U89080 ( .B1(n99024), .B2(n104656), .A(n99185), .ZN(n99184) );
  NAND2_X1 U89081 ( .A1(n69794), .A2(n106927), .ZN(n99185) );
  AOI22_X1 U89082 ( .A1(n105224), .A2(n111074), .B1(n105223), .B2(DataAddr[16]), .ZN(n99182) );
  OAI21_X1 U89083 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [15]), .B2(n105197), .A(
        n99187), .ZN(\DLX_Datapath/ArithLogUnit/N160 ) );
  AOI22_X1 U89084 ( .A1(n99188), .A2(n99189), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [15]), .ZN(n99187) );
  AND2_X2 U89085 ( .A1(n105098), .A2(n99190), .ZN(n99188) );
  NAND2_X1 U89086 ( .A1(n99191), .A2(n99192), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [15]) );
  AOI21_X1 U89087 ( .B1(n69724), .B2(n105225), .A(n99193), .ZN(n99192) );
  OAI21_X1 U89088 ( .B1(n100633), .B2(n99186), .A(n99194), .ZN(n99193) );
  NAND2_X1 U89089 ( .A1(n70872), .A2(n106929), .ZN(n99194) );
  AOI22_X1 U89090 ( .A1(n105224), .A2(n111096), .B1(n105223), .B2(DataAddr[15]), .ZN(n99191) );
  OAI21_X1 U89091 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [14]), .B2(n106946), .A(
        n99195), .ZN(\DLX_Datapath/ArithLogUnit/N159 ) );
  AOI22_X1 U89092 ( .A1(n99196), .A2(n105096), .B1(n105226), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [14]), .ZN(n99195) );
  OAI21_X1 U89093 ( .B1(n107426), .B2(n107511), .A(n99197), .ZN(n99196) );
  OAI21_X1 U89094 ( .B1(n99198), .B2(n99199), .A(n99200), .ZN(n99197) );
  NAND2_X1 U89095 ( .A1(n99201), .A2(n99202), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [14]) );
  AOI21_X1 U89096 ( .B1(n69725), .B2(n105225), .A(n99203), .ZN(n99202) );
  OAI21_X1 U89097 ( .B1(n100634), .B2(n99186), .A(n99204), .ZN(n99203) );
  NAND2_X1 U89098 ( .A1(n71026), .A2(n106929), .ZN(n99204) );
  AOI22_X1 U89099 ( .A1(n105224), .A2(n111079), .B1(n105223), .B2(DataAddr[14]), .ZN(n99201) );
  OAI21_X1 U89100 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [13]), .B2(n105197), .A(
        n99205), .ZN(\DLX_Datapath/ArithLogUnit/N158 ) );
  AOI22_X1 U89101 ( .A1(n99206), .A2(n99207), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [13]), .ZN(n99205) );
  NOR2_X1 U89102 ( .A1(n105900), .A2(n99208), .ZN(n99206) );
  NAND2_X1 U89103 ( .A1(n99209), .A2(n99210), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [13]) );
  AOI21_X1 U89104 ( .B1(n69726), .B2(n105225), .A(n99211), .ZN(n99210) );
  OAI21_X1 U89105 ( .B1(n100635), .B2(n99186), .A(n99212), .ZN(n99211) );
  NAND2_X1 U89106 ( .A1(n71169), .A2(n106929), .ZN(n99212) );
  AOI22_X1 U89107 ( .A1(n105224), .A2(n111080), .B1(n105223), .B2(DataAddr[13]), .ZN(n99209) );
  OAI21_X1 U89108 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [12]), .B2(n105197), .A(
        n99213), .ZN(\DLX_Datapath/ArithLogUnit/N157 ) );
  AOI22_X1 U89109 ( .A1(n99214), .A2(n105096), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [12]), .ZN(n99213) );
  OAI21_X1 U89110 ( .B1(n107427), .B2(n99215), .A(n99216), .ZN(n99214) );
  OAI21_X1 U89111 ( .B1(n107519), .B2(n99217), .A(n99218), .ZN(n99216) );
  NAND2_X1 U89112 ( .A1(n99219), .A2(n99220), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [12]) );
  AOI21_X1 U89113 ( .B1(n69727), .B2(n105225), .A(n99221), .ZN(n99220) );
  OAI21_X1 U89114 ( .B1(n100636), .B2(n99186), .A(n99222), .ZN(n99221) );
  NAND2_X1 U89115 ( .A1(n70130), .A2(n106929), .ZN(n99222) );
  AOI22_X1 U89116 ( .A1(n105224), .A2(n111097), .B1(n105223), .B2(DataAddr[12]), .ZN(n99219) );
  OAI21_X1 U89117 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [11]), .B2(n105197), .A(
        n99223), .ZN(\DLX_Datapath/ArithLogUnit/N156 ) );
  AOI22_X1 U89118 ( .A1(n99224), .A2(n99225), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [11]), .ZN(n99223) );
  NOR2_X1 U89119 ( .A1(n105899), .A2(n99226), .ZN(n99224) );
  NAND2_X1 U89120 ( .A1(n99227), .A2(n99228), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [11]) );
  AOI21_X1 U89121 ( .B1(n69728), .B2(n99022), .A(n99229), .ZN(n99228) );
  OAI21_X1 U89122 ( .B1(n100637), .B2(n99186), .A(n99230), .ZN(n99229) );
  NAND2_X1 U89123 ( .A1(n72661), .A2(n106929), .ZN(n99230) );
  AOI22_X1 U89124 ( .A1(n99026), .A2(n111081), .B1(n99027), .B2(DataAddr[11]), 
        .ZN(n99227) );
  OAI21_X1 U89125 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [10]), .B2(n105197), .A(
        n99231), .ZN(\DLX_Datapath/ArithLogUnit/N155 ) );
  AOI22_X1 U89126 ( .A1(n99232), .A2(n81804), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [10]), .ZN(n99231) );
  OAI21_X1 U89127 ( .B1(n99233), .B2(n99234), .A(n107428), .ZN(n99232) );
  AOI21_X1 U89128 ( .B1(n99234), .B2(n99233), .A(n99236), .ZN(n99235) );
  NAND2_X1 U89129 ( .A1(n99237), .A2(n99238), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [10]) );
  AOI21_X1 U89130 ( .B1(n69729), .B2(n99022), .A(n99239), .ZN(n99238) );
  OAI21_X1 U89131 ( .B1(n100638), .B2(n99186), .A(n99240), .ZN(n99239) );
  NAND2_X1 U89132 ( .A1(n72808), .A2(n106929), .ZN(n99240) );
  AOI22_X1 U89133 ( .A1(n99026), .A2(n111082), .B1(n99027), .B2(DataAddr[10]), 
        .ZN(n99237) );
  OAI21_X1 U89134 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [9]), .B2(n105197), .A(
        n99241), .ZN(\DLX_Datapath/ArithLogUnit/N154 ) );
  AOI22_X1 U89135 ( .A1(n99242), .A2(n99243), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [9]), .ZN(n99241) );
  NOR2_X1 U89136 ( .A1(n105900), .A2(n99244), .ZN(n99242) );
  NAND2_X1 U89137 ( .A1(n99245), .A2(n99246), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [9]) );
  AOI21_X1 U89138 ( .B1(n69706), .B2(n99022), .A(n99247), .ZN(n99246) );
  OAI21_X1 U89139 ( .B1(n100639), .B2(n99186), .A(n99248), .ZN(n99247) );
  NAND2_X1 U89140 ( .A1(n72803), .A2(n106929), .ZN(n99248) );
  AOI22_X1 U89141 ( .A1(n99026), .A2(n111075), .B1(n99027), .B2(DataAddr[9]), 
        .ZN(n99245) );
  OAI21_X1 U89142 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [8]), .B2(n105197), .A(
        n99249), .ZN(\DLX_Datapath/ArithLogUnit/N153 ) );
  AOI22_X1 U89143 ( .A1(n99250), .A2(n105098), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [8]), .ZN(n99249) );
  OAI21_X1 U89144 ( .B1(n99251), .B2(n99252), .A(n107429), .ZN(n99250) );
  AOI21_X1 U89145 ( .B1(n99252), .B2(n99251), .A(n99254), .ZN(n99253) );
  NAND2_X1 U89146 ( .A1(n99255), .A2(n99256), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [8]) );
  AOI21_X1 U89147 ( .B1(n69707), .B2(n105225), .A(n99257), .ZN(n99256) );
  OAI21_X1 U89148 ( .B1(n100640), .B2(n99186), .A(n99258), .ZN(n99257) );
  NAND2_X1 U89149 ( .A1(n72511), .A2(n106929), .ZN(n99258) );
  AOI22_X1 U89150 ( .A1(n99026), .A2(n111076), .B1(n99027), .B2(DataAddr[8]), 
        .ZN(n99255) );
  OAI21_X1 U89151 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [7]), .B2(n105197), .A(
        n99259), .ZN(\DLX_Datapath/ArithLogUnit/N152 ) );
  AOI22_X1 U89152 ( .A1(n99260), .A2(n99261), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [7]), .ZN(n99259) );
  NOR2_X1 U89153 ( .A1(n105900), .A2(n99262), .ZN(n99260) );
  NAND2_X1 U89154 ( .A1(n99263), .A2(n99264), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [7]) );
  AOI21_X1 U89155 ( .B1(n69730), .B2(n105225), .A(n99265), .ZN(n99264) );
  OAI21_X1 U89156 ( .B1(n100641), .B2(n99186), .A(n99266), .ZN(n99265) );
  NAND2_X1 U89157 ( .A1(n71913), .A2(n106929), .ZN(n99266) );
  AOI22_X1 U89158 ( .A1(n99026), .A2(n111088), .B1(n105223), .B2(DataAddr[7]), 
        .ZN(n99263) );
  OAI21_X1 U89159 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [6]), .B2(n105197), .A(
        n99267), .ZN(\DLX_Datapath/ArithLogUnit/N151 ) );
  AOI22_X1 U89160 ( .A1(n99268), .A2(n105097), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [6]), .ZN(n99267) );
  OAI21_X1 U89161 ( .B1(n107551), .B2(n107430), .A(n99269), .ZN(n99268) );
  OAI21_X1 U89162 ( .B1(n99270), .B2(n99271), .A(n99272), .ZN(n99269) );
  NAND2_X1 U89163 ( .A1(n99273), .A2(n99274), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [6]) );
  AOI21_X1 U89164 ( .B1(n69699), .B2(n105225), .A(n99275), .ZN(n99274) );
  OAI21_X1 U89165 ( .B1(n100642), .B2(n99186), .A(n99276), .ZN(n99275) );
  NAND2_X1 U89166 ( .A1(n72362), .A2(n106929), .ZN(n99276) );
  AOI22_X1 U89167 ( .A1(n99026), .A2(n111083), .B1(n105223), .B2(DataAddr[6]), 
        .ZN(n99273) );
  OAI21_X1 U89168 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [5]), .B2(n105197), .A(
        n99277), .ZN(\DLX_Datapath/ArithLogUnit/N150 ) );
  AOI22_X1 U89169 ( .A1(n99278), .A2(n105096), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [5]), .ZN(n99277) );
  OAI21_X1 U89170 ( .B1(n99279), .B2(n99280), .A(n107549), .ZN(n99278) );
  AOI21_X1 U89171 ( .B1(n99280), .B2(n99279), .A(n99282), .ZN(n99281) );
  NAND2_X1 U89172 ( .A1(n99283), .A2(n99284), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [5]) );
  AOI21_X1 U89173 ( .B1(n69700), .B2(n105225), .A(n99285), .ZN(n99284) );
  OAI21_X1 U89174 ( .B1(n100643), .B2(n99186), .A(n99286), .ZN(n99285) );
  NAND2_X1 U89175 ( .A1(n72209), .A2(n106929), .ZN(n99286) );
  AOI22_X1 U89176 ( .A1(n99026), .A2(n111077), .B1(n105223), .B2(DataAddr[5]), 
        .ZN(n99283) );
  OAI21_X1 U89177 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [4]), .B2(n105197), .A(
        n99287), .ZN(\DLX_Datapath/ArithLogUnit/N149 ) );
  AOI22_X1 U89178 ( .A1(n99288), .A2(n99289), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [4]), .ZN(n99287) );
  AND2_X2 U89179 ( .A1(n105097), .A2(n99290), .ZN(n99288) );
  NAND2_X1 U89180 ( .A1(n99291), .A2(n99292), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [4]) );
  AOI21_X1 U89181 ( .B1(n69701), .B2(n105225), .A(n99293), .ZN(n99292) );
  OAI21_X1 U89182 ( .B1(n100644), .B2(n99186), .A(n99294), .ZN(n99293) );
  NAND2_X1 U89183 ( .A1(n72065), .A2(n106929), .ZN(n99294) );
  AOI22_X1 U89184 ( .A1(n105224), .A2(n111089), .B1(n105223), .B2(DataAddr[4]), 
        .ZN(n99291) );
  OAI21_X1 U89185 ( .B1(\DLX_Datapath/MUX_HDU_ALUInB [3]), .B2(n105197), .A(
        n99295), .ZN(\DLX_Datapath/ArithLogUnit/N148 ) );
  AOI22_X1 U89186 ( .A1(n99296), .A2(n99297), .B1(n98996), .B2(
        \DLX_Datapath/MUX_HDU_ALUInB [3]), .ZN(n99295) );
  NOR2_X1 U89187 ( .A1(n105899), .A2(n99298), .ZN(n99296) );
  NAND2_X1 U89188 ( .A1(n99299), .A2(n99300), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [3]) );
  AOI21_X1 U89189 ( .B1(n69702), .B2(n105225), .A(n99301), .ZN(n99300) );
  OAI21_X1 U89190 ( .B1(n100645), .B2(n99186), .A(n99302), .ZN(n99301) );
  NAND2_X1 U89191 ( .A1(n71469), .A2(n106929), .ZN(n99302) );
  AOI22_X1 U89192 ( .A1(n99026), .A2(n111084), .B1(n105223), .B2(DataAddr[3]), 
        .ZN(n99299) );
  OAI21_X1 U89193 ( .B1(n106884), .B2(n105227), .A(n99303), .ZN(
        \DLX_Datapath/ArithLogUnit/N147 ) );
  NAND2_X1 U89194 ( .A1(\DLX_Datapath/ArithLogUnit/N177 ), .A2(n106884), .ZN(
        n99303) );
  NAND2_X1 U89195 ( .A1(n99304), .A2(n99305), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [2]) );
  AOI21_X1 U89196 ( .B1(n69703), .B2(n105225), .A(n99306), .ZN(n99305) );
  OAI21_X1 U89197 ( .B1(n100646), .B2(n99186), .A(n99307), .ZN(n99306) );
  NAND2_X1 U89198 ( .A1(n71762), .A2(n106929), .ZN(n99307) );
  AOI22_X1 U89199 ( .A1(n105224), .A2(n111085), .B1(n105223), .B2(DataAddr[2]), 
        .ZN(n99304) );
  OAI21_X1 U89200 ( .B1(n106882), .B2(n105227), .A(n99308), .ZN(
        \DLX_Datapath/ArithLogUnit/N146 ) );
  NAND2_X1 U89201 ( .A1(\DLX_Datapath/ArithLogUnit/N177 ), .A2(n106882), .ZN(
        n99308) );
  NAND2_X1 U89202 ( .A1(n99309), .A2(n99310), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [1]) );
  AOI21_X1 U89203 ( .B1(n69704), .B2(n105225), .A(n99311), .ZN(n99310) );
  OAI21_X1 U89204 ( .B1(n100647), .B2(n99186), .A(n99312), .ZN(n99311) );
  NAND2_X1 U89205 ( .A1(n71618), .A2(n106929), .ZN(n99312) );
  AOI22_X1 U89206 ( .A1(n99026), .A2(n111086), .B1(n105223), .B2(DataAddr[1]), 
        .ZN(n99309) );
  OAI21_X1 U89207 ( .B1(n106768), .B2(n105227), .A(n99313), .ZN(
        \DLX_Datapath/ArithLogUnit/N145 ) );
  NAND2_X1 U89208 ( .A1(\DLX_Datapath/ArithLogUnit/N177 ), .A2(n106768), .ZN(
        n99313) );
  NAND2_X1 U89209 ( .A1(n99314), .A2(n99315), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInB [0]) );
  AOI21_X1 U89210 ( .B1(n69705), .B2(n105225), .A(n99316), .ZN(n99315) );
  OAI21_X1 U89211 ( .B1(n100648), .B2(n99186), .A(n99317), .ZN(n99316) );
  NAND2_X1 U89212 ( .A1(n69292), .A2(n106929), .ZN(n99317) );
  NAND2_X1 U89213 ( .A1(n99318), .A2(n99319), .ZN(n99024) );
  NOR2_X1 U89214 ( .A1(n61539), .A2(n106930), .ZN(n99318) );
  NAND2_X1 U89215 ( .A1(n99320), .A2(n61539), .ZN(n99186) );
  NOR2_X1 U89216 ( .A1(n106930), .A2(n106928), .ZN(n99320) );
  NOR2_X1 U89217 ( .A1(n99321), .A2(n99319), .ZN(n99022) );
  AOI22_X1 U89218 ( .A1(n105224), .A2(n111087), .B1(n105223), .B2(DataAddr[0]), 
        .ZN(n99314) );
  NOR2_X1 U89219 ( .A1(n99321), .A2(n106928), .ZN(n99027) );
  NOR2_X1 U89220 ( .A1(n99319), .A2(n106930), .ZN(n99026) );
  OAI21_X1 U89221 ( .B1(n99322), .B2(n106938), .A(n106931), .ZN(n99321) );
  NOR2_X1 U89222 ( .A1(n83095), .A2(n106935), .ZN(n99322) );
  NAND2_X1 U89223 ( .A1(n99324), .A2(n106931), .ZN(n99319) );
  NOR2_X1 U89224 ( .A1(n99325), .A2(n106938), .ZN(n99324) );
  AOI22_X1 U89225 ( .A1(n99327), .A2(n99328), .B1(n99329), .B2(n99330), .ZN(
        n99326) );
  NOR4_X1 U89226 ( .A1(n99331), .A2(n82682), .A3(n99332), .A4(n99333), .ZN(
        n99330) );
  XOR2_X1 U89227 ( .A(n100420), .B(n100719), .Z(n99333) );
  XOR2_X1 U89228 ( .A(n100418), .B(n62496), .Z(n99332) );
  XNOR2_X1 U89229 ( .A(n99334), .B(n82686), .ZN(n99331) );
  NOR4_X1 U89230 ( .A1(n99335), .A2(n99336), .A3(n99337), .A4(n99338), .ZN(
        n99329) );
  XOR2_X1 U89231 ( .A(n99339), .B(n82689), .Z(n99338) );
  XOR2_X1 U89232 ( .A(n107061), .B(n107103), .Z(n99337) );
  XOR2_X1 U89233 ( .A(n64247), .B(n62662), .Z(n99336) );
  XOR2_X1 U89234 ( .A(n100419), .B(n100427), .Z(n99335) );
  NOR4_X1 U89235 ( .A1(n106939), .A2(n99341), .A3(n99342), .A4(n99343), .ZN(
        n99328) );
  XOR2_X1 U89236 ( .A(n100423), .B(n100719), .Z(n99343) );
  XOR2_X1 U89237 ( .A(n100796), .B(n62496), .Z(n99342) );
  XOR2_X1 U89238 ( .A(n99334), .B(n107102), .Z(n99341) );
  NOR4_X1 U89239 ( .A1(n99345), .A2(n99346), .A3(n99347), .A4(n99348), .ZN(
        n99327) );
  XOR2_X1 U89240 ( .A(n86281), .B(n99339), .Z(n99348) );
  XOR2_X1 U89241 ( .A(n104723), .B(n99349), .Z(n99347) );
  XOR2_X1 U89242 ( .A(n64267), .B(n64247), .Z(n99346) );
  XOR2_X1 U89243 ( .A(n100422), .B(n100427), .Z(n99345) );
  AOI21_X1 U89244 ( .B1(n107062), .B2(n99350), .A(n83106), .ZN(n99325) );
  NOR4_X1 U89246 ( .A1(n99353), .A2(n86273), .A3(n99354), .A4(n99355), .ZN(
        n99352) );
  XOR2_X1 U89247 ( .A(n100894), .B(n64247), .Z(n99355) );
  XOR2_X1 U89248 ( .A(n100427), .B(n54618), .Z(n99354) );
  XOR2_X1 U89249 ( .A(n99334), .B(n86283), .Z(n99353) );
  NOR4_X1 U89250 ( .A1(n99356), .A2(n99357), .A3(n99358), .A4(n99359), .ZN(
        n99351) );
  XOR2_X1 U89251 ( .A(n62496), .B(n54614), .Z(n99359) );
  XOR2_X1 U89252 ( .A(n100719), .B(n54616), .Z(n99358) );
  XOR2_X1 U89253 ( .A(n99339), .B(n86282), .Z(n99357) );
  XOR2_X1 U89254 ( .A(n99349), .B(n86285), .Z(n99356) );
  NAND2_X1 U89255 ( .A1(n99360), .A2(n99361), .ZN(n83095) );
  NOR4_X1 U89256 ( .A1(n99362), .A2(n99363), .A3(n99364), .A4(n99365), .ZN(
        n99361) );
  XOR2_X1 U89257 ( .A(n100427), .B(n100630), .Z(n99365) );
  XOR2_X1 U89258 ( .A(n100631), .B(n100719), .Z(n99364) );
  XOR2_X1 U89259 ( .A(n100632), .B(n62496), .Z(n99363) );
  XOR2_X1 U89260 ( .A(n99334), .B(n86297), .Z(n99362) );
  NOR3_X1 U89261 ( .A1(n99366), .A2(n99367), .A3(n99368), .ZN(n99360) );
  XOR2_X1 U89262 ( .A(n99339), .B(n86296), .Z(n99368) );
  XOR2_X1 U89263 ( .A(n64247), .B(n54620), .Z(n99367) );
  XOR2_X1 U89264 ( .A(n99349), .B(n86295), .Z(n99366) );
  OAI21_X1 U89265 ( .B1(n105196), .B2(n106875), .A(n99369), .ZN(
        \DLX_Datapath/ArithLogUnit/N141 ) );
  NAND2_X1 U89266 ( .A1(n99370), .A2(n105098), .ZN(n99369) );
  XOR2_X1 U89267 ( .A(n99048), .B(n99371), .Z(n99370) );
  XNOR2_X1 U89268 ( .A(n99051), .B(n99049), .ZN(n99371) );
  OAI21_X1 U89269 ( .B1(n99372), .B2(n99373), .A(n107478), .ZN(n99049) );
  AOI21_X1 U89270 ( .B1(n99372), .B2(n99373), .A(n99034), .ZN(n99374) );
  AOI22_X1 U89272 ( .A1(n99015), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] ), .B2(n105122), .ZN(
        n99376) );
  AOI22_X1 U89273 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] ), .A2(
        n108272), .B1(n99016), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .ZN(n99375) );
  XNOR2_X1 U89274 ( .A(n99034), .B(n99377), .ZN(n99048) );
  XNOR2_X1 U89275 ( .A(n99041), .B(n99036), .ZN(n99377) );
  OAI21_X1 U89276 ( .B1(n99378), .B2(n99379), .A(n99380), .ZN(n99036) );
  AOI21_X1 U89277 ( .B1(n99037), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[16] ), .A(n107559), .ZN(
        n99041) );
  AOI21_X1 U89278 ( .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[16] ), .B2(
        n99039), .A(n99040), .ZN(n99381) );
  AOI21_X1 U89279 ( .B1(n99382), .B2(n99383), .A(n108266), .ZN(n99040) );
  NAND2_X1 U89280 ( .A1(n99384), .A2(n99385), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [28]) );
  AOI22_X1 U89281 ( .A1(n98953), .A2(n69711), .B1(n98954), .B2(n111091), .ZN(
        n99385) );
  AOI22_X1 U89282 ( .A1(n105229), .A2(DataAddr[28]), .B1(n98956), .B2(n107852), 
        .ZN(n99384) );
  OAI21_X1 U89283 ( .B1(n105196), .B2(n106874), .A(n99386), .ZN(
        \DLX_Datapath/ArithLogUnit/N140 ) );
  NAND2_X1 U89284 ( .A1(n99387), .A2(n105096), .ZN(n99386) );
  XNOR2_X1 U89286 ( .A(n99061), .B(n99060), .ZN(n99388) );
  NAND2_X1 U89287 ( .A1(n99389), .A2(n99390), .ZN(n99060) );
  AOI22_X1 U89288 ( .A1(n105121), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] ), .B2(n105122), .ZN(
        n99390) );
  AOI22_X1 U89289 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] ), .A2(
        n108272), .B1(n105120), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .ZN(n99389) );
  AOI21_X1 U89290 ( .B1(n99391), .B2(n99392), .A(n107474), .ZN(n99061) );
  OAI21_X1 U89291 ( .B1(n99392), .B2(n99391), .A(n99394), .ZN(n99393) );
  XNOR2_X1 U89292 ( .A(n99034), .B(n99395), .ZN(n99058) );
  XOR2_X1 U89293 ( .A(n99373), .B(n99372), .Z(n99395) );
  OAI21_X1 U89294 ( .B1(n99396), .B2(n99379), .A(n99380), .ZN(n99372) );
  NAND2_X1 U89295 ( .A1(n99397), .A2(n99398), .ZN(n99380) );
  NOR2_X1 U89296 ( .A1(n99398), .A2(n99397), .ZN(n99379) );
  NAND2_X1 U89297 ( .A1(n99399), .A2(n99400), .ZN(n99373) );
  AOI22_X1 U89298 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] ), .B2(n99037), .ZN(
        n99400) );
  AOI22_X1 U89299 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] ), .A2(
        n105119), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99399) );
  XOR2_X1 U89300 ( .A(n99397), .B(n99401), .Z(n99034) );
  XNOR2_X1 U89301 ( .A(n99378), .B(n99398), .ZN(n99401) );
  AOI21_X1 U89302 ( .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[17] ), .B2(
        n99402), .A(n99403), .ZN(n99378) );
  OAI21_X1 U89303 ( .B1(n99404), .B2(n107556), .A(n99405), .ZN(n99403) );
  NAND2_X1 U89304 ( .A1(n99406), .A2(n99407), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [27]) );
  AOI22_X1 U89305 ( .A1(n98953), .A2(n69712), .B1(n98954), .B2(n111092), .ZN(
        n99407) );
  AOI22_X1 U89306 ( .A1(n105229), .A2(DataAddr[27]), .B1(n98956), .B2(n110747), 
        .ZN(n99406) );
  OAI21_X1 U89307 ( .B1(n105196), .B2(n106873), .A(n99408), .ZN(
        \DLX_Datapath/ArithLogUnit/N139 ) );
  NAND2_X1 U89308 ( .A1(n99409), .A2(n105098), .ZN(n99408) );
  XNOR2_X1 U89309 ( .A(n99069), .B(n99410), .ZN(n99409) );
  XOR2_X1 U89310 ( .A(n99071), .B(n99068), .Z(n99410) );
  AOI22_X1 U89312 ( .A1(n99015), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] ), .B2(n105122), .ZN(
        n99412) );
  AOI22_X1 U89313 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] ), .A2(
        n108272), .B1(n99016), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .ZN(n99411) );
  AOI21_X1 U89314 ( .B1(n99413), .B2(n107471), .A(n99414), .ZN(n99071) );
  AOI21_X1 U89315 ( .B1(n99415), .B2(n107506), .A(n99416), .ZN(n99414) );
  XNOR2_X1 U89316 ( .A(n99394), .B(n99417), .ZN(n99069) );
  XNOR2_X1 U89317 ( .A(n99392), .B(n99391), .ZN(n99417) );
  OAI21_X1 U89318 ( .B1(n99418), .B2(n99419), .A(n107475), .ZN(n99391) );
  AOI21_X1 U89319 ( .B1(n99418), .B2(n99419), .A(n99397), .ZN(n99420) );
  AOI22_X1 U89321 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] ), .B2(n99037), .ZN(
        n99422) );
  AOI22_X1 U89322 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] ), .A2(
        n99039), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .ZN(n99421) );
  XNOR2_X1 U89323 ( .A(n99397), .B(n99423), .ZN(n99394) );
  XNOR2_X1 U89324 ( .A(n99396), .B(n99398), .ZN(n99423) );
  OAI21_X1 U89325 ( .B1(n99424), .B2(n99425), .A(n99426), .ZN(n99398) );
  AOI21_X1 U89326 ( .B1(n99402), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[16] ), .A(n99427), .ZN(n99396) );
  OAI21_X1 U89327 ( .B1(n107558), .B2(n99404), .A(n99405), .ZN(n99427) );
  OAI21_X1 U89328 ( .B1(n99428), .B2(n99429), .A(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99405) );
  NAND2_X1 U89329 ( .A1(n99430), .A2(n99431), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [26]) );
  AOI22_X1 U89330 ( .A1(n98953), .A2(n69713), .B1(n98954), .B2(n111093), .ZN(
        n99431) );
  AOI22_X1 U89331 ( .A1(n105229), .A2(DataAddr[26]), .B1(n98956), .B2(n108152), 
        .ZN(n99430) );
  OAI21_X1 U89332 ( .B1(n105196), .B2(n106872), .A(n99432), .ZN(
        \DLX_Datapath/ArithLogUnit/N138 ) );
  NAND2_X1 U89333 ( .A1(n99433), .A2(n105097), .ZN(n99432) );
  XNOR2_X1 U89334 ( .A(n99081), .B(n99434), .ZN(n99433) );
  XOR2_X1 U89335 ( .A(n107465), .B(n107514), .Z(n99434) );
  NAND2_X1 U89336 ( .A1(n99435), .A2(n99436), .ZN(n99080) );
  AOI22_X1 U89337 ( .A1(n105121), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] ), .B2(n105122), .ZN(
        n99436) );
  AOI22_X1 U89338 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] ), .A2(
        n108272), .B1(n99016), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .ZN(n99435) );
  AOI21_X1 U89339 ( .B1(n99437), .B2(n99438), .A(n107466), .ZN(n99078) );
  OAI21_X1 U89340 ( .B1(n99438), .B2(n99437), .A(n99440), .ZN(n99439) );
  XNOR2_X1 U89341 ( .A(n99441), .B(n99416), .ZN(n99081) );
  XNOR2_X1 U89342 ( .A(n99397), .B(n99442), .ZN(n99416) );
  XOR2_X1 U89343 ( .A(n99419), .B(n99418), .Z(n99442) );
  OAI21_X1 U89344 ( .B1(n99443), .B2(n99425), .A(n99426), .ZN(n99418) );
  NAND2_X1 U89345 ( .A1(n99444), .A2(n99445), .ZN(n99426) );
  NOR2_X1 U89346 ( .A1(n99445), .A2(n99444), .ZN(n99425) );
  NAND2_X1 U89347 ( .A1(n99446), .A2(n99447), .ZN(n99419) );
  AOI22_X1 U89348 ( .A1(n105117), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] ), .B2(n105118), .ZN(
        n99447) );
  AOI22_X1 U89349 ( .A1(n105116), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] ), .B2(n108504), .ZN(
        n99446) );
  XOR2_X1 U89350 ( .A(n99444), .B(n99448), .Z(n99397) );
  XNOR2_X1 U89351 ( .A(n99424), .B(n99445), .ZN(n99448) );
  AOI21_X1 U89352 ( .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[17] ), .B2(
        n99449), .A(n99450), .ZN(n99424) );
  OAI21_X1 U89353 ( .B1(n109087), .B2(n107556), .A(n99451), .ZN(n99450) );
  XOR2_X1 U89354 ( .A(n99413), .B(n107471), .Z(n99441) );
  OAI21_X1 U89355 ( .B1(n107472), .B2(n99452), .A(n99453), .ZN(n99415) );
  OAI21_X1 U89356 ( .B1(n107503), .B2(n99454), .A(n99455), .ZN(n99453) );
  NAND2_X1 U89357 ( .A1(n99456), .A2(n99457), .ZN(n99413) );
  AOI22_X1 U89358 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] ), .B2(n99037), .ZN(
        n99457) );
  AOI22_X1 U89359 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] ), .A2(
        n105119), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .ZN(n99456) );
  NAND2_X1 U89360 ( .A1(n99458), .A2(n99459), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [25]) );
  AOI22_X1 U89361 ( .A1(n98953), .A2(n69714), .B1(n98954), .B2(n111094), .ZN(
        n99459) );
  AOI22_X1 U89362 ( .A1(n105229), .A2(DataAddr[25]), .B1(n98956), .B2(n110850), 
        .ZN(n99458) );
  OAI21_X1 U89363 ( .B1(n105196), .B2(n106871), .A(n99460), .ZN(
        \DLX_Datapath/ArithLogUnit/N137 ) );
  NAND2_X1 U89364 ( .A1(n99461), .A2(n105098), .ZN(n99460) );
  XNOR2_X1 U89365 ( .A(n99089), .B(n99462), .ZN(n99461) );
  XOR2_X1 U89366 ( .A(n99091), .B(n99088), .Z(n99462) );
  AOI21_X1 U89367 ( .B1(n99463), .B2(n99464), .A(n107460), .ZN(n99088) );
  OAI21_X1 U89368 ( .B1(n99464), .B2(n99463), .A(n99466), .ZN(n99465) );
  AOI22_X1 U89370 ( .A1(n99015), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] ), .B2(n105122), .ZN(
        n99468) );
  AOI22_X1 U89371 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] ), .A2(
        n108272), .B1(n99016), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .ZN(n99467) );
  XOR2_X1 U89372 ( .A(n99438), .B(n99469), .Z(n99089) );
  XNOR2_X1 U89373 ( .A(n99440), .B(n99437), .ZN(n99469) );
  NAND2_X1 U89374 ( .A1(n99470), .A2(n99471), .ZN(n99437) );
  AOI22_X1 U89375 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] ), .B2(n99037), .ZN(
        n99471) );
  AOI22_X1 U89376 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] ), .A2(
        n105119), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .ZN(n99470) );
  AOI21_X1 U89377 ( .B1(n99472), .B2(n99473), .A(n107467), .ZN(n99440) );
  OAI21_X1 U89378 ( .B1(n99473), .B2(n99472), .A(n99475), .ZN(n99474) );
  XOR2_X1 U89379 ( .A(n99455), .B(n99476), .Z(n99438) );
  XOR2_X1 U89380 ( .A(n107503), .B(n107472), .Z(n99476) );
  OAI21_X1 U89381 ( .B1(n99477), .B2(n99478), .A(n107473), .ZN(n99454) );
  AOI21_X1 U89382 ( .B1(n99477), .B2(n99478), .A(n99444), .ZN(n99479) );
  NAND2_X1 U89383 ( .A1(n99480), .A2(n99481), .ZN(n99452) );
  AOI22_X1 U89384 ( .A1(n99429), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] ), .B2(n105118), .ZN(
        n99481) );
  AOI22_X1 U89385 ( .A1(n105116), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] ), .B2(n108504), .ZN(
        n99480) );
  XNOR2_X1 U89386 ( .A(n99444), .B(n99482), .ZN(n99455) );
  XNOR2_X1 U89387 ( .A(n99443), .B(n99445), .ZN(n99482) );
  OAI21_X1 U89388 ( .B1(n99483), .B2(n99484), .A(n99485), .ZN(n99445) );
  AOI21_X1 U89389 ( .B1(n99449), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[16] ), .A(n99486), .ZN(n99443) );
  OAI21_X1 U89390 ( .B1(n107558), .B2(n109087), .A(n99451), .ZN(n99486) );
  OAI21_X1 U89391 ( .B1(n109088), .B2(n105114), .A(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99451) );
  NAND2_X1 U89392 ( .A1(n99489), .A2(n99490), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [24]) );
  AOI22_X1 U89393 ( .A1(n98953), .A2(n69715), .B1(n98954), .B2(n111095), .ZN(
        n99490) );
  AOI22_X1 U89394 ( .A1(n105229), .A2(DataAddr[24]), .B1(n98956), .B2(n110951), 
        .ZN(n99489) );
  OAI21_X1 U89395 ( .B1(n105196), .B2(n106870), .A(n99491), .ZN(
        \DLX_Datapath/ArithLogUnit/N136 ) );
  NAND2_X1 U89396 ( .A1(n99492), .A2(n105098), .ZN(n99491) );
  XNOR2_X1 U89397 ( .A(n99493), .B(n99098), .ZN(n99492) );
  XOR2_X1 U89398 ( .A(n99464), .B(n99494), .Z(n99098) );
  XNOR2_X1 U89399 ( .A(n99466), .B(n99463), .ZN(n99494) );
  NAND2_X1 U89400 ( .A1(n99495), .A2(n99496), .ZN(n99463) );
  AOI22_X1 U89401 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] ), .B2(n99037), .ZN(
        n99496) );
  AOI22_X1 U89402 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] ), .A2(
        n99039), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .ZN(n99495) );
  AOI21_X1 U89403 ( .B1(n99497), .B2(n99498), .A(n99499), .ZN(n99466) );
  AOI21_X1 U89404 ( .B1(n107464), .B2(n107461), .A(n99500), .ZN(n99499) );
  XNOR2_X1 U89405 ( .A(n99472), .B(n99501), .ZN(n99464) );
  XOR2_X1 U89406 ( .A(n99475), .B(n99473), .Z(n99501) );
  AOI22_X1 U89408 ( .A1(n105117), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] ), .B2(n105118), .ZN(
        n99503) );
  AOI22_X1 U89409 ( .A1(n99428), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] ), .B2(n108504), .ZN(
        n99502) );
  AOI21_X1 U89410 ( .B1(n99504), .B2(n99505), .A(n99506), .ZN(n99475) );
  AOI21_X1 U89411 ( .B1(n107469), .B2(n107504), .A(n99507), .ZN(n99506) );
  XNOR2_X1 U89412 ( .A(n99444), .B(n99508), .ZN(n99472) );
  XOR2_X1 U89413 ( .A(n99478), .B(n99477), .Z(n99508) );
  OAI21_X1 U89414 ( .B1(n99509), .B2(n99484), .A(n99485), .ZN(n99477) );
  NAND2_X1 U89415 ( .A1(n99510), .A2(n99511), .ZN(n99485) );
  NOR2_X1 U89416 ( .A1(n99511), .A2(n99510), .ZN(n99484) );
  NAND2_X1 U89417 ( .A1(n99512), .A2(n99513), .ZN(n99478) );
  AOI22_X1 U89418 ( .A1(n99487), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] ), .B2(n105115), .ZN(
        n99513) );
  AOI22_X1 U89419 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] ), .B2(n99488), .ZN(n99512) );
  XOR2_X1 U89420 ( .A(n99514), .B(n99483), .Z(n99444) );
  AOI21_X1 U89421 ( .B1(n99515), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[17] ), .A(n99516), .ZN(n99483) );
  OAI21_X1 U89422 ( .B1(n107556), .B2(n99517), .A(n99518), .ZN(n99516) );
  AOI21_X1 U89424 ( .B1(n99519), .B2(n107521), .A(n107455), .ZN(n99100) );
  OAI21_X1 U89425 ( .B1(n99519), .B2(n107521), .A(n99521), .ZN(n99520) );
  NAND2_X1 U89426 ( .A1(n99523), .A2(n99524), .ZN(n99101) );
  AOI22_X1 U89427 ( .A1(n105121), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] ), .B2(n105122), .ZN(
        n99524) );
  AOI22_X1 U89428 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] ), .A2(
        n108272), .B1(n105120), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .ZN(n99523) );
  NAND2_X1 U89429 ( .A1(n99525), .A2(n99526), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [23]) );
  AOI22_X1 U89430 ( .A1(n105231), .A2(n69716), .B1(n105230), .B2(n111071), 
        .ZN(n99526) );
  AOI22_X1 U89431 ( .A1(n98955), .A2(DataAddr[23]), .B1(n105228), .B2(n110544), 
        .ZN(n99525) );
  OAI21_X1 U89432 ( .B1(n105196), .B2(n106869), .A(n99527), .ZN(
        \DLX_Datapath/ArithLogUnit/N135 ) );
  NAND2_X1 U89433 ( .A1(n99528), .A2(n105098), .ZN(n99527) );
  XOR2_X1 U89434 ( .A(n99109), .B(n99529), .Z(n99528) );
  XOR2_X1 U89435 ( .A(n99111), .B(n99110), .Z(n99529) );
  NAND2_X1 U89436 ( .A1(n99530), .A2(n99531), .ZN(n99110) );
  AOI22_X1 U89437 ( .A1(n99015), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] ), .B2(n105122), .ZN(
        n99531) );
  AOI22_X1 U89438 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] ), .A2(
        n108272), .B1(n99016), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .ZN(n99530) );
  AOI21_X1 U89439 ( .B1(n99532), .B2(n99533), .A(n107447), .ZN(n99111) );
  OAI21_X1 U89440 ( .B1(n99533), .B2(n99532), .A(n99535), .ZN(n99534) );
  XOR2_X1 U89441 ( .A(n99536), .B(n99521), .Z(n99109) );
  XOR2_X1 U89442 ( .A(n99537), .B(n99498), .Z(n99521) );
  XOR2_X1 U89443 ( .A(n99538), .B(n107469), .Z(n99498) );
  XOR2_X1 U89444 ( .A(n99514), .B(n99509), .Z(n99505) );
  AOI21_X1 U89445 ( .B1(n99515), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[16] ), .A(n99539), .ZN(n99509) );
  OAI21_X1 U89446 ( .B1(n107558), .B2(n99517), .A(n99518), .ZN(n99539) );
  OAI21_X1 U89447 ( .B1(n105110), .B2(n99541), .A(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99518) );
  XNOR2_X1 U89448 ( .A(n99510), .B(n99511), .ZN(n99514) );
  OAI21_X1 U89449 ( .B1(n99542), .B2(n99543), .A(n99544), .ZN(n99511) );
  XOR2_X1 U89450 ( .A(n107504), .B(n99507), .Z(n99538) );
  OAI21_X1 U89451 ( .B1(n99545), .B2(n99546), .A(n107468), .ZN(n99507) );
  AOI21_X1 U89452 ( .B1(n99545), .B2(n99546), .A(n99510), .ZN(n99547) );
  NAND2_X1 U89453 ( .A1(n99548), .A2(n99549), .ZN(n99504) );
  AOI22_X1 U89454 ( .A1(n99487), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] ), .B2(n105115), .ZN(
        n99549) );
  AOI22_X1 U89455 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] ), .B2(n105113), .ZN(
        n99548) );
  XOR2_X1 U89456 ( .A(n99500), .B(n107461), .Z(n99537) );
  OAI21_X1 U89457 ( .B1(n99550), .B2(n99551), .A(n107462), .ZN(n99497) );
  AOI21_X1 U89458 ( .B1(n99551), .B2(n99550), .A(n99553), .ZN(n99552) );
  NAND2_X1 U89459 ( .A1(n99554), .A2(n99555), .ZN(n99500) );
  AOI22_X1 U89460 ( .A1(n99429), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] ), .B2(n105118), .ZN(
        n99555) );
  AOI22_X1 U89461 ( .A1(n99428), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] ), .B2(n108504), .ZN(
        n99554) );
  XOR2_X1 U89462 ( .A(n99522), .B(n99519), .Z(n99536) );
  AOI21_X1 U89463 ( .B1(n99556), .B2(n99557), .A(n107456), .ZN(n99519) );
  OAI21_X1 U89464 ( .B1(n99557), .B2(n99556), .A(n99559), .ZN(n99558) );
  NAND2_X1 U89465 ( .A1(n99560), .A2(n99561), .ZN(n99522) );
  AOI22_X1 U89466 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] ), .B2(n99037), .ZN(
        n99561) );
  AOI22_X1 U89467 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] ), .A2(
        n99039), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .ZN(n99560) );
  NAND2_X1 U89468 ( .A1(n99562), .A2(n99563), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [22]) );
  AOI22_X1 U89469 ( .A1(n105231), .A2(n69717), .B1(n105230), .B2(n111066), 
        .ZN(n99563) );
  AOI22_X1 U89470 ( .A1(n98955), .A2(DataAddr[22]), .B1(n105228), .B2(n110329), 
        .ZN(n99562) );
  OAI21_X1 U89471 ( .B1(n105196), .B2(n106868), .A(n99564), .ZN(
        \DLX_Datapath/ArithLogUnit/N134 ) );
  NAND2_X1 U89472 ( .A1(n99565), .A2(n105098), .ZN(n99564) );
  XOR2_X1 U89473 ( .A(n99119), .B(n99566), .Z(n99565) );
  XOR2_X1 U89474 ( .A(n99120), .B(n99121), .Z(n99566) );
  AOI21_X1 U89475 ( .B1(n99567), .B2(n99568), .A(n107442), .ZN(n99121) );
  OAI21_X1 U89476 ( .B1(n99567), .B2(n99568), .A(n99570), .ZN(n99569) );
  NAND2_X1 U89477 ( .A1(n99571), .A2(n99572), .ZN(n99120) );
  AOI22_X1 U89478 ( .A1(n105121), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] ), .B2(n105122), .ZN(
        n99572) );
  AOI22_X1 U89479 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] ), .A2(
        n108272), .B1(n99016), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .ZN(n99571) );
  XOR2_X1 U89480 ( .A(n99573), .B(n99532), .Z(n99119) );
  XOR2_X1 U89481 ( .A(n99559), .B(n99574), .Z(n99532) );
  XNOR2_X1 U89482 ( .A(n99556), .B(n99557), .ZN(n99574) );
  AOI21_X1 U89483 ( .B1(n99575), .B2(n99576), .A(n107457), .ZN(n99557) );
  OAI21_X1 U89484 ( .B1(n99576), .B2(n99575), .A(n99578), .ZN(n99577) );
  NAND2_X1 U89485 ( .A1(n99579), .A2(n99580), .ZN(n99556) );
  AOI22_X1 U89486 ( .A1(n105117), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] ), .B2(n105118), .ZN(
        n99580) );
  AOI22_X1 U89487 ( .A1(n105116), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] ), .B2(n108504), .ZN(
        n99579) );
  XNOR2_X1 U89488 ( .A(n99553), .B(n99581), .ZN(n99559) );
  XNOR2_X1 U89489 ( .A(n99551), .B(n99550), .ZN(n99581) );
  AOI21_X1 U89490 ( .B1(n99582), .B2(n99583), .A(n107463), .ZN(n99550) );
  OAI21_X1 U89491 ( .B1(n99582), .B2(n99583), .A(n99585), .ZN(n99584) );
  NAND2_X1 U89492 ( .A1(n99586), .A2(n99587), .ZN(n99551) );
  AOI22_X1 U89493 ( .A1(n105114), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] ), .B2(n105115), .ZN(
        n99587) );
  AOI22_X1 U89494 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] ), .B2(n99488), .ZN(n99586) );
  XOR2_X1 U89495 ( .A(n99510), .B(n99588), .Z(n99553) );
  XOR2_X1 U89496 ( .A(n99546), .B(n99545), .Z(n99588) );
  OAI21_X1 U89497 ( .B1(n99542), .B2(n99589), .A(n99544), .ZN(n99545) );
  NAND2_X1 U89498 ( .A1(n99590), .A2(n99591), .ZN(n99546) );
  AOI22_X1 U89499 ( .A1(n105111), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] ), .B2(n105112), .ZN(
        n99591) );
  AOI22_X1 U89500 ( .A1(n99540), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] ), .B2(n109085), .ZN(
        n99590) );
  XOR2_X1 U89501 ( .A(n99592), .B(n99543), .Z(n99510) );
  AOI21_X1 U89502 ( .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[17] ), .B2(
        n108742), .A(n99593), .ZN(n99543) );
  OAI21_X1 U89503 ( .B1(n108744), .B2(n107484), .A(n99594), .ZN(n99593) );
  XNOR2_X1 U89504 ( .A(n99535), .B(n99533), .ZN(n99573) );
  AOI22_X1 U89506 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] ), .B2(n99037), .ZN(n99596) );
  AOI22_X1 U89507 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] ), .A2(
        n105119), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .ZN(n99595) );
  AOI21_X1 U89508 ( .B1(n99597), .B2(n99598), .A(n107448), .ZN(n99535) );
  OAI21_X1 U89509 ( .B1(n99598), .B2(n99597), .A(n99600), .ZN(n99599) );
  NAND2_X1 U89510 ( .A1(n99601), .A2(n99602), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [21]) );
  AOI22_X1 U89511 ( .A1(n105231), .A2(n69718), .B1(n105230), .B2(n111067), 
        .ZN(n99602) );
  AOI22_X1 U89512 ( .A1(n105229), .A2(DataAddr[21]), .B1(n105228), .B2(n110649), .ZN(n99601) );
  OAI21_X1 U89513 ( .B1(n105196), .B2(n106867), .A(n99603), .ZN(
        \DLX_Datapath/ArithLogUnit/N133 ) );
  NAND2_X1 U89514 ( .A1(n99604), .A2(n105096), .ZN(n99603) );
  XOR2_X1 U89515 ( .A(n99130), .B(n99605), .Z(n99604) );
  XOR2_X1 U89516 ( .A(n99131), .B(n107437), .Z(n99605) );
  AOI21_X1 U89517 ( .B1(n99606), .B2(n99607), .A(n107438), .ZN(n99128) );
  OAI21_X1 U89518 ( .B1(n99607), .B2(n99606), .A(n99609), .ZN(n99608) );
  NAND2_X1 U89519 ( .A1(n99610), .A2(n99611), .ZN(n99131) );
  AOI22_X1 U89520 ( .A1(n99015), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] ), .B2(n81819), .ZN(n99611) );
  AOI22_X1 U89521 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] ), .A2(
        n108272), .B1(n105120), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .ZN(n99610) );
  XOR2_X1 U89522 ( .A(n99612), .B(n99570), .Z(n99130) );
  XNOR2_X1 U89523 ( .A(n99598), .B(n99613), .ZN(n99570) );
  XOR2_X1 U89524 ( .A(n99600), .B(n99597), .Z(n99613) );
  NAND2_X1 U89525 ( .A1(n99614), .A2(n99615), .ZN(n99597) );
  AOI22_X1 U89526 ( .A1(n99429), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] ), .B2(n105118), .ZN(
        n99615) );
  AOI22_X1 U89527 ( .A1(n99428), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] ), .B2(n108504), .ZN(
        n99614) );
  OAI21_X1 U89528 ( .B1(n99616), .B2(n99617), .A(n107449), .ZN(n99600) );
  AOI21_X1 U89529 ( .B1(n99617), .B2(n99616), .A(n99619), .ZN(n99618) );
  XOR2_X1 U89530 ( .A(n99620), .B(n99575), .Z(n99598) );
  XNOR2_X1 U89531 ( .A(n99621), .B(n99585), .ZN(n99575) );
  XNOR2_X1 U89532 ( .A(n99592), .B(n99589), .ZN(n99585) );
  AOI21_X1 U89533 ( .B1(n108742), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[16] ), .A(n99622), .ZN(n99589)
         );
  OAI21_X1 U89534 ( .B1(n107490), .B2(n108744), .A(n99594), .ZN(n99622) );
  OAI21_X1 U89535 ( .B1(n99623), .B2(n105107), .A(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99594) );
  XNOR2_X1 U89536 ( .A(n99582), .B(n99583), .ZN(n99621) );
  AOI22_X1 U89538 ( .A1(n99541), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] ), .B2(n105112), .ZN(
        n99627) );
  AOI22_X1 U89539 ( .A1(n99540), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] ), .B2(n109085), .ZN(
        n99626) );
  XNOR2_X1 U89541 ( .A(n99578), .B(n99576), .ZN(n99620) );
  AND2_X2 U89542 ( .A1(n99629), .A2(n99630), .ZN(n99576) );
  AOI22_X1 U89543 ( .A1(n99487), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] ), .B2(n105115), .ZN(
        n99630) );
  AOI22_X1 U89544 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] ), .B2(n105113), .ZN(
        n99629) );
  AOI21_X1 U89545 ( .B1(n99631), .B2(n99632), .A(n99633), .ZN(n99578) );
  XNOR2_X1 U89547 ( .A(n99568), .B(n99567), .ZN(n99612) );
  AOI22_X1 U89549 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] ), .B2(n99037), .ZN(n99636) );
  AOI22_X1 U89550 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] ), .A2(
        n99039), .B1(n107737), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .ZN(n99635) );
  AOI21_X1 U89551 ( .B1(n99637), .B2(n99638), .A(n107443), .ZN(n99568) );
  OAI21_X1 U89552 ( .B1(n99638), .B2(n99637), .A(n99640), .ZN(n99639) );
  NAND2_X1 U89553 ( .A1(n99641), .A2(n99642), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [20]) );
  AOI22_X1 U89554 ( .A1(n105231), .A2(n69719), .B1(n105230), .B2(n111068), 
        .ZN(n99642) );
  AOI22_X1 U89555 ( .A1(n105229), .A2(DataAddr[20]), .B1(n105228), .B2(n110438), .ZN(n99641) );
  OAI21_X1 U89556 ( .B1(n105196), .B2(n106866), .A(n99643), .ZN(
        \DLX_Datapath/ArithLogUnit/N132 ) );
  NAND2_X1 U89557 ( .A1(n99644), .A2(n105096), .ZN(n99643) );
  XOR2_X1 U89558 ( .A(n99645), .B(n99140), .Z(n99644) );
  XNOR2_X1 U89559 ( .A(n99607), .B(n99646), .ZN(n99140) );
  XNOR2_X1 U89560 ( .A(n99609), .B(n99606), .ZN(n99646) );
  NAND2_X1 U89561 ( .A1(n99647), .A2(n99648), .ZN(n99606) );
  AOI22_X1 U89562 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] ), .B2(n99037), .ZN(n99648) );
  AOI22_X1 U89563 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] ), .A2(
        n105119), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .ZN(n99647) );
  AOI21_X1 U89565 ( .B1(n99650), .B2(n99651), .A(n99652), .ZN(n99649) );
  XOR2_X1 U89566 ( .A(n99653), .B(n99638), .Z(n99607) );
  XOR2_X1 U89567 ( .A(n99654), .B(n99617), .Z(n99638) );
  XOR2_X1 U89568 ( .A(n99632), .B(n99655), .Z(n99617) );
  XOR2_X1 U89569 ( .A(n99634), .B(n99631), .Z(n99655) );
  NAND2_X1 U89570 ( .A1(n99656), .A2(n99657), .ZN(n99631) );
  AOI22_X1 U89571 ( .A1(n105111), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] ), .B2(n105112), .ZN(
        n99657) );
  AOI22_X1 U89572 ( .A1(n105110), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] ), .B2(n109085), .ZN(
        n99656) );
  OAI21_X1 U89573 ( .B1(n99658), .B2(n99659), .A(n107483), .ZN(n99634) );
  AOI21_X1 U89574 ( .B1(n99658), .B2(n99659), .A(n99661), .ZN(n99660) );
  XNOR2_X1 U89575 ( .A(n99592), .B(n99628), .ZN(n99632) );
  NAND2_X1 U89576 ( .A1(n99662), .A2(n99663), .ZN(n99628) );
  AOI22_X1 U89577 ( .A1(n105108), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] ), .B2(n105109), .ZN(
        n99663) );
  AOI22_X1 U89578 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] ), .A2(
        n108742), .B1(n105107), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99662) );
  NAND2_X1 U89579 ( .A1(n107482), .A2(n99544), .ZN(n99592) );
  NAND2_X1 U89580 ( .A1(n99664), .A2(n99661), .ZN(n99544) );
  NOR2_X1 U89581 ( .A1(n99661), .A2(n99664), .ZN(n99542) );
  OAI21_X1 U89582 ( .B1(n107556), .B2(n99665), .A(n99666), .ZN(n99664) );
  AOI21_X1 U89583 ( .B1(n99667), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[17] ), .A(n108268), .ZN(
        n99666) );
  XNOR2_X1 U89584 ( .A(n99616), .B(n99619), .ZN(n99654) );
  AOI21_X1 U89585 ( .B1(n99668), .B2(n107450), .A(n99669), .ZN(n99619) );
  AOI21_X1 U89586 ( .B1(n99670), .B2(n107510), .A(n99671), .ZN(n99669) );
  AOI22_X1 U89588 ( .A1(n99487), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] ), .B2(n105115), .ZN(
        n99673) );
  AOI22_X1 U89589 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] ), .B2(n99488), .ZN(n99672) );
  XOR2_X1 U89590 ( .A(n99640), .B(n99637), .Z(n99653) );
  NAND2_X1 U89591 ( .A1(n99674), .A2(n99675), .ZN(n99637) );
  AOI22_X1 U89592 ( .A1(n105117), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] ), .B2(n105118), .ZN(
        n99675) );
  AOI22_X1 U89593 ( .A1(n105116), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] ), .B2(n108504), .ZN(n99674) );
  AOI21_X1 U89594 ( .B1(n107444), .B2(n99676), .A(n99677), .ZN(n99640) );
  AOI21_X1 U89595 ( .B1(n107451), .B2(n99678), .A(n99679), .ZN(n99677) );
  XOR2_X1 U89596 ( .A(n107434), .B(n99141), .Z(n99645) );
  NAND2_X1 U89597 ( .A1(n99680), .A2(n99681), .ZN(n99141) );
  AOI22_X1 U89598 ( .A1(n105121), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] ), .B2(n81819), .ZN(n99681) );
  AOI22_X1 U89599 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] ), .A2(
        n108272), .B1(n105120), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .ZN(n99680) );
  OAI21_X1 U89600 ( .B1(n99682), .B2(n99683), .A(n99684), .ZN(n99138) );
  OAI21_X1 U89601 ( .B1(n107540), .B2(n107439), .A(n99685), .ZN(n99684) );
  NAND2_X1 U89602 ( .A1(n99686), .A2(n99687), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [19]) );
  AOI22_X1 U89603 ( .A1(n105231), .A2(n69720), .B1(n105230), .B2(n111072), 
        .ZN(n99687) );
  AOI22_X1 U89604 ( .A1(n105229), .A2(DataAddr[19]), .B1(n105228), .B2(n110116), .ZN(n99686) );
  OAI21_X1 U89605 ( .B1(n105196), .B2(n106865), .A(n99688), .ZN(
        \DLX_Datapath/ArithLogUnit/N131 ) );
  NAND2_X1 U89606 ( .A1(n99689), .A2(n105098), .ZN(n99688) );
  XNOR2_X1 U89607 ( .A(n99148), .B(n99690), .ZN(n99689) );
  XOR2_X1 U89608 ( .A(n99149), .B(n99151), .Z(n99690) );
  AOI22_X1 U89610 ( .A1(n99015), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] ), .B2(n81819), .ZN(n99692) );
  AOI22_X1 U89611 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] ), .A2(
        n108272), .B1(n105120), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .ZN(n99691) );
  OAI21_X1 U89612 ( .B1(n99693), .B2(n99694), .A(n107433), .ZN(n99149) );
  AOI21_X1 U89613 ( .B1(n99694), .B2(n99693), .A(n99696), .ZN(n99695) );
  XOR2_X1 U89614 ( .A(n99682), .B(n99697), .Z(n99148) );
  XOR2_X1 U89615 ( .A(n99685), .B(n99683), .Z(n99697) );
  NAND2_X1 U89616 ( .A1(n99698), .A2(n99699), .ZN(n99683) );
  AOI22_X1 U89617 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] ), .B2(n99037), .ZN(n99699) );
  AOI22_X1 U89618 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] ), .A2(
        n105119), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .ZN(n99698) );
  OAI21_X1 U89619 ( .B1(n99700), .B2(n99701), .A(n107435), .ZN(n99685) );
  AOI21_X1 U89620 ( .B1(n99701), .B2(n99700), .A(n99703), .ZN(n99702) );
  XOR2_X1 U89621 ( .A(n99704), .B(n99650), .Z(n99682) );
  XOR2_X1 U89622 ( .A(n99676), .B(n99705), .Z(n99650) );
  XOR2_X1 U89623 ( .A(n99679), .B(n107444), .Z(n99705) );
  AOI21_X1 U89624 ( .B1(n99706), .B2(n99707), .A(n107445), .ZN(n99678) );
  OAI21_X1 U89625 ( .B1(n99707), .B2(n99706), .A(n99709), .ZN(n99708) );
  NAND2_X1 U89626 ( .A1(n99710), .A2(n99711), .ZN(n99679) );
  AOI22_X1 U89627 ( .A1(n105114), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] ), .B2(n105115), .ZN(
        n99711) );
  AOI22_X1 U89628 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] ), .B2(n105113), .ZN(
        n99710) );
  XOR2_X1 U89629 ( .A(n99712), .B(n99671), .Z(n99676) );
  XOR2_X1 U89630 ( .A(n99713), .B(n99658), .Z(n99671) );
  NAND2_X1 U89631 ( .A1(n99714), .A2(n99715), .ZN(n99658) );
  AOI22_X1 U89632 ( .A1(n99623), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] ), .B2(n105109), .ZN(
        n99715) );
  AOI22_X1 U89633 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] ), .A2(
        n108742), .B1(n105107), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .ZN(n99714) );
  XNOR2_X1 U89634 ( .A(n99659), .B(n99661), .ZN(n99713) );
  OAI21_X1 U89635 ( .B1(n99665), .B2(n107558), .A(n99716), .ZN(n99659) );
  AOI21_X1 U89636 ( .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[16] ), .B2(
        n99667), .A(n108268), .ZN(n99716) );
  OAI21_X1 U89637 ( .B1(n99718), .B2(n105104), .A(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99717) );
  XOR2_X1 U89638 ( .A(n99670), .B(n107510), .Z(n99712) );
  NAND2_X1 U89639 ( .A1(n99720), .A2(n99721), .ZN(n99668) );
  AOI22_X1 U89640 ( .A1(n99541), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] ), .B2(n105112), .ZN(
        n99721) );
  AOI22_X1 U89641 ( .A1(n99540), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] ), .B2(n109085), .ZN(
        n99720) );
  OAI21_X1 U89642 ( .B1(n99722), .B2(n99723), .A(n107452), .ZN(n99670) );
  AOI21_X1 U89643 ( .B1(n99722), .B2(n99723), .A(n99661), .ZN(n99724) );
  XOR2_X1 U89644 ( .A(n99651), .B(n99652), .Z(n99704) );
  NAND2_X1 U89645 ( .A1(n99725), .A2(n99726), .ZN(n99652) );
  AOI22_X1 U89646 ( .A1(n99429), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] ), .B2(n105118), .ZN(
        n99726) );
  AOI22_X1 U89647 ( .A1(n105116), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] ), .B2(n108504), .ZN(n99725) );
  AOI21_X1 U89648 ( .B1(n99727), .B2(n99728), .A(n107440), .ZN(n99651) );
  OAI21_X1 U89649 ( .B1(n99728), .B2(n99727), .A(n99730), .ZN(n99729) );
  NAND2_X1 U89650 ( .A1(n99731), .A2(n99732), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [18]) );
  AOI22_X1 U89651 ( .A1(n105231), .A2(n69721), .B1(n105230), .B2(n111073), 
        .ZN(n99732) );
  AOI22_X1 U89652 ( .A1(n105229), .A2(DataAddr[18]), .B1(n105228), .B2(n110223), .ZN(n99731) );
  OAI21_X1 U89653 ( .B1(n105196), .B2(n106864), .A(n99733), .ZN(
        \DLX_Datapath/ArithLogUnit/N130 ) );
  NAND2_X1 U89654 ( .A1(n99734), .A2(n105096), .ZN(n99733) );
  XOR2_X1 U89655 ( .A(n99159), .B(n99735), .Z(n99734) );
  AOI22_X1 U89658 ( .A1(n105121), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] ), .B2(n81819), .ZN(n99737) );
  AOI22_X1 U89659 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] ), .A2(
        n108272), .B1(n105120), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .ZN(n99736) );
  OAI21_X1 U89660 ( .B1(n99738), .B2(n99739), .A(n99740), .ZN(n99161) );
  OAI21_X1 U89661 ( .B1(n107545), .B2(n107486), .A(n99741), .ZN(n99740) );
  XOR2_X1 U89662 ( .A(n99742), .B(n99693), .Z(n99159) );
  XNOR2_X1 U89663 ( .A(n99703), .B(n99743), .ZN(n99693) );
  XNOR2_X1 U89664 ( .A(n99700), .B(n99701), .ZN(n99743) );
  NAND2_X1 U89665 ( .A1(n99744), .A2(n99745), .ZN(n99701) );
  AOI22_X1 U89666 ( .A1(n105117), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] ), .B2(n105118), .ZN(
        n99745) );
  AOI22_X1 U89667 ( .A1(n99428), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] ), .B2(n108504), .ZN(n99744) );
  AOI21_X1 U89668 ( .B1(n99746), .B2(n99747), .A(n107488), .ZN(n99700) );
  OAI21_X1 U89669 ( .B1(n99747), .B2(n99746), .A(n99749), .ZN(n99748) );
  XNOR2_X1 U89670 ( .A(n99727), .B(n99750), .ZN(n99703) );
  XOR2_X1 U89671 ( .A(n99730), .B(n99728), .Z(n99750) );
  AOI22_X1 U89673 ( .A1(n99487), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] ), .B2(n105115), .ZN(
        n99752) );
  AOI22_X1 U89674 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] ), .B2(n99488), .ZN(n99751)
         );
  AOI21_X1 U89675 ( .B1(n99753), .B2(n107496), .A(n99754), .ZN(n99730) );
  AOI21_X1 U89676 ( .B1(n99755), .B2(n107522), .A(n99756), .ZN(n99754) );
  XOR2_X1 U89677 ( .A(n99757), .B(n99709), .Z(n99727) );
  XOR2_X1 U89678 ( .A(n99758), .B(n99722), .Z(n99709) );
  NAND2_X1 U89679 ( .A1(n99759), .A2(n99760), .ZN(n99722) );
  AOI22_X1 U89680 ( .A1(n105108), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] ), .B2(n105109), .ZN(
        n99760) );
  AOI22_X1 U89681 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] ), .A2(
        n108742), .B1(n105107), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .ZN(n99759) );
  XNOR2_X1 U89682 ( .A(n99661), .B(n99723), .ZN(n99758) );
  NAND2_X1 U89683 ( .A1(n99761), .A2(n99762), .ZN(n99723) );
  AOI22_X1 U89684 ( .A1(n105105), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] ), .B2(n105106), .ZN(
        n99762) );
  AOI22_X1 U89685 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] ), .A2(
        n108741), .B1(n99719), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(n99761) );
  OAI21_X1 U89686 ( .B1(n107484), .B2(n107570), .A(n99763), .ZN(n99661) );
  AOI21_X1 U89687 ( .B1(n99764), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[17] ), .A(n99765), .ZN(n99763)
         );
  XOR2_X1 U89688 ( .A(n99706), .B(n99707), .Z(n99757) );
  AOI22_X1 U89690 ( .A1(n105111), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] ), .B2(n105112), .ZN(
        n99767) );
  AOI22_X1 U89691 ( .A1(n105110), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] ), .B2(n109085), .ZN(
        n99766) );
  OAI21_X1 U89692 ( .B1(n99768), .B2(n99769), .A(n107489), .ZN(n99706) );
  AOI21_X1 U89693 ( .B1(n99768), .B2(n99769), .A(n99771), .ZN(n99770) );
  XNOR2_X1 U89694 ( .A(n99696), .B(n99694), .ZN(n99742) );
  NAND2_X1 U89695 ( .A1(n99772), .A2(n99773), .ZN(n99694) );
  AOI22_X1 U89696 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] ), .B2(n99037), .ZN(n99773) );
  AOI22_X1 U89697 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] ), .A2(
        n99039), .B1(n107737), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .ZN(n99772) );
  OAI21_X1 U89698 ( .B1(n99774), .B2(n99775), .A(n107487), .ZN(n99696) );
  AOI21_X1 U89699 ( .B1(n99775), .B2(n99774), .A(n99777), .ZN(n99776) );
  NAND2_X1 U89700 ( .A1(n99778), .A2(n99779), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [17]) );
  AOI22_X1 U89701 ( .A1(n105231), .A2(n69722), .B1(n105230), .B2(n111078), 
        .ZN(n99779) );
  AOI22_X1 U89702 ( .A1(n105229), .A2(DataAddr[17]), .B1(n105228), .B2(n110008), .ZN(n99778) );
  OAI21_X1 U89703 ( .B1(n106945), .B2(n106863), .A(n99780), .ZN(
        \DLX_Datapath/ArithLogUnit/N129 ) );
  NAND2_X1 U89704 ( .A1(n99781), .A2(n105096), .ZN(n99780) );
  XNOR2_X1 U89705 ( .A(n99169), .B(n99782), .ZN(n99781) );
  XOR2_X1 U89706 ( .A(n99171), .B(n107552), .Z(n99782) );
  NAND2_X1 U89707 ( .A1(n99783), .A2(n99784), .ZN(n99170) );
  AOI22_X1 U89708 ( .A1(n99015), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] ), .B2(n81819), .ZN(n99784) );
  AOI22_X1 U89709 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] ), .A2(
        n108272), .B1(n105120), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .ZN(n99783) );
  AOI21_X1 U89710 ( .B1(n99785), .B2(n99786), .A(n107493), .ZN(n99171) );
  OAI21_X1 U89711 ( .B1(n99786), .B2(n99785), .A(n99788), .ZN(n99787) );
  XOR2_X1 U89712 ( .A(n107486), .B(n99789), .Z(n99169) );
  XOR2_X1 U89713 ( .A(n99741), .B(n99739), .Z(n99789) );
  NAND2_X1 U89714 ( .A1(n99790), .A2(n99791), .ZN(n99739) );
  AOI22_X1 U89715 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] ), .B2(n99037), .ZN(n99791) );
  AOI22_X1 U89716 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] ), .A2(
        n99039), .B1(n107737), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .ZN(n99790) );
  OAI21_X1 U89717 ( .B1(n99792), .B2(n99793), .A(n107494), .ZN(n99741) );
  AOI21_X1 U89718 ( .B1(n99793), .B2(n99792), .A(n99795), .ZN(n99794) );
  XOR2_X1 U89719 ( .A(n99796), .B(n99775), .Z(n99738) );
  XNOR2_X1 U89720 ( .A(n99797), .B(n99746), .ZN(n99775) );
  XOR2_X1 U89721 ( .A(n99798), .B(n99756), .Z(n99746) );
  XOR2_X1 U89722 ( .A(n99799), .B(n99768), .Z(n99756) );
  NAND2_X1 U89723 ( .A1(n99800), .A2(n99801), .ZN(n99768) );
  AOI22_X1 U89724 ( .A1(n99623), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] ), .B2(n105109), .ZN(
        n99801) );
  AOI22_X1 U89725 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] ), .A2(
        n108742), .B1(n105107), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .ZN(n99800) );
  XNOR2_X1 U89726 ( .A(n99771), .B(n99769), .ZN(n99799) );
  NAND2_X1 U89727 ( .A1(n99802), .A2(n99803), .ZN(n99769) );
  AOI22_X1 U89728 ( .A1(n99718), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] ), .B2(n105106), .ZN(
        n99803) );
  AOI22_X1 U89729 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] ), .A2(
        n108741), .B1(n105104), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .ZN(n99802) );
  OAI21_X1 U89730 ( .B1(n107570), .B2(n107490), .A(n99804), .ZN(n99771) );
  AOI21_X1 U89731 ( .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[16] ), .B2(
        n99764), .A(n99765), .ZN(n99804) );
  XOR2_X1 U89732 ( .A(n99755), .B(n107522), .Z(n99798) );
  NAND2_X1 U89733 ( .A1(n99805), .A2(n99806), .ZN(n99753) );
  AOI22_X1 U89734 ( .A1(n99541), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] ), .B2(n105112), .ZN(
        n99806) );
  AOI22_X1 U89735 ( .A1(n105110), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] ), .B2(n109085), .ZN(
        n99805) );
  OAI21_X1 U89736 ( .B1(n99807), .B2(n99808), .A(n99809), .ZN(n99755) );
  OAI21_X1 U89737 ( .B1(n107515), .B2(n107507), .A(n99810), .ZN(n99809) );
  XNOR2_X1 U89738 ( .A(n99749), .B(n99747), .ZN(n99797) );
  AOI22_X1 U89740 ( .A1(n105114), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] ), .B2(n105115), .ZN(
        n99812) );
  AOI22_X1 U89741 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] ), .B2(n105113), .ZN(n99811) );
  AOI21_X1 U89742 ( .B1(n99813), .B2(n99814), .A(n99815), .ZN(n99749) );
  XNOR2_X1 U89744 ( .A(n99774), .B(n99777), .ZN(n99796) );
  AOI22_X1 U89746 ( .A1(n99429), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] ), .B2(n99402), .ZN(n99818) );
  AOI22_X1 U89747 ( .A1(n99428), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] ), .B2(n108504), .ZN(n99817) );
  AOI21_X1 U89748 ( .B1(n99819), .B2(n99820), .A(n107495), .ZN(n99774) );
  OAI21_X1 U89749 ( .B1(n99820), .B2(n99819), .A(n99822), .ZN(n99821) );
  NAND2_X1 U89750 ( .A1(n99823), .A2(n99824), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [16]) );
  AOI22_X1 U89751 ( .A1(n105231), .A2(n69723), .B1(n105230), .B2(n111074), 
        .ZN(n99824) );
  AOI22_X1 U89752 ( .A1(n105229), .A2(DataAddr[16]), .B1(n105228), .B2(n109891), .ZN(n99823) );
  OAI21_X1 U89753 ( .B1(n106945), .B2(n106862), .A(n99825), .ZN(
        \DLX_Datapath/ArithLogUnit/N128 ) );
  NAND2_X1 U89754 ( .A1(n99826), .A2(n105098), .ZN(n99825) );
  XNOR2_X1 U89755 ( .A(n99827), .B(n99178), .ZN(n99826) );
  XOR2_X1 U89756 ( .A(n99785), .B(n99828), .Z(n99178) );
  XOR2_X1 U89757 ( .A(n99788), .B(n99786), .Z(n99828) );
  AOI22_X1 U89759 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] ), .B2(n99037), .ZN(n99830) );
  AOI22_X1 U89760 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] ), .A2(
        n105119), .B1(n107737), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .ZN(n99829) );
  AOI21_X1 U89761 ( .B1(n99831), .B2(n99832), .A(n107498), .ZN(n99788) );
  OAI21_X1 U89762 ( .B1(n99832), .B2(n99831), .A(n99834), .ZN(n99833) );
  XOR2_X1 U89763 ( .A(n99835), .B(n99792), .Z(n99785) );
  XOR2_X1 U89764 ( .A(n99820), .B(n99836), .Z(n99792) );
  XOR2_X1 U89765 ( .A(n99822), .B(n99819), .Z(n99836) );
  NAND2_X1 U89766 ( .A1(n99837), .A2(n99838), .ZN(n99819) );
  AOI22_X1 U89767 ( .A1(n105114), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] ), .B2(n105115), .ZN(
        n99838) );
  AOI22_X1 U89768 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] ), .B2(n105113), .ZN(n99837) );
  OAI21_X1 U89769 ( .B1(n99839), .B2(n99840), .A(n107500), .ZN(n99822) );
  AOI21_X1 U89770 ( .B1(n99840), .B2(n99839), .A(n99842), .ZN(n99841) );
  XOR2_X1 U89771 ( .A(n99843), .B(n99814), .Z(n99820) );
  XOR2_X1 U89772 ( .A(n99844), .B(n107515), .Z(n99814) );
  NAND2_X1 U89773 ( .A1(n99845), .A2(n99846), .ZN(n99807) );
  AOI22_X1 U89774 ( .A1(n105108), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] ), .B2(n105109), .ZN(
        n99846) );
  AOI22_X1 U89775 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] ), .A2(
        n108742), .B1(n105107), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .ZN(n99845) );
  XOR2_X1 U89776 ( .A(n99810), .B(n99808), .Z(n99844) );
  NAND2_X1 U89777 ( .A1(n99847), .A2(n99848), .ZN(n99808) );
  AOI22_X1 U89778 ( .A1(n105105), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] ), .B2(n105106), .ZN(
        n99848) );
  AOI22_X1 U89779 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] ), .A2(
        n108741), .B1(n99719), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .ZN(n99847) );
  AOI21_X1 U89780 ( .B1(n105102), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] ), .A(n107560), .ZN(
        n99810) );
  AOI21_X1 U89781 ( .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] ), .B2(
        n99764), .A(n99765), .ZN(n99850) );
  NOR2_X1 U89782 ( .A1(n99851), .A2(n108266), .ZN(n99765) );
  XNOR2_X1 U89783 ( .A(n99816), .B(n99813), .ZN(n99843) );
  NAND2_X1 U89784 ( .A1(n99852), .A2(n99853), .ZN(n99813) );
  AOI22_X1 U89785 ( .A1(n105111), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] ), .B2(n105112), .ZN(
        n99853) );
  AOI22_X1 U89786 ( .A1(n99540), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] ), .B2(n109085), .ZN(n99852) );
  OAI21_X1 U89787 ( .B1(n99854), .B2(n99855), .A(n107501), .ZN(n99816) );
  AOI21_X1 U89788 ( .B1(n99854), .B2(n99855), .A(n99857), .ZN(n99856) );
  XNOR2_X1 U89789 ( .A(n99793), .B(n99795), .ZN(n99835) );
  NAND2_X1 U89790 ( .A1(n99858), .A2(n99859), .ZN(n99795) );
  AOI22_X1 U89791 ( .A1(n105117), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] ), .B2(n99402), .ZN(n99859) );
  AOI22_X1 U89792 ( .A1(n105116), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] ), .B2(n108504), .ZN(n99858) );
  OAI21_X1 U89793 ( .B1(n99860), .B2(n99861), .A(n107499), .ZN(n99793) );
  AOI21_X1 U89794 ( .B1(n99861), .B2(n99860), .A(n99863), .ZN(n99862) );
  NAND2_X1 U89796 ( .A1(n99864), .A2(n99865), .ZN(n99180) );
  AOI22_X1 U89797 ( .A1(n105121), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[1] ), .B2(n81819), .ZN(n99865) );
  NOR2_X1 U89798 ( .A1(n99866), .A2(n108273), .ZN(n81819) );
  NOR2_X1 U89799 ( .A1(n99867), .A2(n108271), .ZN(n99015) );
  AOI22_X1 U89800 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] ), .A2(
        n108272), .B1(n105120), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .ZN(n99864) );
  AOI21_X1 U89801 ( .B1(n99869), .B2(n99870), .A(n107497), .ZN(n99181) );
  OAI21_X1 U89802 ( .B1(n99870), .B2(n99869), .A(n99872), .ZN(n99871) );
  NAND2_X1 U89803 ( .A1(n99873), .A2(n99874), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [15]) );
  AOI22_X1 U89804 ( .A1(n105231), .A2(n69724), .B1(n105230), .B2(n111096), 
        .ZN(n99874) );
  AOI22_X1 U89805 ( .A1(n105229), .A2(DataAddr[15]), .B1(n105228), .B2(n108265), .ZN(n99873) );
  OAI21_X1 U89806 ( .B1(n106945), .B2(n106861), .A(n99875), .ZN(
        \DLX_Datapath/ArithLogUnit/N127 ) );
  NAND2_X1 U89807 ( .A1(n99876), .A2(n105098), .ZN(n99875) );
  XOR2_X1 U89808 ( .A(n99190), .B(n99189), .Z(n99876) );
  XNOR2_X1 U89809 ( .A(n99869), .B(n99877), .ZN(n99189) );
  XOR2_X1 U89810 ( .A(n99872), .B(n99870), .Z(n99877) );
  AOI22_X1 U89812 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] ), .B2(n99037), .ZN(n99879) );
  AOI22_X1 U89813 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] ), .A2(
        n99039), .B1(n107737), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .ZN(n99878) );
  AOI21_X1 U89814 ( .B1(n99880), .B2(n99881), .A(n107508), .ZN(n99872) );
  OAI21_X1 U89815 ( .B1(n99881), .B2(n99880), .A(n99883), .ZN(n99882) );
  XOR2_X1 U89816 ( .A(n99884), .B(n99832), .Z(n99869) );
  XNOR2_X1 U89817 ( .A(n99861), .B(n99885), .ZN(n99832) );
  XOR2_X1 U89818 ( .A(n99863), .B(n99860), .Z(n99885) );
  AOI22_X1 U89820 ( .A1(n99487), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] ), .B2(n99449), .ZN(n99887) );
  AOI22_X1 U89821 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] ), .B2(n105113), .ZN(n99886) );
  AOI21_X1 U89822 ( .B1(n99888), .B2(n107513), .A(n99889), .ZN(n99863) );
  AOI21_X1 U89823 ( .B1(n99890), .B2(n107536), .A(n99891), .ZN(n99889) );
  XOR2_X1 U89824 ( .A(n99892), .B(n99842), .Z(n99861) );
  XOR2_X1 U89825 ( .A(n99893), .B(n99854), .Z(n99842) );
  NAND2_X1 U89826 ( .A1(n99894), .A2(n99895), .ZN(n99854) );
  AOI22_X1 U89827 ( .A1(n99718), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] ), .B2(n105106), .ZN(
        n99895) );
  AOI22_X1 U89828 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] ), .A2(
        n108741), .B1(n105104), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .ZN(n99894) );
  XNOR2_X1 U89829 ( .A(n99857), .B(n99855), .ZN(n99893) );
  NAND2_X1 U89830 ( .A1(n99896), .A2(n99897), .ZN(n99855) );
  AOI22_X1 U89831 ( .A1(n99623), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] ), .B2(n105109), .ZN(
        n99897) );
  AOI22_X1 U89832 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] ), .A2(
        n108742), .B1(n105107), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .ZN(n99896) );
  OAI21_X1 U89833 ( .B1(n107570), .B2(n107502), .A(n99898), .ZN(n99857) );
  AOI22_X1 U89834 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] ), .A2(
        n99764), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .ZN(n99898) );
  XOR2_X1 U89835 ( .A(n99840), .B(n99839), .Z(n99892) );
  AOI22_X1 U89837 ( .A1(n99541), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] ), .B2(n105112), .ZN(
        n99900) );
  AOI22_X1 U89838 ( .A1(n99540), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] ), .B2(n109085), .ZN(n99899) );
  OAI21_X1 U89839 ( .B1(n99901), .B2(n99902), .A(n99903), .ZN(n99840) );
  OAI21_X1 U89840 ( .B1(n107516), .B2(n107526), .A(n99904), .ZN(n99903) );
  XNOR2_X1 U89841 ( .A(n99831), .B(n99834), .ZN(n99884) );
  NAND2_X1 U89842 ( .A1(n99905), .A2(n99906), .ZN(n99834) );
  AOI22_X1 U89843 ( .A1(n99429), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] ), .B2(n99402), .ZN(n99906) );
  AOI22_X1 U89844 ( .A1(n99428), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] ), .B2(n108504), .ZN(n99905) );
  OAI21_X1 U89845 ( .B1(n99907), .B2(n99908), .A(n107509), .ZN(n99831) );
  AOI21_X1 U89846 ( .B1(n99908), .B2(n99907), .A(n99910), .ZN(n99909) );
  OAI21_X1 U89847 ( .B1(n81817), .B2(n107568), .A(n99911), .ZN(n99190) );
  NAND2_X1 U89848 ( .A1(n105120), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .ZN(n99911) );
  NOR2_X1 U89849 ( .A1(n99868), .A2(n99867), .ZN(n99016) );
  NAND2_X1 U89850 ( .A1(n99868), .A2(n99867), .ZN(n81817) );
  NAND2_X1 U89851 ( .A1(n99866), .A2(n108273), .ZN(n99867) );
  OR2_X1 U89852 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [14]), .A2(
        \DLX_Datapath/ArithLogUnit/B_mul [13]), .ZN(n99866) );
  OAI21_X1 U89853 ( .B1(n108392), .B2(n99912), .A(n99913), .ZN(n99868) );
  NAND2_X1 U89854 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [15]), .A2(n99914), 
        .ZN(n99913) );
  XOR2_X1 U89855 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [14]), .B(
        \DLX_Datapath/ArithLogUnit/B_mul [13]), .Z(n99914) );
  NAND2_X1 U89856 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [13]), .A2(n108273), 
        .ZN(n99912) );
  NAND2_X1 U89857 ( .A1(n99915), .A2(n99916), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [14]) );
  AOI22_X1 U89858 ( .A1(n105231), .A2(n69725), .B1(n105230), .B2(n111079), 
        .ZN(n99916) );
  AOI22_X1 U89859 ( .A1(n105229), .A2(DataAddr[14]), .B1(n105228), .B2(n108388), .ZN(n99915) );
  OAI21_X1 U89860 ( .B1(n106945), .B2(n106860), .A(n99917), .ZN(
        \DLX_Datapath/ArithLogUnit/N126 ) );
  NAND2_X1 U89861 ( .A1(n99918), .A2(n105097), .ZN(n99917) );
  XNOR2_X1 U89862 ( .A(n99200), .B(n99919), .ZN(n99918) );
  XOR2_X1 U89863 ( .A(n99198), .B(n107426), .Z(n99919) );
  NAND2_X1 U89864 ( .A1(n99920), .A2(n99921), .ZN(n99199) );
  AOI22_X1 U89865 ( .A1(n107739), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[1] ), .B2(n99037), .ZN(n99921) );
  NAND2_X1 U89867 ( .A1(n99923), .A2(n99924), .ZN(n99383) );
  AOI22_X1 U89868 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] ), .A2(
        n99039), .B1(n107737), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .ZN(n99920) );
  AOI21_X1 U89869 ( .B1(n107553), .B2(n99925), .A(n99926), .ZN(n99198) );
  AOI21_X1 U89870 ( .B1(n99927), .B2(n107517), .A(n99928), .ZN(n99926) );
  XNOR2_X1 U89871 ( .A(n99929), .B(n99881), .ZN(n99200) );
  XNOR2_X1 U89872 ( .A(n99908), .B(n99930), .ZN(n99881) );
  XOR2_X1 U89873 ( .A(n99910), .B(n99907), .Z(n99930) );
  AOI22_X1 U89875 ( .A1(n99487), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] ), .B2(n99449), .ZN(n99932) );
  AOI22_X1 U89876 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] ), .B2(n99488), .ZN(n99931)
         );
  AOI21_X1 U89877 ( .B1(n99933), .B2(n107520), .A(n99934), .ZN(n99910) );
  AOI21_X1 U89878 ( .B1(n99935), .B2(n107541), .A(n99936), .ZN(n99934) );
  XOR2_X1 U89879 ( .A(n99937), .B(n99891), .Z(n99908) );
  NAND2_X1 U89881 ( .A1(n99939), .A2(n99940), .ZN(n99901) );
  AOI22_X1 U89882 ( .A1(n105105), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] ), .B2(n105106), .ZN(
        n99940) );
  AOI22_X1 U89883 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] ), .A2(
        n108741), .B1(n99719), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .ZN(n99939) );
  XOR2_X1 U89884 ( .A(n99904), .B(n99902), .Z(n99938) );
  NAND2_X1 U89885 ( .A1(n99941), .A2(n99942), .ZN(n99902) );
  AOI22_X1 U89886 ( .A1(n105108), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] ), .B2(n105109), .ZN(
        n99942) );
  AOI22_X1 U89887 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] ), .A2(
        n108742), .B1(n105107), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .ZN(n99941) );
  AOI21_X1 U89888 ( .B1(n105102), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] ), .A(n107561), .ZN(
        n99904) );
  AOI22_X1 U89889 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] ), .A2(
        n99764), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .ZN(n99943) );
  XOR2_X1 U89890 ( .A(n99890), .B(n107536), .Z(n99937) );
  NAND2_X1 U89891 ( .A1(n99944), .A2(n99945), .ZN(n99888) );
  AOI22_X1 U89892 ( .A1(n105111), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] ), .B2(n105112), .ZN(
        n99945) );
  AOI22_X1 U89893 ( .A1(n105110), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] ), .B2(n109085), .ZN(n99944) );
  OAI21_X1 U89894 ( .B1(n99946), .B2(n99947), .A(n99948), .ZN(n99890) );
  OAI21_X1 U89895 ( .B1(n107523), .B2(n107533), .A(n99949), .ZN(n99948) );
  XNOR2_X1 U89896 ( .A(n99880), .B(n99883), .ZN(n99929) );
  NAND2_X1 U89897 ( .A1(n99950), .A2(n99951), .ZN(n99883) );
  AOI22_X1 U89898 ( .A1(n105117), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] ), .B2(n99402), .ZN(n99951) );
  AOI22_X1 U89899 ( .A1(n105116), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] ), .B2(n108504), .ZN(n99950) );
  OAI21_X1 U89900 ( .B1(n99952), .B2(n99953), .A(n107512), .ZN(n99880) );
  AOI21_X1 U89901 ( .B1(n99953), .B2(n99952), .A(n99955), .ZN(n99954) );
  NAND2_X1 U89902 ( .A1(n99956), .A2(n99957), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [13]) );
  AOI22_X1 U89903 ( .A1(n105231), .A2(n69726), .B1(n105230), .B2(n111080), 
        .ZN(n99957) );
  AOI22_X1 U89904 ( .A1(n105229), .A2(DataAddr[13]), .B1(n105228), .B2(n108499), .ZN(n99956) );
  OAI21_X1 U89905 ( .B1(n106945), .B2(n106859), .A(n99958), .ZN(
        \DLX_Datapath/ArithLogUnit/N125 ) );
  NAND2_X1 U89906 ( .A1(n99959), .A2(n105097), .ZN(n99958) );
  XNOR2_X1 U89907 ( .A(n99207), .B(n99208), .ZN(n99959) );
  AOI21_X1 U89908 ( .B1(n105119), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[0] ), .A(n99960), .ZN(n99208)
         );
  NOR2_X1 U89909 ( .A1(n99382), .A2(n107568), .ZN(n99960) );
  NAND2_X1 U89910 ( .A1(n99923), .A2(n107738), .ZN(n99382) );
  NOR2_X1 U89911 ( .A1(n107738), .A2(n99923), .ZN(n99039) );
  NOR2_X1 U89912 ( .A1(n99922), .A2(\DLX_Datapath/ArithLogUnit/B_mul [13]), 
        .ZN(n99923) );
  NOR2_X1 U89913 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [12]), .A2(
        \DLX_Datapath/ArithLogUnit/B_mul [11]), .ZN(n99922) );
  OAI21_X1 U89914 ( .B1(n107740), .B2(n99961), .A(n99962), .ZN(n99924) );
  NAND2_X1 U89915 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [13]), .A2(n99963), 
        .ZN(n99962) );
  XOR2_X1 U89916 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [12]), .B(
        \DLX_Datapath/ArithLogUnit/B_mul [11]), .Z(n99963) );
  OR2_X1 U89917 ( .A1(n108505), .A2(\DLX_Datapath/ArithLogUnit/B_mul [13]), 
        .ZN(n99961) );
  XNOR2_X1 U89918 ( .A(n99964), .B(n99928), .ZN(n99207) );
  XNOR2_X1 U89919 ( .A(n99953), .B(n99965), .ZN(n99928) );
  XOR2_X1 U89920 ( .A(n99955), .B(n99952), .Z(n99965) );
  AOI22_X1 U89922 ( .A1(n105114), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] ), .B2(n99449), .ZN(n99967) );
  AOI22_X1 U89923 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] ), .B2(n105113), .ZN(n99966) );
  AOI21_X1 U89924 ( .B1(n99968), .B2(n107525), .A(n99969), .ZN(n99955) );
  AOI21_X1 U89925 ( .B1(n99970), .B2(n107544), .A(n99971), .ZN(n99969) );
  XOR2_X1 U89926 ( .A(n99972), .B(n99936), .Z(n99953) );
  NAND2_X1 U89928 ( .A1(n99974), .A2(n99975), .ZN(n99946) );
  AOI22_X1 U89929 ( .A1(n99718), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] ), .B2(n105106), .ZN(
        n99975) );
  AOI22_X1 U89930 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] ), .A2(
        n108741), .B1(n105104), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .ZN(n99974) );
  XOR2_X1 U89931 ( .A(n99949), .B(n99947), .Z(n99973) );
  NAND2_X1 U89932 ( .A1(n99976), .A2(n99977), .ZN(n99947) );
  AOI22_X1 U89933 ( .A1(n99623), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] ), .B2(n105109), .ZN(
        n99977) );
  AOI22_X1 U89934 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] ), .A2(
        n108742), .B1(n105107), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .ZN(n99976) );
  AOI21_X1 U89935 ( .B1(n105102), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] ), .A(n107562), .ZN(
        n99949) );
  AOI22_X1 U89936 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] ), .A2(
        n99764), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .ZN(n99978) );
  XOR2_X1 U89937 ( .A(n99935), .B(n107541), .Z(n99972) );
  NAND2_X1 U89938 ( .A1(n99979), .A2(n99980), .ZN(n99933) );
  AOI22_X1 U89939 ( .A1(n99541), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] ), .B2(n99515), .ZN(n99980) );
  AOI22_X1 U89940 ( .A1(n99540), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] ), .B2(n109085), .ZN(n99979) );
  OAI21_X1 U89941 ( .B1(n99981), .B2(n99982), .A(n99983), .ZN(n99935) );
  OAI21_X1 U89942 ( .B1(n107527), .B2(n107537), .A(n99984), .ZN(n99983) );
  XOR2_X1 U89943 ( .A(n107517), .B(n107553), .Z(n99964) );
  NAND2_X1 U89944 ( .A1(n99985), .A2(n99986), .ZN(n99927) );
  AOI22_X1 U89945 ( .A1(n99429), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] ), .B2(n99402), .ZN(n99986) );
  AOI22_X1 U89946 ( .A1(n105116), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] ), .B2(n108504), .ZN(n99985) );
  AOI21_X1 U89947 ( .B1(n99987), .B2(n107518), .A(n99988), .ZN(n99925) );
  AOI21_X1 U89948 ( .B1(n99989), .B2(n107550), .A(n99990), .ZN(n99988) );
  NAND2_X1 U89949 ( .A1(n99991), .A2(n99992), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [12]) );
  AOI22_X1 U89950 ( .A1(n105231), .A2(n69727), .B1(n105230), .B2(n111097), 
        .ZN(n99992) );
  AOI22_X1 U89951 ( .A1(n105229), .A2(DataAddr[12]), .B1(n105228), .B2(n107736), .ZN(n99991) );
  OAI21_X1 U89952 ( .B1(n106945), .B2(n106858), .A(n99993), .ZN(
        \DLX_Datapath/ArithLogUnit/N124 ) );
  NAND2_X1 U89953 ( .A1(n99994), .A2(n105097), .ZN(n99993) );
  XNOR2_X1 U89954 ( .A(n99995), .B(n99215), .ZN(n99994) );
  XOR2_X1 U89955 ( .A(n99989), .B(n99996), .Z(n99215) );
  XOR2_X1 U89956 ( .A(n99990), .B(n107550), .Z(n99996) );
  NAND2_X1 U89957 ( .A1(n99997), .A2(n99998), .ZN(n99987) );
  AOI22_X1 U89958 ( .A1(n105114), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] ), .B2(n99449), .ZN(n99998) );
  AOI22_X1 U89959 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] ), .B2(n105113), .ZN(n99997) );
  AOI21_X1 U89960 ( .B1(n99999), .B2(n107529), .A(n100000), .ZN(n99990) );
  AOI21_X1 U89961 ( .B1(n100001), .B2(n107546), .A(n100002), .ZN(n100000) );
  XOR2_X1 U89962 ( .A(n100003), .B(n99971), .Z(n99989) );
  NAND2_X1 U89964 ( .A1(n100005), .A2(n100006), .ZN(n99981) );
  AOI22_X1 U89965 ( .A1(n105105), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] ), .B2(n105106), .ZN(
        n100006) );
  AOI22_X1 U89966 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] ), .A2(
        n108741), .B1(n99719), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .ZN(n100005) );
  XOR2_X1 U89967 ( .A(n99984), .B(n99982), .Z(n100004) );
  NAND2_X1 U89968 ( .A1(n100007), .A2(n100008), .ZN(n99982) );
  AOI22_X1 U89969 ( .A1(n105108), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] ), .B2(n105109), .ZN(
        n100008) );
  AOI22_X1 U89970 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] ), .A2(
        n108742), .B1(n99624), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .ZN(n100007) );
  AOI21_X1 U89971 ( .B1(n105102), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] ), .A(n107563), .ZN(
        n99984) );
  AOI22_X1 U89972 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] ), .A2(
        n99764), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .ZN(n100009) );
  XOR2_X1 U89973 ( .A(n99970), .B(n107544), .Z(n100003) );
  NAND2_X1 U89974 ( .A1(n100010), .A2(n100011), .ZN(n99968) );
  AOI22_X1 U89975 ( .A1(n105111), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] ), .B2(n99515), .ZN(
        n100011) );
  AOI22_X1 U89976 ( .A1(n105110), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] ), .B2(n109085), .ZN(
        n100010) );
  OAI21_X1 U89977 ( .B1(n100012), .B2(n100013), .A(n100014), .ZN(n99970) );
  OAI21_X1 U89978 ( .B1(n107534), .B2(n107542), .A(n100015), .ZN(n100014) );
  NAND2_X1 U89980 ( .A1(n100016), .A2(n100017), .ZN(n99217) );
  AOI22_X1 U89981 ( .A1(n105117), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[1] ), .B2(n99402), .ZN(
        n100017) );
  NOR2_X1 U89982 ( .A1(n100018), .A2(n108505), .ZN(n99402) );
  NOR2_X1 U89983 ( .A1(n100019), .A2(n108503), .ZN(n99429) );
  AOI22_X1 U89984 ( .A1(n99428), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] ), .B2(n108504), .ZN(
        n100016) );
  AOI21_X1 U89985 ( .B1(n100021), .B2(n100022), .A(n107524), .ZN(n99218) );
  OAI21_X1 U89986 ( .B1(n100022), .B2(n100021), .A(n100024), .ZN(n100023) );
  NAND2_X1 U89987 ( .A1(n100025), .A2(n100026), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [11]) );
  AOI22_X1 U89988 ( .A1(n98953), .A2(n69728), .B1(n98954), .B2(n111081), .ZN(
        n100026) );
  AOI22_X1 U89989 ( .A1(n98955), .A2(DataAddr[11]), .B1(n98956), .B2(n109651), 
        .ZN(n100025) );
  OAI21_X1 U89990 ( .B1(n106945), .B2(n106857), .A(n100027), .ZN(
        \DLX_Datapath/ArithLogUnit/N123 ) );
  NAND2_X1 U89991 ( .A1(n100028), .A2(n105098), .ZN(n100027) );
  XNOR2_X1 U89992 ( .A(n99225), .B(n99226), .ZN(n100028) );
  AOI21_X1 U89993 ( .B1(n108504), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[0] ), .A(n100029), .ZN(n99226)
         );
  NOR2_X1 U89995 ( .A1(n100019), .A2(n100020), .ZN(n99428) );
  NAND2_X1 U89996 ( .A1(n100020), .A2(n100019), .ZN(n99404) );
  NAND2_X1 U89997 ( .A1(n100018), .A2(n108505), .ZN(n100019) );
  OR2_X1 U89998 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [9]), .A2(
        \DLX_Datapath/ArithLogUnit/B_mul [10]), .ZN(n100018) );
  OAI21_X1 U89999 ( .B1(n108505), .B2(n100030), .A(n100031), .ZN(n100020) );
  NAND2_X1 U90000 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [9]), .A2(n100032), 
        .ZN(n100031) );
  XOR2_X1 U90001 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [11]), .B(
        \DLX_Datapath/ArithLogUnit/B_mul [10]), .Z(n100032) );
  NAND2_X1 U90002 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [10]), .A2(n109762), 
        .ZN(n100030) );
  XOR2_X1 U90003 ( .A(n100033), .B(n100021), .Z(n99225) );
  XOR2_X1 U90004 ( .A(n100034), .B(n100002), .Z(n100021) );
  NAND2_X1 U90006 ( .A1(n100036), .A2(n100037), .ZN(n100012) );
  AOI22_X1 U90007 ( .A1(n99718), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] ), .B2(n105106), .ZN(
        n100037) );
  AOI22_X1 U90008 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] ), .A2(
        n108741), .B1(n105104), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .ZN(n100036) );
  XOR2_X1 U90009 ( .A(n100015), .B(n100013), .Z(n100035) );
  NAND2_X1 U90010 ( .A1(n100038), .A2(n100039), .ZN(n100013) );
  AOI22_X1 U90011 ( .A1(n99623), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] ), .B2(n105109), .ZN(
        n100039) );
  AOI22_X1 U90012 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] ), .A2(
        n108742), .B1(n99624), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .ZN(n100038) );
  AOI21_X1 U90013 ( .B1(n105102), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] ), .A(n107564), .ZN(
        n100015) );
  AOI22_X1 U90014 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] ), .A2(
        n99764), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .ZN(n100040) );
  XOR2_X1 U90015 ( .A(n100001), .B(n107546), .Z(n100034) );
  NAND2_X1 U90016 ( .A1(n100041), .A2(n100042), .ZN(n99999) );
  AOI22_X1 U90017 ( .A1(n99541), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] ), .B2(n99515), .ZN(
        n100042) );
  AOI22_X1 U90018 ( .A1(n105110), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] ), .B2(n109085), .ZN(
        n100041) );
  OAI21_X1 U90019 ( .B1(n100043), .B2(n100044), .A(n107530), .ZN(n100001) );
  AOI21_X1 U90020 ( .B1(n100043), .B2(n100044), .A(n100046), .ZN(n100045) );
  XNOR2_X1 U90021 ( .A(n100024), .B(n100022), .ZN(n100033) );
  AOI22_X1 U90023 ( .A1(n99487), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] ), .B2(n99449), .ZN(
        n100048) );
  AOI22_X1 U90024 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] ), .B2(n105113), .ZN(
        n100047) );
  AOI21_X1 U90025 ( .B1(n100049), .B2(n100050), .A(n107528), .ZN(n100024) );
  OAI21_X1 U90026 ( .B1(n100050), .B2(n100049), .A(n100052), .ZN(n100051) );
  NAND2_X1 U90027 ( .A1(n100053), .A2(n100054), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [10]) );
  AOI22_X1 U90028 ( .A1(n98953), .A2(n69729), .B1(n98954), .B2(n111082), .ZN(
        n100054) );
  AOI22_X1 U90029 ( .A1(n98955), .A2(DataAddr[10]), .B1(n98956), .B2(n108613), 
        .ZN(n100053) );
  OAI21_X1 U90030 ( .B1(n106945), .B2(n106856), .A(n100055), .ZN(
        \DLX_Datapath/ArithLogUnit/N122 ) );
  NAND2_X1 U90031 ( .A1(n100056), .A2(n105097), .ZN(n100055) );
  XNOR2_X1 U90032 ( .A(n99234), .B(n100057), .ZN(n100056) );
  XOR2_X1 U90033 ( .A(n99236), .B(n99233), .Z(n100057) );
  AOI22_X1 U90035 ( .A1(n105114), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[1] ), .B2(n99449), .ZN(
        n100059) );
  NOR2_X1 U90036 ( .A1(n100060), .A2(n109762), .ZN(n99449) );
  OR2_X1 U90037 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [8]), .A2(
        \DLX_Datapath/ArithLogUnit/B_mul [7]), .ZN(n100060) );
  NOR2_X1 U90038 ( .A1(n100061), .A2(n100062), .ZN(n99487) );
  AOI22_X1 U90039 ( .A1(n109088), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] ), .B2(n99488), .ZN(n100058) );
  AOI21_X1 U90040 ( .B1(n100064), .B2(n107538), .A(n100065), .ZN(n99236) );
  AOI21_X1 U90041 ( .B1(n100066), .B2(n107554), .A(n100067), .ZN(n100065) );
  XNOR2_X1 U90042 ( .A(n100068), .B(n100050), .ZN(n99234) );
  XNOR2_X1 U90043 ( .A(n100069), .B(n100043), .ZN(n100050) );
  NAND2_X1 U90044 ( .A1(n100070), .A2(n100071), .ZN(n100043) );
  AOI22_X1 U90045 ( .A1(n105108), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] ), .B2(n105109), .ZN(
        n100071) );
  AOI22_X1 U90046 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] ), .A2(
        n108742), .B1(n99624), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .ZN(n100070) );
  XNOR2_X1 U90047 ( .A(n100046), .B(n100044), .ZN(n100069) );
  NAND2_X1 U90048 ( .A1(n100072), .A2(n100073), .ZN(n100044) );
  AOI22_X1 U90049 ( .A1(n105105), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] ), .B2(n105106), .ZN(
        n100073) );
  AOI22_X1 U90050 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] ), .A2(
        n108741), .B1(n105104), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .ZN(n100072) );
  OAI21_X1 U90051 ( .B1(n109759), .B2(n99851), .A(n100074), .ZN(n100046) );
  AOI22_X1 U90052 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] ), .A2(
        n105103), .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] ), .B2(
        n105102), .ZN(n100074) );
  XOR2_X1 U90053 ( .A(n100052), .B(n100049), .Z(n100068) );
  NAND2_X1 U90054 ( .A1(n100075), .A2(n100076), .ZN(n100049) );
  AOI22_X1 U90055 ( .A1(n105111), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] ), .B2(n99515), .ZN(
        n100076) );
  AOI22_X1 U90056 ( .A1(n99540), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] ), .B2(n109085), .ZN(
        n100075) );
  AOI21_X1 U90057 ( .B1(n107543), .B2(n107547), .A(n100077), .ZN(n100052) );
  AOI21_X1 U90058 ( .B1(n100078), .B2(n100079), .A(n100080), .ZN(n100077) );
  NAND2_X1 U90059 ( .A1(n100081), .A2(n100082), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [9]) );
  AOI22_X1 U90060 ( .A1(n98953), .A2(n69706), .B1(n98954), .B2(n111075), .ZN(
        n100082) );
  AOI22_X1 U90061 ( .A1(n98955), .A2(DataAddr[9]), .B1(n98956), .B2(n109758), 
        .ZN(n100081) );
  OAI21_X1 U90062 ( .B1(n106945), .B2(n106855), .A(n100083), .ZN(
        \DLX_Datapath/ArithLogUnit/N121 ) );
  NAND2_X1 U90063 ( .A1(n100084), .A2(n105097), .ZN(n100083) );
  XNOR2_X1 U90064 ( .A(n99243), .B(n99244), .ZN(n100084) );
  AOI21_X1 U90065 ( .B1(n99488), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[0] ), .A(n100085), .ZN(n99244)
         );
  NOR2_X1 U90066 ( .A1(n100063), .A2(n107568), .ZN(n100085) );
  NAND2_X1 U90067 ( .A1(n109090), .A2(n100062), .ZN(n100063) );
  NOR2_X1 U90068 ( .A1(n109090), .A2(n100062), .ZN(n99488) );
  NOR2_X1 U90072 ( .A1(n109089), .A2(\DLX_Datapath/ArithLogUnit/B_mul [9]), 
        .ZN(n100086) );
  OAI21_X1 U90073 ( .B1(\DLX_Datapath/ArithLogUnit/B_mul [8]), .B2(
        \DLX_Datapath/ArithLogUnit/B_mul [7]), .A(n109762), .ZN(n100061) );
  XNOR2_X1 U90074 ( .A(n100089), .B(n100067), .ZN(n99243) );
  NAND2_X1 U90076 ( .A1(n100091), .A2(n100092), .ZN(n100078) );
  AOI22_X1 U90077 ( .A1(n99718), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] ), .B2(n99667), .ZN(
        n100092) );
  AOI22_X1 U90078 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] ), .A2(
        n108741), .B1(n105104), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .ZN(n100091) );
  XOR2_X1 U90079 ( .A(n100080), .B(n107547), .Z(n100090) );
  NAND2_X1 U90080 ( .A1(n100093), .A2(n100094), .ZN(n100079) );
  AOI22_X1 U90081 ( .A1(n99623), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] ), .B2(n105109), .ZN(
        n100094) );
  AOI22_X1 U90082 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] ), .A2(
        n108742), .B1(n99624), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .ZN(n100093) );
  OAI21_X1 U90083 ( .B1(n107570), .B2(n107531), .A(n100095), .ZN(n100080) );
  AOI22_X1 U90084 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] ), .A2(
        n105103), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .ZN(n100095) );
  XOR2_X1 U90085 ( .A(n100066), .B(n107554), .Z(n100089) );
  NAND2_X1 U90086 ( .A1(n100096), .A2(n100097), .ZN(n100064) );
  AOI22_X1 U90087 ( .A1(n99541), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] ), .B2(n99515), .ZN(
        n100097) );
  AOI22_X1 U90088 ( .A1(n99540), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] ), .B2(n109085), .ZN(
        n100096) );
  OAI21_X1 U90089 ( .B1(n100098), .B2(n100099), .A(n107539), .ZN(n100066) );
  AOI21_X1 U90090 ( .B1(n100098), .B2(n100099), .A(n100101), .ZN(n100100) );
  NAND2_X1 U90091 ( .A1(n100102), .A2(n100103), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [8]) );
  AOI22_X1 U90092 ( .A1(n105231), .A2(n69707), .B1(n98954), .B2(n111076), .ZN(
        n100103) );
  AOI22_X1 U90093 ( .A1(n98955), .A2(DataAddr[8]), .B1(n98956), .B2(n109543), 
        .ZN(n100102) );
  OAI21_X1 U90094 ( .B1(n106945), .B2(n106854), .A(n100104), .ZN(
        \DLX_Datapath/ArithLogUnit/N120 ) );
  NAND2_X1 U90095 ( .A1(n100105), .A2(n105096), .ZN(n100104) );
  XOR2_X1 U90096 ( .A(n99254), .B(n100106), .Z(n100105) );
  XNOR2_X1 U90097 ( .A(n99252), .B(n99251), .ZN(n100106) );
  AOI22_X1 U90099 ( .A1(n105111), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[1] ), .B2(n99515), .ZN(
        n100108) );
  NOR2_X1 U90100 ( .A1(n100109), .A2(n109089), .ZN(n99515) );
  NAND2_X1 U90101 ( .A1(n109432), .A2(n109310), .ZN(n100109) );
  NOR2_X1 U90102 ( .A1(n100110), .A2(n109086), .ZN(n99541) );
  AOI22_X1 U90103 ( .A1(n105110), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] ), .B2(n109085), .ZN(
        n100107) );
  OAI21_X1 U90104 ( .B1(n100112), .B2(n100113), .A(n100114), .ZN(n99252) );
  OAI21_X1 U90105 ( .B1(n107548), .B2(n107555), .A(n100115), .ZN(n100114) );
  XOR2_X1 U90106 ( .A(n100116), .B(n100098), .Z(n99254) );
  NAND2_X1 U90107 ( .A1(n100117), .A2(n100118), .ZN(n100098) );
  AOI22_X1 U90108 ( .A1(n105108), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] ), .B2(n99625), .ZN(
        n100118) );
  AOI22_X1 U90109 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] ), .A2(
        n108742), .B1(n99624), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .ZN(n100117) );
  XNOR2_X1 U90110 ( .A(n100101), .B(n100099), .ZN(n100116) );
  NAND2_X1 U90111 ( .A1(n100119), .A2(n100120), .ZN(n100099) );
  AOI22_X1 U90112 ( .A1(n105105), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] ), .B2(n99667), .ZN(
        n100120) );
  AOI22_X1 U90113 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] ), .A2(
        n108741), .B1(n99719), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .ZN(n100119) );
  OAI21_X1 U90114 ( .B1(n109082), .B2(n99851), .A(n100121), .ZN(n100101) );
  AOI22_X1 U90115 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] ), .A2(
        n105103), .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] ), .B2(
        n105102), .ZN(n100121) );
  NAND2_X1 U90116 ( .A1(n100122), .A2(n100123), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [7]) );
  AOI22_X1 U90117 ( .A1(n105231), .A2(n69730), .B1(n105230), .B2(n111088), 
        .ZN(n100123) );
  AOI22_X1 U90118 ( .A1(n98955), .A2(DataAddr[7]), .B1(n105228), .B2(n109081), 
        .ZN(n100122) );
  OAI21_X1 U90119 ( .B1(n106945), .B2(n106853), .A(n100124), .ZN(
        \DLX_Datapath/ArithLogUnit/N119 ) );
  NAND2_X1 U90120 ( .A1(n100125), .A2(n105097), .ZN(n100124) );
  XNOR2_X1 U90121 ( .A(n99262), .B(n99261), .ZN(n100125) );
  XOR2_X1 U90122 ( .A(n100126), .B(n107548), .Z(n99261) );
  NAND2_X1 U90123 ( .A1(n100127), .A2(n100128), .ZN(n100112) );
  AOI22_X1 U90124 ( .A1(n99718), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] ), .B2(n99667), .ZN(
        n100128) );
  AOI22_X1 U90125 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] ), .A2(
        n108741), .B1(n99719), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .ZN(n100127) );
  XOR2_X1 U90126 ( .A(n100115), .B(n100113), .Z(n100126) );
  NAND2_X1 U90127 ( .A1(n100129), .A2(n100130), .ZN(n100113) );
  AOI22_X1 U90128 ( .A1(n99623), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] ), .B2(n99625), .ZN(
        n100130) );
  AOI22_X1 U90129 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] ), .A2(
        n108742), .B1(n99624), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .ZN(n100129) );
  AOI21_X1 U90130 ( .B1(n105102), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] ), .A(n107565), .ZN(
        n100115) );
  AOI22_X1 U90131 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] ), .A2(
        n105103), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .ZN(n100131) );
  AOI21_X1 U90132 ( .B1(n109085), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[0] ), .A(n100132), .ZN(n99262)
         );
  NOR2_X1 U90134 ( .A1(n100110), .A2(n100111), .ZN(n99540) );
  NAND2_X1 U90135 ( .A1(n100110), .A2(n100111), .ZN(n99517) );
  OAI21_X1 U90136 ( .B1(n109432), .B2(n100133), .A(n100134), .ZN(n100111) );
  NAND2_X1 U90137 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [7]), .A2(n100135), 
        .ZN(n100134) );
  XOR2_X1 U90138 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [6]), .B(
        \DLX_Datapath/ArithLogUnit/B_mul [5]), .Z(n100135) );
  NAND2_X1 U90139 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [5]), .A2(n109089), 
        .ZN(n100133) );
  OAI21_X1 U90140 ( .B1(\DLX_Datapath/ArithLogUnit/B_mul [6]), .B2(
        \DLX_Datapath/ArithLogUnit/B_mul [5]), .A(n109089), .ZN(n100110) );
  NAND2_X1 U90141 ( .A1(n100136), .A2(n100137), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [6]) );
  AOI22_X1 U90142 ( .A1(n105231), .A2(n69699), .B1(n105230), .B2(n111083), 
        .ZN(n100137) );
  AOI22_X1 U90143 ( .A1(n98955), .A2(DataAddr[6]), .B1(n105228), .B2(n109428), 
        .ZN(n100136) );
  OAI21_X1 U90144 ( .B1(n106945), .B2(n106852), .A(n100138), .ZN(
        \DLX_Datapath/ArithLogUnit/N118 ) );
  NAND2_X1 U90145 ( .A1(n100139), .A2(n105098), .ZN(n100138) );
  XNOR2_X1 U90146 ( .A(n100140), .B(n99270), .ZN(n100139) );
  NAND2_X1 U90147 ( .A1(n100141), .A2(n100142), .ZN(n99270) );
  AOI22_X1 U90148 ( .A1(n105108), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[1] ), .B2(n99625), .ZN(
        n100142) );
  NOR2_X1 U90151 ( .A1(n100144), .A2(n100145), .ZN(n99623) );
  AOI22_X1 U90152 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] ), .A2(
        n108742), .B1(n99624), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .ZN(n100141) );
  XNOR2_X1 U90153 ( .A(n99272), .B(n99271), .ZN(n100140) );
  NAND2_X1 U90154 ( .A1(n100147), .A2(n100148), .ZN(n99271) );
  AOI22_X1 U90155 ( .A1(n105105), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] ), .B2(n99667), .ZN(
        n100148) );
  AOI22_X1 U90156 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] ), .A2(
        n108741), .B1(n105104), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .ZN(n100147) );
  OAI21_X1 U90157 ( .B1(n109313), .B2(n99851), .A(n100149), .ZN(n99272) );
  AOI22_X1 U90158 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] ), .A2(
        n105103), .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] ), .B2(
        n105102), .ZN(n100149) );
  NAND2_X1 U90159 ( .A1(n100150), .A2(n100151), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [5]) );
  AOI22_X1 U90160 ( .A1(n105231), .A2(n69700), .B1(n105230), .B2(n111077), 
        .ZN(n100151) );
  AOI22_X1 U90161 ( .A1(n98955), .A2(DataAddr[5]), .B1(n105228), .B2(n109309), 
        .ZN(n100150) );
  XNOR2_X1 U90164 ( .A(n99280), .B(n100154), .ZN(n100153) );
  XOR2_X1 U90165 ( .A(n99282), .B(n99279), .Z(n100154) );
  NAND2_X1 U90168 ( .A1(n108743), .A2(n100145), .ZN(n100146) );
  NOR2_X1 U90169 ( .A1(n100145), .A2(n108743), .ZN(n99624) );
  OAI21_X1 U90170 ( .B1(n109310), .B2(n100156), .A(n100157), .ZN(n100144) );
  OAI21_X1 U90171 ( .B1(n108745), .B2(n109202), .A(n109310), .ZN(n100157) );
  XOR2_X1 U90172 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [4]), .B(
        \DLX_Datapath/ArithLogUnit/B_mul [3]), .Z(n100156) );
  OAI21_X1 U90173 ( .B1(\DLX_Datapath/ArithLogUnit/B_mul [4]), .B2(
        \DLX_Datapath/ArithLogUnit/B_mul [3]), .A(n109310), .ZN(n100145) );
  AOI21_X1 U90174 ( .B1(n99849), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] ), .A(n107566), .ZN(n99282) );
  AOI22_X1 U90175 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] ), .A2(
        n105103), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .ZN(n100158) );
  AOI22_X1 U90177 ( .A1(n99718), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] ), .B2(n99667), .ZN(
        n100160) );
  AOI22_X1 U90178 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] ), .A2(
        n108741), .B1(n99719), .B2(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .ZN(n100159) );
  NAND2_X1 U90179 ( .A1(n100161), .A2(n100162), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [4]) );
  AOI22_X1 U90180 ( .A1(n105231), .A2(n69701), .B1(n105230), .B2(n111089), 
        .ZN(n100162) );
  AOI22_X1 U90181 ( .A1(n105229), .A2(DataAddr[4]), .B1(n105228), .B2(n109201), 
        .ZN(n100161) );
  OAI21_X1 U90182 ( .B1(n105196), .B2(n106851), .A(n100163), .ZN(
        \DLX_Datapath/ArithLogUnit/N116 ) );
  NAND2_X1 U90183 ( .A1(n100164), .A2(n105096), .ZN(n100163) );
  XOR2_X1 U90184 ( .A(n99290), .B(n99289), .Z(n100164) );
  OAI21_X1 U90185 ( .B1(n108737), .B2(n99851), .A(n100165), .ZN(n99289) );
  AOI22_X1 U90186 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] ), .A2(
        n105103), .B1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] ), .B2(
        n105102), .ZN(n100165) );
  NAND2_X1 U90187 ( .A1(n100166), .A2(n100167), .ZN(n99290) );
  AOI22_X1 U90188 ( .A1(n105105), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .B1(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[1] ), .B2(n99667), .ZN(
        n100167) );
  NOR2_X1 U90189 ( .A1(n100168), .A2(n108745), .ZN(n99667) );
  NAND2_X1 U90190 ( .A1(n108968), .A2(n108857), .ZN(n100168) );
  NOR2_X1 U90191 ( .A1(n100169), .A2(n108740), .ZN(n99718) );
  AOI22_X1 U90192 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] ), .A2(
        n108741), .B1(n105104), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .ZN(n100166) );
  NAND2_X1 U90193 ( .A1(n100171), .A2(n100172), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [3]) );
  AOI22_X1 U90194 ( .A1(n105231), .A2(n69702), .B1(n105230), .B2(n111084), 
        .ZN(n100172) );
  AOI22_X1 U90195 ( .A1(n98955), .A2(DataAddr[3]), .B1(n105228), .B2(n108736), 
        .ZN(n100171) );
  OAI21_X1 U90196 ( .B1(n106945), .B2(n106850), .A(n100173), .ZN(
        \DLX_Datapath/ArithLogUnit/N115 ) );
  NAND2_X1 U90197 ( .A1(n100174), .A2(n105098), .ZN(n100173) );
  XNOR2_X1 U90198 ( .A(n99298), .B(n99297), .ZN(n100174) );
  OAI21_X1 U90199 ( .B1(n99665), .B2(n107568), .A(n100175), .ZN(n99297) );
  NAND2_X1 U90200 ( .A1(n99719), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .ZN(n100175) );
  NOR2_X1 U90201 ( .A1(n100170), .A2(n100169), .ZN(n99719) );
  NAND2_X1 U90202 ( .A1(n100170), .A2(n100169), .ZN(n99665) );
  OAI21_X1 U90203 ( .B1(\DLX_Datapath/ArithLogUnit/B_mul [2]), .B2(
        \DLX_Datapath/ArithLogUnit/B_mul [1]), .A(n108745), .ZN(n100169) );
  OAI21_X1 U90204 ( .B1(n108968), .B2(n100176), .A(n100177), .ZN(n100170) );
  NAND2_X1 U90205 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [3]), .A2(n100178), 
        .ZN(n100177) );
  XOR2_X1 U90206 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [2]), .B(
        \DLX_Datapath/ArithLogUnit/B_mul [1]), .Z(n100178) );
  NAND2_X1 U90207 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [1]), .A2(n108745), 
        .ZN(n100176) );
  AOI21_X1 U90208 ( .B1(n99849), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] ), .A(n107567), .ZN(n99298) );
  AOI22_X1 U90209 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] ), .A2(
        n105103), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .ZN(n100179) );
  NAND2_X1 U90210 ( .A1(n100180), .A2(n100181), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [2]) );
  AOI22_X1 U90211 ( .A1(n105231), .A2(n69703), .B1(n105230), .B2(n111085), 
        .ZN(n100181) );
  AOI22_X1 U90212 ( .A1(n105229), .A2(DataAddr[2]), .B1(n105228), .B2(n108964), 
        .ZN(n100180) );
  OAI21_X1 U90213 ( .B1(n105196), .B2(n106849), .A(n100182), .ZN(
        \DLX_Datapath/ArithLogUnit/N114 ) );
  NAND2_X1 U90214 ( .A1(n100183), .A2(n105098), .ZN(n100182) );
  OAI21_X1 U90215 ( .B1(n108855), .B2(n99851), .A(n100184), .ZN(n100183) );
  AOI22_X1 U90216 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] ), .A2(
        n105103), .B1(n105102), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .ZN(n100184) );
  NAND2_X1 U90217 ( .A1(n100185), .A2(n100186), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [1]) );
  AOI22_X1 U90218 ( .A1(n105231), .A2(n69704), .B1(n105230), .B2(n111086), 
        .ZN(n100186) );
  AOI22_X1 U90219 ( .A1(n98955), .A2(DataAddr[1]), .B1(n105228), .B2(n108853), 
        .ZN(n100185) );
  OAI21_X1 U90220 ( .B1(n105899), .B2(n100187), .A(n100188), .ZN(
        \DLX_Datapath/ArithLogUnit/N113 ) );
  NAND2_X1 U90221 ( .A1(\DLX_Datapath/MUX_HDU_ALUInA [0]), .A2(n81805), .ZN(
        n100188) );
  NAND2_X1 U90222 ( .A1(n100189), .A2(n100190), .ZN(
        \DLX_Datapath/MUX_HDU_ALUInA [0]) );
  AOI22_X1 U90223 ( .A1(n105231), .A2(n69705), .B1(n105230), .B2(n111087), 
        .ZN(n100190) );
  NOR2_X1 U90224 ( .A1(n100191), .A2(n100192), .ZN(n98954) );
  NOR2_X1 U90225 ( .A1(n106878), .A2(n100191), .ZN(n98953) );
  AOI22_X1 U90226 ( .A1(n105229), .A2(DataAddr[0]), .B1(n105228), .B2(n107419), 
        .ZN(n100189) );
  NOR2_X1 U90227 ( .A1(n106879), .A2(n100192), .ZN(n98956) );
  NOR2_X1 U90228 ( .A1(n106878), .A2(n106879), .ZN(n98955) );
  NAND2_X1 U90229 ( .A1(n100193), .A2(n100194), .ZN(n100191) );
  NOR2_X1 U90230 ( .A1(n100195), .A2(n100196), .ZN(n100193) );
  AOI22_X1 U90231 ( .A1(n100197), .A2(n100198), .B1(n100199), .B2(n99350), 
        .ZN(n100196) );
  OR2_X1 U90232 ( .A1(n83105), .A2(n99323), .ZN(n99350) );
  OAI21_X1 U90233 ( .B1(n100200), .B2(n100201), .A(n100202), .ZN(n83105) );
  NAND2_X1 U90234 ( .A1(n69380), .A2(n100203), .ZN(n100202) );
  OAI21_X1 U90235 ( .B1(n69382), .B2(n100204), .A(n100205), .ZN(n100203) );
  AOI22_X1 U90236 ( .A1(n100206), .A2(n69319), .B1(n100204), .B2(n111055), 
        .ZN(n100205) );
  NOR2_X1 U90237 ( .A1(n69324), .A2(n111055), .ZN(n100206) );
  NAND2_X1 U90239 ( .A1(n69324), .A2(n69319), .ZN(n100201) );
  OAI21_X1 U90240 ( .B1(n69378), .B2(n100762), .A(n100207), .ZN(n100200) );
  NOR2_X1 U90241 ( .A1(n69382), .A2(n69380), .ZN(n100207) );
  NOR4_X1 U90242 ( .A1(n86273), .A2(n100208), .A3(n100209), .A4(n100210), .ZN(
        n100198) );
  XOR2_X1 U90243 ( .A(n100429), .B(n54618), .Z(n100210) );
  XOR2_X1 U90244 ( .A(n100430), .B(n54616), .Z(n100209) );
  XOR2_X1 U90245 ( .A(n100428), .B(n54614), .Z(n100208) );
  NAND2_X1 U90246 ( .A1(n100211), .A2(n100212), .ZN(n86273) );
  NOR3_X1 U90247 ( .A1(n69378), .A2(n69382), .A3(n69380), .ZN(n100212) );
  NOR3_X1 U90248 ( .A1(n106944), .A2(n69324), .A3(n69319), .ZN(n100211) );
  NOR4_X1 U90249 ( .A1(n100213), .A2(n100214), .A3(n100215), .A4(n100216), 
        .ZN(n100197) );
  XOR2_X1 U90250 ( .A(n100217), .B(n86282), .Z(n100216) );
  OAI21_X1 U90251 ( .B1(n104497), .B2(n107129), .A(n100218), .ZN(n86282) );
  XOR2_X1 U90252 ( .A(n100219), .B(n107107), .Z(n100218) );
  XNOR2_X1 U90253 ( .A(n86283), .B(n100220), .ZN(n100215) );
  NOR2_X1 U90254 ( .A1(n100219), .A2(n100221), .ZN(n86283) );
  AOI21_X1 U90255 ( .B1(n107105), .B2(n107129), .A(n104497), .ZN(n100221) );
  XOR2_X1 U90256 ( .A(n86285), .B(n100222), .Z(n100214) );
  OAI21_X1 U90257 ( .B1(n104497), .B2(n107129), .A(n100223), .ZN(n86285) );
  XOR2_X1 U90258 ( .A(n107109), .B(n100224), .Z(n100223) );
  NAND2_X1 U90259 ( .A1(n100219), .A2(n107107), .ZN(n100224) );
  NOR2_X1 U90260 ( .A1(n58722), .A2(n54623), .ZN(n100219) );
  XOR2_X1 U90261 ( .A(n100893), .B(n100894), .Z(n100213) );
  AOI21_X1 U90262 ( .B1(n100225), .B2(n100194), .A(n100195), .ZN(n100192) );
  NOR3_X1 U90265 ( .A1(n106880), .A2(n69326), .A3(n100230), .ZN(n100229) );
  AOI21_X1 U90266 ( .B1(n59415), .B2(n106937), .A(n59419), .ZN(n100230) );
  AOI22_X1 U90268 ( .A1(n100234), .A2(n100235), .B1(n100236), .B2(n100237), 
        .ZN(n100194) );
  NOR4_X1 U90269 ( .A1(n82682), .A2(n100238), .A3(n100239), .A4(n100240), .ZN(
        n100237) );
  XOR2_X1 U90270 ( .A(n100419), .B(n100429), .Z(n100240) );
  XOR2_X1 U90271 ( .A(n100418), .B(n100428), .Z(n100239) );
  XOR2_X1 U90272 ( .A(n100420), .B(n100430), .Z(n100238) );
  NAND2_X1 U90273 ( .A1(n100241), .A2(n100242), .ZN(n82682) );
  NOR3_X1 U90274 ( .A1(\DLX_Datapath/IR_EXMEM[29] ), .A2(n69323), .A3(
        \DLX_Datapath/IR_EXMEM[27] ), .ZN(n100242) );
  NOR3_X1 U90275 ( .A1(n111022), .A2(\DLX_Datapath/IR_EXMEM[31] ), .A3(n106943), .ZN(n100241) );
  NOR4_X1 U90276 ( .A1(n100243), .A2(n100244), .A3(n100245), .A4(n100246), 
        .ZN(n100236) );
  XOR2_X1 U90277 ( .A(n100217), .B(n82689), .Z(n100246) );
  NAND2_X1 U90278 ( .A1(n100247), .A2(n100248), .ZN(n82689) );
  XOR2_X1 U90279 ( .A(n104950), .B(n100249), .Z(n100247) );
  XOR2_X1 U90280 ( .A(n82686), .B(n100220), .Z(n100245) );
  NAND2_X1 U90281 ( .A1(n100249), .A2(n100250), .ZN(n82686) );
  XOR2_X1 U90283 ( .A(n104722), .B(n100222), .Z(n100244) );
  NAND2_X1 U90284 ( .A1(n100251), .A2(n100248), .ZN(n99340) );
  NAND2_X1 U90285 ( .A1(n62661), .A2(n62662), .ZN(n100248) );
  NOR2_X1 U90287 ( .A1(n104950), .A2(n100249), .ZN(n100252) );
  OR2_X1 U90288 ( .A1(n107104), .A2(n62661), .ZN(n100249) );
  XOR2_X1 U90289 ( .A(n100893), .B(n62662), .Z(n100243) );
  NOR4_X1 U90290 ( .A1(n106939), .A2(n100253), .A3(n100254), .A4(n100255), 
        .ZN(n100235) );
  XOR2_X1 U90291 ( .A(n100422), .B(n100429), .Z(n100255) );
  XOR2_X1 U90292 ( .A(n100423), .B(n100430), .Z(n100254) );
  XOR2_X1 U90293 ( .A(n100428), .B(n100796), .Z(n100253) );
  OAI21_X1 U90294 ( .B1(n59325), .B2(n100257), .A(n100258), .ZN(n100256) );
  NAND2_X1 U90295 ( .A1(n100259), .A2(n69323), .ZN(n100258) );
  NOR2_X1 U90296 ( .A1(n57379), .A2(n100260), .ZN(n100259) );
  AOI22_X1 U90297 ( .A1(n100261), .A2(n59326), .B1(n59323), .B2(
        \DLX_Datapath/IR_EXMEM[29] ), .ZN(n100260) );
  AOI21_X1 U90298 ( .B1(n59323), .B2(n106943), .A(\DLX_Datapath/IR_EXMEM[29] ), 
        .ZN(n100261) );
  AOI22_X1 U90299 ( .A1(n107148), .A2(n106940), .B1(n59326), .B2(n100262), 
        .ZN(n100257) );
  NAND2_X1 U90300 ( .A1(\DLX_Datapath/IR_EXMEM[27] ), .A2(n111022), .ZN(
        n100262) );
  NOR4_X1 U90301 ( .A1(n100263), .A2(n100264), .A3(n100265), .A4(n100266), 
        .ZN(n100234) );
  XOR2_X1 U90302 ( .A(n86281), .B(n100217), .Z(n100266) );
  XOR2_X1 U90303 ( .A(n99344), .B(n100220), .Z(n100265) );
  XOR2_X1 U90304 ( .A(n86284), .B(n100222), .Z(n100264) );
  XOR2_X1 U90305 ( .A(n100893), .B(n64267), .Z(n100263) );
  NAND2_X1 U90306 ( .A1(n99323), .A2(n100199), .ZN(n100225) );
  NOR4_X1 U90308 ( .A1(n100269), .A2(n100270), .A3(n100271), .A4(n100272), 
        .ZN(n100268) );
  XOR2_X1 U90309 ( .A(n100893), .B(n54620), .Z(n100272) );
  XOR2_X1 U90310 ( .A(n100429), .B(n100630), .Z(n100271) );
  XOR2_X1 U90311 ( .A(n100430), .B(n100631), .Z(n100270) );
  XOR2_X1 U90312 ( .A(n100428), .B(n100632), .Z(n100269) );
  XOR2_X1 U90314 ( .A(n86295), .B(n100222), .Z(n100275) );
  OAI21_X1 U90315 ( .B1(n61799), .B2(n100276), .A(n100277), .ZN(n100222) );
  NOR2_X1 U90316 ( .A1(n100278), .A2(n107108), .ZN(n100277) );
  OAI21_X1 U90318 ( .B1(n107143), .B2(n105037), .A(n100280), .ZN(n86295) );
  XOR2_X1 U90319 ( .A(n107109), .B(n100281), .Z(n100280) );
  NAND2_X1 U90320 ( .A1(n100282), .A2(n107107), .ZN(n100281) );
  XOR2_X1 U90321 ( .A(n100217), .B(n86296), .Z(n100274) );
  OAI21_X1 U90322 ( .B1(n107143), .B2(n105037), .A(n100283), .ZN(n86296) );
  XOR2_X1 U90323 ( .A(n100282), .B(n107107), .Z(n100283) );
  NAND2_X1 U90324 ( .A1(n100284), .A2(n100285), .ZN(n100217) );
  AOI21_X1 U90325 ( .B1(n105052), .B2(n111028), .A(n81901), .ZN(n100285) );
  AOI22_X1 U90326 ( .A1(n61799), .A2(n105012), .B1(n61799), .B2(n100893), .ZN(
        n100284) );
  OAI21_X1 U90328 ( .B1(n61799), .B2(n59516), .A(n100286), .ZN(n100220) );
  OAI21_X1 U90329 ( .B1(n59516), .B2(n100893), .A(n61799), .ZN(n100286) );
  NOR2_X1 U90330 ( .A1(n100282), .A2(n100287), .ZN(n86297) );
  AOI21_X1 U90331 ( .B1(n105037), .B2(n107105), .A(n107143), .ZN(n100287) );
  NOR2_X1 U90332 ( .A1(n100892), .A2(n58722), .ZN(n100282) );
  NOR4_X1 U90333 ( .A1(n69380), .A2(n69319), .A3(n111054), .A4(n100288), .ZN(
        n99323) );
  XOR2_X1 U90334 ( .A(n69378), .B(n100289), .Z(n100288) );
  NOR2_X1 U90335 ( .A1(n69324), .A2(n100762), .ZN(n100289) );
  AOI22_X1 U90336 ( .A1(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[0] ), .A2(
        n105103), .B1(n107569), .B2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .ZN(n100187) );
  NAND2_X1 U90337 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [0]), .A2(n108857), 
        .ZN(n99851) );
  NOR2_X1 U90338 ( .A1(n108857), .A2(n99849), .ZN(n99764) );
  NOR2_X1 U90339 ( .A1(n108857), .A2(\DLX_Datapath/ArithLogUnit/B_mul [0]), 
        .ZN(n99849) );
  NAND2_X1 U90340 ( .A1(n105196), .A2(n105900), .ZN(
        \DLX_Datapath/ArithLogUnit/N112 ) );
  NOR4_X1 U90341 ( .A1(n69330), .A2(n107422), .A3(n107423), .A4(n99001), .ZN(
        n81804) );
  NAND2_X1 U90342 ( .A1(n105227), .A2(n105197), .ZN(n81805) );
  NAND2_X1 U90343 ( .A1(n106359), .A2(n98995), .ZN(
        \DLX_Datapath/ArithLogUnit/N177 ) );
  OR2_X1 U90344 ( .A1(n98973), .A2(n98999), .ZN(n98995) );
  NOR2_X1 U90345 ( .A1(n100290), .A2(n100291), .ZN(n60159) );
  OAI21_X1 U90346 ( .B1(n98978), .B2(n106956), .A(n106955), .ZN(n100291) );
  NOR4_X1 U90347 ( .A1(n69801), .A2(n69330), .A3(n107422), .A4(n99001), .ZN(
        n100292) );
  NAND2_X1 U90348 ( .A1(n98980), .A2(n99003), .ZN(n100290) );
  AOI22_X1 U90351 ( .A1(n69802), .A2(n98976), .B1(n107424), .B2(n98978), .ZN(
        n100295) );
  NAND2_X1 U90352 ( .A1(n100296), .A2(n69801), .ZN(n98978) );
  NOR2_X1 U90353 ( .A1(n106953), .A2(n107422), .ZN(n100296) );
  NAND2_X1 U90355 ( .A1(n100297), .A2(n69801), .ZN(n98971) );
  NOR2_X1 U90356 ( .A1(n69800), .A2(n106953), .ZN(n100297) );
  NAND2_X1 U90357 ( .A1(n100298), .A2(n69800), .ZN(n98973) );
  NOR2_X1 U90358 ( .A1(n69801), .A2(n106953), .ZN(n100298) );
  NAND2_X1 U90360 ( .A1(n107424), .A2(n106956), .ZN(n99001) );
  NOR2_X1 U90362 ( .A1(n98999), .A2(n98976), .ZN(n98996) );
  NAND2_X1 U90363 ( .A1(n100300), .A2(n69330), .ZN(n98976) );
  NOR2_X1 U90364 ( .A1(n69801), .A2(n69800), .ZN(n100300) );
  NAND2_X1 U90365 ( .A1(n69802), .A2(n106956), .ZN(n98999) );
  NOR2_X1 U90366 ( .A1(net113156), .A2(n111029), .ZN(\DLX_ControlUnit/N2798 )
         );
  NOR2_X1 U90367 ( .A1(net113159), .A2(n111030), .ZN(\DLX_ControlUnit/N2789 )
         );
  NOR2_X1 U90368 ( .A1(net113155), .A2(n111031), .ZN(\DLX_ControlUnit/N2787 )
         );
  NOR2_X1 U90369 ( .A1(net113156), .A2(n111032), .ZN(\DLX_ControlUnit/N2785 )
         );
  NAND2_X1 U90370 ( .A1(n100301), .A2(n100302), .ZN(n80001) );
  AOI21_X1 U90371 ( .B1(n100303), .B2(n100304), .A(n100305), .ZN(n100302) );
  OR2_X1 U90372 ( .A1(FILL), .A2(SPILL), .ZN(n100305) );
  OAI21_X1 U90373 ( .B1(n111026), .B2(n106327), .A(n81888), .ZN(SPILL) );
  NAND2_X1 U90374 ( .A1(n81903), .A2(n106958), .ZN(n81888) );
  NOR2_X1 U90375 ( .A1(n106695), .A2(n81915), .ZN(n81903) );
  NAND2_X1 U90376 ( .A1(n100306), .A2(n100307), .ZN(n81915) );
  XOR2_X1 U90377 ( .A(n100308), .B(n59518), .Z(n100307) );
  NAND2_X1 U90378 ( .A1(n81909), .A2(n86228), .ZN(n100308) );
  NAND2_X1 U90379 ( .A1(n59515), .A2(n59514), .ZN(n86228) );
  NAND2_X1 U90380 ( .A1(n106764), .A2(n106753), .ZN(n81909) );
  NOR2_X1 U90381 ( .A1(n106762), .A2(n100309), .ZN(n100306) );
  NAND2_X1 U90382 ( .A1(n100717), .A2(n107021), .ZN(n80203) );
  NAND2_X1 U90383 ( .A1(n98368), .A2(n86300), .ZN(FILL) );
  OR2_X1 U90384 ( .A1(n100311), .A2(n106957), .ZN(n86300) );
  NAND2_X1 U90385 ( .A1(n106958), .A2(n81882), .ZN(n100311) );
  NOR4_X1 U90386 ( .A1(n69283), .A2(n100309), .A3(n100310), .A4(n100312), .ZN(
        n81882) );
  XOR2_X1 U90387 ( .A(n59518), .B(n59515), .Z(n100312) );
  XNOR2_X1 U90388 ( .A(n106764), .B(n59517), .ZN(n100310) );
  XOR2_X1 U90389 ( .A(n59516), .B(
        \dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .Z(n100309) );
  NAND2_X1 U90390 ( .A1(n107023), .A2(n107021), .ZN(n86222) );
  NAND2_X1 U90391 ( .A1(n105206), .A2(n86230), .ZN(n98368) );
  NAND2_X1 U90392 ( .A1(n62212), .A2(n62190), .ZN(n86230) );
  NAND2_X1 U90393 ( .A1(n69343), .A2(n107023), .ZN(n94366) );
  NOR4_X1 U90394 ( .A1(n100313), .A2(n100314), .A3(n100315), .A4(n100316), 
        .ZN(n100304) );
  XOR2_X1 U90395 ( .A(n64247), .B(n59453), .Z(n100316) );
  XOR2_X1 U90396 ( .A(n100427), .B(n59452), .Z(n100315) );
  AOI22_X1 U90398 ( .A1(n100317), .A2(n100318), .B1(n100228), .B2(n106846), 
        .ZN(n100313) );
  NOR3_X1 U90399 ( .A1(n100320), .A2(n100321), .A3(n100322), .ZN(n100319) );
  NOR2_X1 U90400 ( .A1(n69321), .A2(n100323), .ZN(n100322) );
  AOI21_X1 U90401 ( .B1(n100324), .B2(n106942), .A(n100325), .ZN(n100323) );
  NOR3_X1 U90402 ( .A1(n100326), .A2(n69313), .A3(n107149), .ZN(n100325) );
  XOR2_X1 U90403 ( .A(n69377), .B(n69325), .Z(n100326) );
  NOR3_X1 U90404 ( .A1(n104498), .A2(n100327), .A3(n106847), .ZN(n100321) );
  XOR2_X1 U90405 ( .A(n104496), .B(n69321), .Z(n100327) );
  OAI21_X1 U90406 ( .B1(n100328), .B2(n106936), .A(n100329), .ZN(n100320) );
  OAI21_X1 U90407 ( .B1(n100330), .B2(n100331), .A(n107149), .ZN(n100329) );
  OAI33_X1 U90408 ( .A1(n106936), .A2(n69377), .A3(n69325), .B1(n104496), .B2(
        n69379), .B3(n106847), .ZN(n100331) );
  AOI21_X1 U90409 ( .B1(n100332), .B2(n69321), .A(n104498), .ZN(n100330) );
  AOI21_X1 U90410 ( .B1(n106847), .B2(n106942), .A(n104496), .ZN(n100332) );
  OAI21_X1 U90411 ( .B1(\DLX_Datapath/IR_IDEX[31] ), .B2(n106880), .A(n106848), 
        .ZN(n100317) );
  OAI21_X1 U90412 ( .B1(\DLX_Datapath/IR_IDEX[31] ), .B2(n100333), .A(n100334), 
        .ZN(n100232) );
  NAND2_X1 U90413 ( .A1(n69315), .A2(n100335), .ZN(n100334) );
  OAI21_X1 U90414 ( .B1(n100336), .B2(n106937), .A(n100233), .ZN(n100335) );
  NAND2_X1 U90415 ( .A1(n100337), .A2(\DLX_Datapath/IR_IDEX[27] ), .ZN(n100233) );
  NOR2_X1 U90416 ( .A1(n69322), .A2(n59417), .ZN(n100337) );
  AOI22_X1 U90417 ( .A1(n100338), .A2(n59419), .B1(n59415), .B2(
        \DLX_Datapath/IR_IDEX[29] ), .ZN(n100336) );
  NAND2_X1 U90419 ( .A1(n69326), .A2(n59415), .ZN(n83104) );
  NAND2_X1 U90420 ( .A1(n59415), .A2(\DLX_Datapath/IR_IDEX[29] ), .ZN(n100333)
         );
  NOR2_X1 U90421 ( .A1(n59417), .A2(n69315), .ZN(n83102) );
  NOR4_X1 U90422 ( .A1(n100339), .A2(n100340), .A3(n100341), .A4(n100342), 
        .ZN(n100303) );
  XOR2_X1 U90423 ( .A(n100719), .B(n59451), .Z(n100342) );
  XOR2_X1 U90424 ( .A(n62496), .B(n59445), .Z(n100341) );
  XOR2_X1 U90425 ( .A(n104700), .B(n99339), .Z(n100340) );
  XOR2_X1 U90426 ( .A(n104786), .B(n107061), .Z(n100339) );
  AOI22_X1 U90427 ( .A1(n100343), .A2(n100344), .B1(n106932), .B2(n100318), 
        .ZN(n100301) );
  NAND2_X1 U90429 ( .A1(n100345), .A2(n100346), .ZN(n82280) );
  NOR3_X1 U90430 ( .A1(n69321), .A2(n69381), .A3(n69379), .ZN(n100346) );
  NOR2_X1 U90431 ( .A1(n106847), .A2(n104496), .ZN(n100345) );
  NOR2_X1 U90432 ( .A1(n106936), .A2(n106845), .ZN(n82656) );
  AOI22_X1 U90433 ( .A1(n100348), .A2(n100349), .B1(n100350), .B2(n100351), 
        .ZN(n100347) );
  NOR3_X1 U90434 ( .A1(\DLX_Datapath/IR_EXMEM[29] ), .A2(n59326), .A3(n100352), 
        .ZN(n100351) );
  XOR2_X1 U90435 ( .A(\DLX_Datapath/IR_EXMEM[27] ), .B(n100353), .Z(n100352)
         );
  NOR2_X1 U90436 ( .A1(n57378), .A2(n69323), .ZN(n100353) );
  NOR2_X1 U90437 ( .A1(n111022), .A2(n82678), .ZN(n100350) );
  NAND2_X1 U90438 ( .A1(n100354), .A2(n100355), .ZN(n82678) );
  XOR2_X1 U90440 ( .A(n99344), .B(n82687), .Z(n100359) );
  NAND2_X1 U90441 ( .A1(n104995), .A2(n100361), .ZN(n99344) );
  OAI21_X1 U90442 ( .B1(n107141), .B2(n104996), .A(n104874), .ZN(n100361) );
  XNOR2_X1 U90443 ( .A(n82694), .B(n86284), .ZN(n100358) );
  NAND2_X1 U90444 ( .A1(n100363), .A2(n100362), .ZN(n86284) );
  XOR2_X1 U90447 ( .A(n100422), .B(n59452), .Z(n100357) );
  XOR2_X1 U90448 ( .A(n64267), .B(n59453), .Z(n100356) );
  XOR2_X1 U90450 ( .A(n82688), .B(n86281), .Z(n100367) );
  NAND2_X1 U90451 ( .A1(n100368), .A2(n100362), .ZN(n86281) );
  NAND2_X1 U90452 ( .A1(n104874), .A2(n64267), .ZN(n100362) );
  XOR2_X1 U90455 ( .A(n100423), .B(n59451), .Z(n100366) );
  XOR2_X1 U90456 ( .A(n100796), .B(n59445), .Z(n100365) );
  NOR4_X1 U90457 ( .A1(n100231), .A2(n100369), .A3(n100370), .A4(n100371), 
        .ZN(n100349) );
  XOR2_X1 U90458 ( .A(n82687), .B(n100372), .Z(n100371) );
  OAI21_X1 U90459 ( .B1(n107096), .B2(\DLX_Datapath/IR_IDEX[15] ), .A(n100373), 
        .ZN(n100372) );
  OAI21_X1 U90460 ( .B1(n62574), .B2(\DLX_Datapath/IR_IDEX[15] ), .A(n107096), 
        .ZN(n100373) );
  NAND2_X1 U90461 ( .A1(n94068), .A2(n94253), .ZN(n82687) );
  XOR2_X1 U90463 ( .A(n104786), .B(n100374), .Z(n100370) );
  NOR3_X1 U90464 ( .A1(n100375), .A2(n100278), .A3(n100376), .ZN(n100374) );
  AOI21_X1 U90465 ( .B1(\DLX_Datapath/HazardDetUnit/N112 ), .B2(
        \DLX_Datapath/CWP_IDEX[2] ), .A(\DLX_Datapath/IR_IDEX[15] ), .ZN(
        n100376) );
  NOR2_X1 U90466 ( .A1(n62573), .A2(n100276), .ZN(n100375) );
  AOI21_X1 U90469 ( .B1(n104899), .B2(n104495), .A(n100278), .ZN(n100377) );
  XOR2_X1 U90470 ( .A(n104700), .B(n100378), .Z(n100369) );
  OAI21_X1 U90471 ( .B1(n62573), .B2(n81890), .A(n100379), .ZN(n100378) );
  NOR2_X1 U90472 ( .A1(n81901), .A2(n100380), .ZN(n100379) );
  AOI21_X1 U90473 ( .B1(\DLX_Datapath/HazardDetUnit/N112 ), .B2(n104898), .A(
        \DLX_Datapath/IR_IDEX[15] ), .ZN(n100380) );
  NOR2_X1 U90474 ( .A1(n104898), .A2(n107096), .ZN(n81901) );
  NAND2_X1 U90475 ( .A1(n94257), .A2(n94068), .ZN(n82688) );
  NAND2_X1 U90476 ( .A1(n59454), .A2(n59453), .ZN(n94068) );
  AOI21_X1 U90478 ( .B1(n81899), .B2(n104495), .A(n100382), .ZN(n100381) );
  NAND2_X1 U90479 ( .A1(n100383), .A2(n100384), .ZN(n100231) );
  NOR3_X1 U90480 ( .A1(n69315), .A2(n69326), .A3(n69322), .ZN(n100384) );
  NOR3_X1 U90481 ( .A1(\DLX_Datapath/IR_IDEX[31] ), .A2(
        \DLX_Datapath/IR_IDEX[27] ), .A3(\DLX_Datapath/IR_IDEX[29] ), .ZN(
        n100383) );
  NOR4_X1 U90482 ( .A1(n100385), .A2(n100386), .A3(n100387), .A4(n100388), 
        .ZN(n100348) );
  XOR2_X1 U90483 ( .A(n100426), .B(n59451), .Z(n100388) );
  XOR2_X1 U90484 ( .A(n100424), .B(n59445), .Z(n100387) );
  XOR2_X1 U90485 ( .A(n62574), .B(n59453), .Z(n100386) );
  NOR4_X1 U90487 ( .A1(n100389), .A2(n100390), .A3(n69325), .A4(n69321), .ZN(
        n100344) );
  AOI21_X1 U90488 ( .B1(n100391), .B2(n99339), .A(n90110), .ZN(n100390) );
  OAI21_X1 U90489 ( .B1(n62496), .B2(n107132), .A(n100392), .ZN(n100389) );
  AOI22_X1 U90490 ( .A1(n100393), .A2(n90110), .B1(n107061), .B2(n107060), 
        .ZN(n100392) );
  NAND2_X1 U90491 ( .A1(n100395), .A2(n100391), .ZN(n100393) );
  AOI22_X1 U90493 ( .A1(n62496), .A2(n107132), .B1(n100719), .B2(n107134), 
        .ZN(n100397) );
  AOI22_X1 U90494 ( .A1(n100427), .A2(n107137), .B1(n64247), .B2(n107139), 
        .ZN(n100396) );
  AOI22_X1 U90495 ( .A1(n90291), .A2(n99339), .B1(n100394), .B2(n99349), .ZN(
        n100395) );
  NAND2_X1 U90496 ( .A1(n100398), .A2(n100399), .ZN(n99349) );
  AOI22_X1 U90499 ( .A1(n104899), .A2(\DLX_Datapath/IR_IDEX[20] ), .B1(n64246), 
        .B2(n59518), .ZN(n100398) );
  XOR2_X1 U90501 ( .A(n100401), .B(n59518), .Z(n100394) );
  NAND2_X1 U90502 ( .A1(n105052), .A2(n107142), .ZN(n100401) );
  OAI21_X1 U90504 ( .B1(n100402), .B2(n107094), .A(n100400), .ZN(n99339) );
  AOI21_X1 U90505 ( .B1(\DLX_Datapath/IR_IDEX[20] ), .B2(n81899), .A(n100382), 
        .ZN(n100403) );
  NOR2_X1 U90506 ( .A1(n59517), .A2(\DLX_Datapath/IR_IDEX[20] ), .ZN(n100402)
         );
  OAI21_X1 U90507 ( .B1(n105012), .B2(n107142), .A(n100404), .ZN(n90291) );
  AOI21_X1 U90508 ( .B1(n105031), .B2(n107142), .A(n100382), .ZN(n100404) );
  NOR2_X1 U90510 ( .A1(n107106), .A2(n59516), .ZN(n81899) );
  NOR4_X1 U90511 ( .A1(n100405), .A2(n100406), .A3(n106845), .A4(n106933), 
        .ZN(n100343) );
  NOR4_X1 U90512 ( .A1(n69315), .A2(n59419), .A3(n100407), .A4(
        \DLX_Datapath/IR_IDEX[29] ), .ZN(n100228) );
  XOR2_X1 U90513 ( .A(n100408), .B(n59415), .Z(n100407) );
  NAND2_X1 U90514 ( .A1(n69326), .A2(n106937), .ZN(n100408) );
  NOR2_X1 U90515 ( .A1(n100328), .A2(n69381), .ZN(n100324) );
  NAND2_X1 U90516 ( .A1(n100409), .A2(n106847), .ZN(n100328) );
  NOR2_X1 U90517 ( .A1(n69379), .A2(n69377), .ZN(n100409) );
  XOR2_X1 U90518 ( .A(n99334), .B(n100410), .Z(n100406) );
  NOR2_X1 U90519 ( .A1(n107140), .A2(n90293), .ZN(n100410) );
  XOR2_X1 U90520 ( .A(n107142), .B(n59516), .Z(n90293) );
  NAND2_X1 U90521 ( .A1(n59444), .A2(n59443), .ZN(n90110) );
  XOR2_X1 U90522 ( .A(n100411), .B(n64246), .Z(n99334) );
  NAND2_X1 U90523 ( .A1(n107096), .A2(n100400), .ZN(n100411) );
  NAND2_X1 U90524 ( .A1(n64246), .A2(n64247), .ZN(n100400) );
  OAI21_X1 U90525 ( .B1(n64247), .B2(n107139), .A(n100412), .ZN(n100405) );
  AOI22_X1 U90526 ( .A1(n59441), .A2(\DLX_Datapath/HazardDetUnit/N96 ), .B1(
        n59442), .B2(\DLX_Datapath/HazardDetUnit/N97 ), .ZN(n100412) );
  DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW_sra_0 \DLX_Datapath/ArithLogUnit/ALU_shift/sra_39  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_shf ), .SH(
        \DLX_Datapath/ArithLogUnit/B_shf ), .SH_TC(1'b0), .B({
        \DLX_Datapath/ArithLogUnit/ALU_shift/N103 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N102 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N101 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N100 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N99 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N98 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N97 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N96 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N95 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N94 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N93 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N92 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N91 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N90 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N89 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N88 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N87 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N86 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N85 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N84 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N83 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N82 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N81 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N80 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N79 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N78 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N77 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N76 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N75 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N74 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N73 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N72 }) );
  DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW_rash_0 \DLX_Datapath/ArithLogUnit/ALU_shift/srl_39  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_shf ), .DATA_TC(1'b0), .SH(
        \DLX_Datapath/ArithLogUnit/B_shf ), .SH_TC(1'b0), .B({
        \DLX_Datapath/ArithLogUnit/ALU_shift/N71 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N70 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N69 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N68 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N67 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N66 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N65 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N64 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N63 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N62 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N61 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N60 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N59 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N58 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N57 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N56 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N55 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N54 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N53 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N52 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N51 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N50 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N49 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N48 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N47 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N46 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N45 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N44 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N43 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N42 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N41 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N40 }) );
  DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW01_ash_0 \DLX_Datapath/ArithLogUnit/ALU_shift/sll_39  ( 
        .A(\DLX_Datapath/ArithLogUnit/A_shf ), .DATA_TC(1'b0), .SH(
        \DLX_Datapath/ArithLogUnit/B_shf ), .SH_TC(1'b0), .B({
        \DLX_Datapath/ArithLogUnit/ALU_shift/N39 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N38 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N37 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N36 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N35 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N34 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N33 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N32 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N31 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N30 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N29 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N28 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N27 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N26 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N25 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N24 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N23 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N22 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N21 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N20 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N19 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N18 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N17 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N16 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N15 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N14 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N13 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N12 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N11 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N10 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N9 , 
        \DLX_Datapath/ArithLogUnit/ALU_shift/N8 }) );
  DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW01_inc_0 \DLX_Datapath/ArithLogUnit/ALU_mult/boothCalc/add_52  ( 
        .A({n108266, n108266, n108389, n108501, n107742, n109652, n108614, 
        n109759, n109545, n109082, n109429, n109313, n109204, n108737, n108966, 
        n108855, n107568, 1'b1}), .SUM({
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[17] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[16] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[15] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[13] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[12] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[11] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[10] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[9] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[7] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[6] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[5] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[4] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[3] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[2] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[1] , SYNOPSYS_UNCONNECTED__0}) );
  DLX_ADDR_SIZE32_DATA_SIZE32_IR_SIZE32_OPC_SIZE6_REGADDR_SIZE5_STACKBUS_WIDTH4_DW01_inc_1 \DLX_Datapath/ArithLogUnit/ALU_mult/boothCalc/add_50  ( 
        .A({n108266, n108266, n108266, n108389, n108501, n107742, n109652, 
        n108614, n109759, n109545, n109082, n109429, n109313, n109204, n108737, 
        n108966, n108855, n107568}), .SUM({
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[17] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[16] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[15] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[14] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[13] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[12] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[11] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[10] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[9] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[8] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[7] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[6] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[5] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[4] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[3] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[2] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[1] , 
        \DLX_Datapath/ArithLogUnit/ALU_mult/m_A[0] }) );
  NAND2_X1 U68045 ( .A1(IR_in[5]), .A2(n104755), .ZN(n81967) );
  AOI22_X1 U67722 ( .A1(n82423), .A2(n62200), .B1(n82424), .B2(n104755), .ZN(
        n82422) );
  SDFFR_X2 \DLX_ControlUnit/ALUop3_reg[4]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/ALUop2 [4]), .SE(net113091), .CK(Clk), .RN(Rst), .Q(
        n106953), .QN(n69330) );
  SDFFR_X2 \DLX_Datapath/IR_IDEX_reg[13]  ( .D(1'b0), .SI(net113091), .SE(
        \DLX_Datapath/IR_IFID[13] ), .CK(Clk), .RN(Rst), .Q(
        \DLX_Datapath/HazardDetUnit/N111 ) );
  SDFFR_X2 \DLX_ControlUnit/ALUop3_reg[2]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/ALUop2 [2]), .SE(n104753), .CK(Clk), .RN(Rst), .Q(
        n69802), .QN(n107424) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[11]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [11]), .SE(net113081), .CK(Clk), .RN(n106508), 
        .Q(\DLX_ControlUnit/cw3 [11]) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[2]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [2]), .SE(n104753), .CK(Clk), .RN(n106508), .Q(
        \DLX_ControlUnit/cw3 [2]) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[17]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [17]), .SE(net113091), .CK(Clk), .RN(n106508), 
        .Q(n61539) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[13]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [13]), .SE(net113102), .CK(Clk), .RN(n106508), 
        .Q(\DLX_ControlUnit/cw3 [13]) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[9]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [9]), .SE(net113153), .CK(Clk), .RN(Rst), .Q(
        \DLX_ControlUnit/cw3 [9]) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[15]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [15]), .SE(net113091), .CK(Clk), .RN(n106508), 
        .Q(n62027), .QN(n107413) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[12]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [12]), .SE(net113081), .CK(Clk), .RN(n106508), 
        .Q(\DLX_ControlUnit/cw3 [12]) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[7]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [7]), .SE(net113102), .CK(Clk), .RN(n106508), .Q(
        \DLX_ControlUnit/cw3 [7]) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[6]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [6]), .SE(n104753), .CK(Clk), .RN(n106508), .Q(
        \DLX_ControlUnit/cw3 [6]) );
  SDFFR_X2 \DLX_ControlUnit/ALUop3_reg[3]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/ALUop2 [3]), .SE(net113153), .CK(Clk), .RN(n106508), 
        .Q(n69339), .QN(n106956) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[10]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [10]), .SE(net113081), .CK(Clk), .RN(Rst), .Q(
        \DLX_ControlUnit/cw3 [10]) );
  SDFFR_X2 \DLX_ControlUnit/cw3_reg[0]  ( .D(1'b0), .SI(
        \DLX_ControlUnit/cw2 [0]), .SE(net113091), .CK(Clk), .RN(n106508), .Q(
        \DLX_ControlUnit/cw3 [0]) );
  DFF_X2 \DLX_Datapath/CWP_EXMEM_reg[2]  ( .D(n59069), .CK(Clk), .Q(n69348), 
        .QN(n104741) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[13]  ( .D(\DLX_ControlUnit/cw3 [13]), .CK(
        Clk), .RN(n106471), .Q(DRAM_WE) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[12]  ( .D(\DLX_ControlUnit/cw3 [12]), .CK(
        Clk), .RN(n106471), .Q(DRAM_RE) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[11]  ( .D(\DLX_ControlUnit/cw3 [11]), .CK(
        Clk), .RN(n106471), .Q(DRAMOP_SEL) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[10]  ( .D(\DLX_ControlUnit/cw3 [10]), .CK(
        Clk), .RN(n106465), .Q(n100415), .QN(n111050) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[9]  ( .D(\DLX_ControlUnit/cw3 [9]), .CK(Clk), .RN(n106465), .Q(n69698), .QN(n104450) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[7]  ( .D(\DLX_ControlUnit/cw3 [7]), .CK(Clk), .RN(n106465), .Q(n69697), .QN(n111053) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[6]  ( .D(\DLX_ControlUnit/cw3 [6]), .CK(Clk), .RN(n106465), .Q(n100414) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[2]  ( .D(\DLX_ControlUnit/cw3 [2]), .CK(Clk), .RN(n106471), .Q(\DLX_ControlUnit/cw4 [2]) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[0]  ( .D(\DLX_ControlUnit/cw3 [0]), .CK(Clk), .RN(n106471), .Q(\DLX_ControlUnit/cw4 [0]) );
  DFFR_X2 \DLX_Datapath/RegisterFile/old_CWP2_reg[2]  ( .D(
        \DLX_Datapath/RegisterFile/old_CWP1 [2]), .CK(Clk), .RN(n106470), .Q(
        \DLX_Datapath/RegisterFile/old_CWP2[2] ) );
  DFFR_X2 \DLX_Datapath/RegisterFile/old_CWP2_reg[1]  ( .D(
        \DLX_Datapath/RegisterFile/old_CWP1 [1]), .CK(Clk), .RN(n106470), .Q(
        \DLX_Datapath/RegisterFile/old_CWP2[1] ) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[31]  ( .D(\DLX_Datapath/IR_EXMEM[31] ), 
        .CK(Clk), .RN(n106465), .Q(n69382), .QN(n111054) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[29]  ( .D(\DLX_Datapath/IR_EXMEM[29] ), 
        .CK(Clk), .RN(n106465), .Q(n69380) );
  DFFR_X2 \DLX_Datapath/IR_MEMWB_reg[27]  ( .D(\DLX_Datapath/IR_EXMEM[27] ), 
        .CK(Clk), .RN(n106465), .Q(n69378), .QN(n111055) );
  DFFR_X2 \DLX_ControlUnit/cw5_reg[4]  ( .D(\DLX_ControlUnit/cw4 [4]), .CK(Clk), .RN(n106465), .Q(n69424), .QN(n111056) );
  DFFR_X2 \DLX_ControlUnit/cw5_reg[1]  ( .D(\DLX_ControlUnit/cw4 [1]), .CK(Clk), .RN(n106465), .Q(n64655), .QN(n111064) );
  DFFR_X2 \DLX_ControlUnit/cw5_reg[0]  ( .D(\DLX_ControlUnit/cw4 [0]), .CK(Clk), .RN(n106465), .Q(n100629) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[8]  ( .D(\DLX_ControlUnit/cw3 [8]), .CK(Clk), .RN(n106465), .Q(n104434), .QN(n111065) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[5]  ( .D(\DLX_ControlUnit/cw3 [5]), .CK(Clk), .RN(n106465), .Q(n64652) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[4]  ( .D(\DLX_ControlUnit/cw3 [4]), .CK(Clk), .RN(n106470), .Q(\DLX_ControlUnit/cw4 [4]) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[3]  ( .D(\DLX_ControlUnit/cw3 [3]), .CK(Clk), .RN(n106470), .Q(\DLX_ControlUnit/cw4 [3]) );
  DFFR_X2 \DLX_ControlUnit/cw4_reg[1]  ( .D(\DLX_ControlUnit/cw3 [1]), .CK(Clk), .RN(n106470), .Q(\DLX_ControlUnit/cw4 [1]) );
  DFFR_X2 \DLX_Datapath/RegisterFile/old_CWP1_reg[2]  ( .D(
        \DLX_Datapath/CWP_IDEX[2] ), .CK(Clk), .RN(n106469), .Q(
        \DLX_Datapath/RegisterFile/old_CWP1 [2]) );
  DFFR_X2 \DLX_Datapath/RegisterFile/old_CWP1_reg[1]  ( .D(n104898), .CK(Clk), 
        .RN(n106469), .Q(\DLX_Datapath/RegisterFile/old_CWP1 [1]) );
  DFFR_X2 \DLX_Datapath/RegisterFile/old_CWP1_reg[0]  ( .D(n107096), .CK(Clk), 
        .RN(n106469), .Q(\DLX_Datapath/RegisterFile/old_CWP1 [0]) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[0]  ( .D(n59080), .CK(Clk), .RN(n106462), 
        .QN(n111106) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[1]  ( .D(n58951), .CK(Clk), .RN(n106462), 
        .QN(n111109) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[2]  ( .D(n58950), .CK(Clk), .RN(n106462), 
        .QN(n111108) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[3]  ( .D(n58949), .CK(Clk), .RN(n106462), 
        .QN(n111107) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[31]  ( .D(n59041), .CK(Clk), .RN(Rst), 
        .Q(n69708), .QN(n107370) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[30]  ( .D(n59040), .CK(Clk), .RN(Rst), 
        .Q(n69709), .QN(n107372) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[29]  ( .D(n59039), .CK(Clk), .RN(Rst), 
        .Q(n69710), .QN(n107374) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[28]  ( .D(n59038), .CK(Clk), .RN(Rst), 
        .Q(n69711), .QN(n107375) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[20]  ( .D(n59030), .CK(Clk), .RN(Rst), 
        .Q(n69719), .QN(n107391) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[18]  ( .D(n59028), .CK(Clk), .RN(Rst), 
        .Q(n69721), .QN(n107395) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[17]  ( .D(n59027), .CK(Clk), .RN(Rst), 
        .Q(n69722), .QN(n107397) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[16]  ( .D(n59026), .CK(Clk), .RN(Rst), 
        .Q(n69723), .QN(n107399) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[4]  ( .D(n58931), .CK(Clk), .RN(n106475), 
        .QN(n111115) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[8]  ( .D(n58917), .CK(Clk), .RN(n106462), 
        .QN(n111112) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[12]  ( .D(n59008), .CK(Clk), .RN(n106429), .QN(n107631) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[15]  ( .D(n59025), .CK(Clk), .RN(Rst), 
        .Q(n69724), .QN(n107401) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[13]  ( .D(n59023), .CK(Clk), .RN(n106430), .Q(n69726), .QN(n107405) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[12]  ( .D(n59022), .CK(Clk), .RN(n106430), .Q(n69727), .QN(n107407) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[11]  ( .D(n59021), .CK(Clk), .RN(n106430), .Q(n69728), .QN(n107409) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[14]  ( .D(n59024), .CK(Clk), .RN(Rst), 
        .Q(n69725), .QN(n107403) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[10]  ( .D(n59020), .CK(Clk), .RN(n106430), .Q(n69729), .QN(n107411) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[9]  ( .D(n59043), .CK(Clk), .RN(Rst), 
        .Q(n69706), .QN(n107366) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[8]  ( .D(n59042), .CK(Clk), .RN(Rst), 
        .Q(n69707), .QN(n107368) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[7]  ( .D(n59019), .CK(Clk), .RN(n106463), 
        .Q(n69730), .QN(n111098) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[6]  ( .D(n59050), .CK(Clk), .RN(n106463), 
        .Q(n69699), .QN(n111099) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[5]  ( .D(n59049), .CK(Clk), .RN(n106463), 
        .Q(n69700), .QN(n111100) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[4]  ( .D(n59048), .CK(Clk), .RN(n106463), 
        .Q(n69701), .QN(n111101) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[3]  ( .D(n59047), .CK(Clk), .RN(n106462), 
        .Q(n69702), .QN(n111102) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[2]  ( .D(n59046), .CK(Clk), .RN(n106462), 
        .Q(n69703), .QN(n111103) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[1]  ( .D(n59045), .CK(Clk), .RN(n106462), 
        .Q(n69704), .QN(n111104) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[0]  ( .D(n59044), .CK(Clk), .RN(n106462), 
        .Q(n69705), .QN(n111105) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[27]  ( .D(n59037), .CK(Clk), .RN(Rst), 
        .Q(n69712), .QN(n107377) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[26]  ( .D(n59036), .CK(Clk), .RN(Rst), 
        .Q(n69713), .QN(n107379) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[25]  ( .D(n59035), .CK(Clk), .RN(Rst), 
        .Q(n69714), .QN(n107381) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[24]  ( .D(n59034), .CK(Clk), .RN(Rst), 
        .Q(n69715), .QN(n107383) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[23]  ( .D(n59033), .CK(Clk), .RN(Rst), 
        .Q(n69716), .QN(n107385) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[22]  ( .D(n59032), .CK(Clk), .RN(Rst), 
        .Q(n69717), .QN(n107387) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[21]  ( .D(n59031), .CK(Clk), .RN(Rst), 
        .Q(n69718), .QN(n107389) );
  DFFR_X2 \DLX_Datapath/LMD_MEMWB_reg[19]  ( .D(n59029), .CK(Clk), .RN(Rst), 
        .Q(n69720), .QN(n107393) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[16]  ( .D(n58901), .CK(Clk), .RN(Rst), 
        .QN(n109785) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[9]  ( .D(n58911), .CK(Clk), .RN(n106462), 
        .QN(n111111) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[13]  ( .D(n58968), .CK(Clk), .RN(n106387), .QN(n108282) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[5]  ( .D(n58927), .CK(Clk), .RN(n106457), 
        .QN(n111114) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[6]  ( .D(n58923), .CK(Clk), .RN(n106462), 
        .QN(n111113) );
  DFFR_X2 \DLX_Datapath/RegisterFile/RF_state_reg[1]  ( .D(n60377), .CK(Clk), 
        .RN(Rst), .Q(n69343), .QN(n107021) );
  DFFR_X2 \DLX_Datapath/RegisterFile/RF_state_reg[0]  ( .D(n60375), .CK(Clk), 
        .RN(Rst), .Q(n100717), .QN(n107023) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[20]  ( .D(n58878), .CK(Clk), .RN(Rst), 
        .QN(n110338) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[17]  ( .D(n58895), .CK(Clk), .RN(n106507), .QN(n109903) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[7]  ( .D(n58938), .CK(Clk), .RN(n106403), 
        .QN(n108975) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[10]  ( .D(n58957), .CK(Clk), .RN(n106414), .QN(n108510) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[14]  ( .D(n58967), .CK(Clk), .RN(n106467), .QN(n111117) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[11]  ( .D(n58913), .CK(Clk), .RN(n106462), .QN(n111110) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[15]  ( .D(n58975), .CK(Clk), .RN(n106458), .QN(n111116) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[18]  ( .D(n58891), .CK(Clk), .RN(n106497), .QN(n110120) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[19]  ( .D(n58893), .CK(Clk), .RN(n106444), .QN(n110012) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[24]  ( .D(n58866), .CK(Clk), .RN(n106477), .QN(n110852) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[21]  ( .D(n58872), .CK(Clk), .RN(Rst), 
        .QN(n110547) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[22]  ( .D(n58884), .CK(Clk), .RN(Rst), 
        .QN(n110230) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[23]  ( .D(n58874), .CK(Clk), .RN(Rst), 
        .QN(n110447) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[28]  ( .D(n59001), .CK(Clk), .RN(Rst), 
        .QN(n107751) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[25]  ( .D(n58868), .CK(Clk), .RN(Rst), 
        .QN(n110751) );
  DFFR_X2 \DLX_ControlUnit/cw3_reg[5]  ( .D(\DLX_ControlUnit/N2789 ), .CK(Clk), 
        .RN(n106468), .Q(\DLX_ControlUnit/cw3 [5]) );
  DFFR_X2 \DLX_ControlUnit/ALUop3_reg[1]  ( .D(n103926), .CK(Clk), .RN(n106429), .Q(n69801), .QN(n107423) );
  DFFR_X2 \DLX_ControlUnit/cw3_reg[4]  ( .D(n103924), .CK(Clk), .RN(n106468), 
        .Q(\DLX_ControlUnit/cw3 [4]) );
  DFFR_X2 \DLX_ControlUnit/cw3_reg[16]  ( .D(n103925), .CK(Clk), .RN(n106430), 
        .Q(n62189) );
  DFFR_X2 \DLX_ControlUnit/cw3_reg[14]  ( .D(\DLX_ControlUnit/N2798 ), .CK(Clk), .RN(Rst), .Q(n100417) );
  DFFR_X2 \DLX_ControlUnit/cw3_reg[1]  ( .D(\DLX_ControlUnit/N2785 ), .CK(Clk), 
        .RN(n106469), .Q(\DLX_ControlUnit/cw3 [1]) );
  DFFR_X2 \DLX_ControlUnit/ALUop3_reg[0]  ( .D(n103922), .CK(Clk), .RN(n106429), .Q(n69800), .QN(n107422) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[29]  ( .D(n59077), .CK(Clk), .RN(Rst), 
        .QN(n106837) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[26]  ( .D(n58984), .CK(Clk), .RN(n106439), .QN(n108053) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[27]  ( .D(n58870), .CK(Clk), .RN(Rst), 
        .QN(n110654) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[30]  ( .D(n59002), .CK(Clk), .RN(Rst), 
        .QN(n107750) );
  DFFR_X2 \DLX_ControlUnit/cw3_reg[3]  ( .D(\DLX_ControlUnit/N2787 ), .CK(Clk), 
        .RN(n106468), .Q(\DLX_ControlUnit/cw3 [3]) );
  DFFR_X2 \DLX_ControlUnit/cw3_reg[8]  ( .D(n103923), .CK(Clk), .RN(n106468), 
        .Q(\DLX_ControlUnit/cw3 [8]) );
  DFFR_X2 \DLX_Datapath/LPC_MEMWB_reg[31]  ( .D(n59003), .CK(Clk), .RN(Rst), 
        .QN(n107749) );
  DFFR_X2 \DLX_ControlUnit/ALUop2_reg[2]  ( .D(n59090), .CK(Clk), .RN(n106429), 
        .Q(\DLX_ControlUnit/ALUop2 [2]) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[23]  ( .D(n59082), .CK(Clk), .RN(Rst), .Q(
        n100496) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[24]  ( .D(n59088), .CK(Clk), .RN(Rst), .Q(
        n61670) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[3]  ( .D(n60364), .CK(Clk), .RN(n106468), 
        .QN(n111031) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[18]  ( .D(n60358), .CK(Clk), .RN(Rst), .Q(
        n100718), .QN(n107151) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[14]  ( .D(n60360), .CK(Clk), .RN(n106468), 
        .QN(n111029) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[5]  ( .D(n60362), .CK(Clk), .RN(n106468), 
        .QN(n111030) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[1]  ( .D(n60365), .CK(Clk), .RN(n106468), 
        .QN(n111032) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26826 ), .CK(Clk), .RN(n106426), .Q(n70424), .QN(n107945) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26825 ), .CK(Clk), .RN(Rst), .Q(n70566), 
        .QN(n108041) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26824 ), .CK(Clk), .RN(Rst), .Q(n69425), 
        .QN(n107166) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26823 ), .CK(Clk), .RN(n106448), .Q(n70280), .QN(n107850) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26822 ), .CK(Clk), .RN(n106473), .Q(n74126), .QN(n110745) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26821 ), .CK(Clk), .RN(Rst), .Q(n70713), 
        .QN(n108150) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26820 ), .CK(Clk), .RN(n106477), .Q(n74267), .QN(n110848) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26819 ), .CK(Clk), .RN(n106418), .Q(n74407), .QN(n110949) );
  DFFR_X2 \DLX_ControlUnit/RMLcw2_reg[1]  ( .D(n103928), .CK(Clk), .RN(n106503), .Q(n69283), .QN(n106695) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26818 ), .CK(Clk), .RN(Rst), .Q(n73843), 
        .QN(n110542) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26817 ), .CK(Clk), .RN(n106406), .Q(n73547), .QN(n110327) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26816 ), .CK(Clk), .RN(n106412), .Q(n73984), .QN(n110647) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26815 ), .CK(Clk), .RN(n106450), .Q(n73696), .QN(n110436) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26814 ), .CK(Clk), .RN(n106498), .Q(n73258), .QN(n110114) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26813 ), .CK(Clk), .RN(n106456), .Q(n73400), .QN(n110221) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26812 ), .CK(Clk), .RN(Rst), .Q(n73116), 
        .QN(n110006) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26811 ), .CK(Clk), .RN(Rst), .Q(n72966), 
        .QN(n109889) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26810 ), .CK(Clk), .RN(n106389), .Q(n70862), .QN(n108263) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26809 ), .CK(Clk), .RN(Rst), .Q(n71021), 
        .QN(n108386) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26808 ), .CK(Clk), .RN(n106375), .Q(n71166), .QN(n108497) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26807 ), .CK(Clk), .RN(Rst), .Q(n70127), 
        .QN(n107734) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26806 ), .CK(Clk), .RN(n106485), .Q(n72656), .QN(n109649) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26805 ), .CK(Clk), .RN(Rst), .Q(n71315), 
        .QN(n108611) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26804 ), .CK(Clk), .RN(n106371), .Q(n72798), .QN(n109756) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26803 ), .CK(Clk), .RN(n106479), .Q(n72508), .QN(n109541) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26802 ), .CK(Clk), .RN(Rst), .Q(n71908), 
        .QN(n109079) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26801 ), .CK(Clk), .RN(Rst), .Q(n72357), 
        .QN(n109426) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26800 ), .CK(Clk), .RN(n106488), .Q(n72206), .QN(n109307) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26799 ), .CK(Clk), .RN(n106405), .Q(n72062), .QN(n109199) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26798 ), .CK(Clk), .RN(n106420), .Q(n71464), .QN(n108734) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26797 ), .CK(Clk), .RN(n106404), .Q(n71759), .QN(n108962) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26796 ), .CK(Clk), .RN(Rst), .Q(n71615), 
        .QN(n108850) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[2][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26795 ), .CK(Clk), .RN(Rst), .Q(n69426), 
        .QN(n107167) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25718 ), .CK(Clk), .RN(Rst), .Q(n72527) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25712 ), .CK(Clk), .RN(Rst), .Q(n72077) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25707 ), .CK(Clk), .RN(Rst), .Q(n69595) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25728 ), .CK(Clk), .RN(n106452), .Q(n73855) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][29]  ( .D(n104225), 
        .CK(Clk), .RN(n106443), .Q(n69492) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25644 ), .CK(Clk), .RN(n106486), .Q(n71488) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][30]  ( .D(n104224), 
        .CK(Clk), .RN(Rst), .Q(n70439) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25653 ), .CK(Clk), .RN(n106407), .Q(n71188) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25651 ), .CK(Clk), .RN(n106489), .Q(n72381) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25646 ), .CK(Clk), .RN(n106382), .Q(n71337) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25738 ), .CK(Clk), .RN(n106447), .Q(n70295) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][29]  ( .D(n104314), 
        .CK(Clk), .RN(Rst), .Q(n69490) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25719 ), .CK(Clk), .RN(Rst), .Q(n69998) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25737 ), .CK(Clk), .RN(Rst), .Q(n70437) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25733 ), .CK(Clk), .RN(n106438), .Q(n70584) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25714 ), .CK(Clk), .RN(n106403), .Q(n71779) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25711 ), .CK(Clk), .RN(n106483), .Q(n71933) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25710 ), .CK(Clk), .RN(n106382), .Q(n71335) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25709 ), .CK(Clk), .RN(n106428), .Q(n71630) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25668 ), .CK(Clk), .RN(Rst), .Q(n74140) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25665 ), .CK(Clk), .RN(n106455), .Q(n73420) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25664 ), .CK(Clk), .RN(n106453), .Q(n73857) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25660 ), .CK(Clk), .RN(n106406), .Q(n72989) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25655 ), .CK(Clk), .RN(Rst), .Q(n70000) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][25]  ( .D(n104315), 
        .CK(Clk), .RN(Rst), .Q(n74138) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25729 ), .CK(Clk), .RN(n106455), .Q(n73418) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25724 ), .CK(Clk), .RN(n106371), .Q(n72987) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25720 ), .CK(Clk), .RN(n106395), .Q(n71037) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25731 ), .CK(Clk), .RN(Rst), .Q(n74278) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25725 ), .CK(Clk), .RN(n106497), .Q(n73271) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25723 ), .CK(Clk), .RN(n106503), .Q(n72837) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][31]  ( .D(n104223), 
        .CK(Clk), .RN(n106447), .Q(n70297) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25650 ), .CK(Clk), .RN(n106402), .Q(n71781) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25671 ), .CK(Clk), .RN(Rst), .Q(n70153) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25670 ), .CK(Clk), .RN(n106413), .Q(n73999) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25669 ), .CK(Clk), .RN(n106438), .Q(n70586) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][15]  ( .D(n104222), 
        .CK(Clk), .RN(Rst), .Q(n70735) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25654 ), .CK(Clk), .RN(Rst), .Q(n72529) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25652 ), .CK(Clk), .RN(n106484), .Q(n72671) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25649 ), .CK(Clk), .RN(Rst), .Q(n72230) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25648 ), .CK(Clk), .RN(n106488), .Q(n72079) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25647 ), .CK(Clk), .RN(n106482), .Q(n71935) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][2]  ( .D(n104221), 
        .CK(Clk), .RN(n106428), .Q(n71632) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25643 ), .CK(Clk), .RN(Rst), .Q(n69597) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25735 ), .CK(Clk), .RN(Rst), .Q(n70151) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25734 ), .CK(Clk), .RN(Rst), .Q(n73997) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][10]  ( .D(n104313), 
        .CK(Clk), .RN(n106412), .Q(n71186) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25716 ), .CK(Clk), .RN(n106484), .Q(n72669) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25715 ), .CK(Clk), .RN(n106489), .Q(n72379) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][6]  ( .D(n104312), 
        .CK(Clk), .RN(Rst), .Q(n72228) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25708 ), .CK(Clk), .RN(n106443), .Q(n71486) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25667 ), .CK(Clk), .RN(Rst), .Q(n74280) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25662 ), .CK(Clk), .RN(Rst), .Q(n73131) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25666 ), .CK(Clk), .RN(n106402), .Q(n73716) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25663 ), .CK(Clk), .RN(Rst), .Q(n73569) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25661 ), .CK(Clk), .RN(n106497), .Q(n73273) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25659 ), .CK(Clk), .RN(n106503), .Q(n72839) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25657 ), .CK(Clk), .RN(n106387), .Q(n70894) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[38][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25656 ), .CK(Clk), .RN(n106395), .Q(n71039) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25730 ), .CK(Clk), .RN(n106437), .Q(n73714) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25727 ), .CK(Clk), .RN(n106444), .Q(n73567) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25726 ), .CK(Clk), .RN(Rst), .Q(n73129) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25722 ), .CK(Clk), .RN(Rst), .Q(n70733) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[36][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25721 ), .CK(Clk), .RN(n106387), .Q(n70892) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23850 ), .CK(Clk), .RN(n106476), .Q(n70354) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23848 ), .CK(Clk), .RN(Rst), .Q(n69549) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23846 ), .CK(Clk), .RN(Rst), .Q(n74056) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23844 ), .CK(Clk), .RN(Rst), .Q(n74197) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23829 ), .CK(Clk), .RN(n106375), .Q(n71245) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][8]  ( .D(
        \DLX_Datapath/RegisterFile/N23827 ), .CK(Clk), .RN(n106481), .Q(n72438) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][6]  ( .D(
        \DLX_Datapath/RegisterFile/N23825 ), .CK(Clk), .RN(Rst), .Q(n72287) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][4]  ( .D(
        \DLX_Datapath/RegisterFile/N23823 ), .CK(Clk), .RN(n106408), .Q(n71992) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][2]  ( .D(
        \DLX_Datapath/RegisterFile/N23821 ), .CK(Clk), .RN(n106425), .Q(n71689) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][1]  ( .D(
        \DLX_Datapath/RegisterFile/N23820 ), .CK(Clk), .RN(n106416), .Q(n71545) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[73][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24553 ), .CK(Clk), .RN(Rst), .Q(n70474) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23849 ), .CK(Clk), .RN(n106468), .Q(n70496) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23847 ), .CK(Clk), .RN(n106417), .Q(n70210) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23845 ), .CK(Clk), .RN(n106377), .Q(n70643) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][24]  ( .D(
        \DLX_Datapath/RegisterFile/N23843 ), .CK(Clk), .RN(Rst), .Q(n74337) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][23]  ( .D(
        \DLX_Datapath/RegisterFile/N23842 ), .CK(Clk), .RN(n106497), .Q(n73773) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23828 ), .CK(Clk), .RN(n106505), .Q(n72728) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][7]  ( .D(
        \DLX_Datapath/RegisterFile/N23826 ), .CK(Clk), .RN(n106399), .Q(n71838) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][5]  ( .D(
        \DLX_Datapath/RegisterFile/N23824 ), .CK(Clk), .RN(n106487), .Q(n72136) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][3]  ( .D(
        \DLX_Datapath/RegisterFile/N23822 ), .CK(Clk), .RN(Rst), .Q(n71394) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][0]  ( .D(
        \DLX_Datapath/RegisterFile/N23819 ), .CK(Clk), .RN(Rst), .Q(n69654) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][22]  ( .D(
        \DLX_Datapath/RegisterFile/N23841 ), .CK(Clk), .RN(n106449), .Q(n73477) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][21]  ( .D(
        \DLX_Datapath/RegisterFile/N23840 ), .CK(Clk), .RN(n106453), .Q(n73914) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][20]  ( .D(
        \DLX_Datapath/RegisterFile/N23839 ), .CK(Clk), .RN(n106391), .Q(n73626) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][19]  ( .D(
        \DLX_Datapath/RegisterFile/N23838 ), .CK(Clk), .RN(Rst), .Q(n73188) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][18]  ( .D(
        \DLX_Datapath/RegisterFile/N23837 ), .CK(Clk), .RN(n106494), .Q(n73330) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][17]  ( .D(
        \DLX_Datapath/RegisterFile/N23836 ), .CK(Clk), .RN(n106435), .Q(n73046) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][16]  ( .D(
        \DLX_Datapath/RegisterFile/N23835 ), .CK(Clk), .RN(Rst), .Q(n72896) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][15]  ( .D(
        \DLX_Datapath/RegisterFile/N23834 ), .CK(Clk), .RN(n106392), .Q(n70792) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][14]  ( .D(
        \DLX_Datapath/RegisterFile/N23833 ), .CK(Clk), .RN(Rst), .Q(n70951) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][13]  ( .D(
        \DLX_Datapath/RegisterFile/N23832 ), .CK(Clk), .RN(n106373), .Q(n71096) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][12]  ( .D(
        \DLX_Datapath/RegisterFile/N23831 ), .CK(Clk), .RN(n106431), .Q(n70057) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[95][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23830 ), .CK(Clk), .RN(n106486), .Q(n72586) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][23]  ( .D(
        \DLX_Datapath/RegisterFile/N22562 ), .CK(Clk), .RN(n106449), .Q(n73813), .QN(n110518) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][24]  ( .D(
        \DLX_Datapath/RegisterFile/N22563 ), .CK(Clk), .RN(Rst), .Q(n74377), 
        .QN(n110925) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][22]  ( .D(
        \DLX_Datapath/RegisterFile/N22561 ), .CK(Clk), .RN(Rst), .Q(n73517), 
        .QN(n110303) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][21]  ( .D(
        \DLX_Datapath/RegisterFile/N22560 ), .CK(Clk), .RN(Rst), .Q(n73954), 
        .QN(n110623) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][20]  ( .D(
        \DLX_Datapath/RegisterFile/N22559 ), .CK(Clk), .RN(n106457), .Q(n73666), .QN(n110412) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][19]  ( .D(
        \DLX_Datapath/RegisterFile/N22558 ), .CK(Clk), .RN(Rst), .Q(n73228), 
        .QN(n110090) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][18]  ( .D(
        \DLX_Datapath/RegisterFile/N22557 ), .CK(Clk), .RN(Rst), .Q(n73370), 
        .QN(n110197) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][17]  ( .D(
        \DLX_Datapath/RegisterFile/N22556 ), .CK(Clk), .RN(n106461), .Q(n73086), .QN(n109982) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][16]  ( .D(
        \DLX_Datapath/RegisterFile/N22555 ), .CK(Clk), .RN(Rst), .Q(n72936), 
        .QN(n109865) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][15]  ( .D(
        \DLX_Datapath/RegisterFile/N22554 ), .CK(Clk), .RN(n106439), .Q(n70832), .QN(n108239) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][14]  ( .D(
        \DLX_Datapath/RegisterFile/N22553 ), .CK(Clk), .RN(n106396), .Q(n70991), .QN(n108362) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][13]  ( .D(
        \DLX_Datapath/RegisterFile/N22552 ), .CK(Clk), .RN(Rst), .Q(n71136), 
        .QN(n108473) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24581 ), .CK(Clk), .RN(Rst), .Q(n70620) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24576 ), .CK(Clk), .RN(Rst), .Q(n73891) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24573 ), .CK(Clk), .RN(n106495), .Q(n73307) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24571 ), .CK(Clk), .RN(n106500), .Q(n72873) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24579 ), .CK(Clk), .RN(Rst), .Q(n74314) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24566 ), .CK(Clk), .RN(Rst), .Q(n72563) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24562 ), .CK(Clk), .RN(n106400), .Q(n71815) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24560 ), .CK(Clk), .RN(n106421), .Q(n72113) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24559 ), .CK(Clk), .RN(n106410), .Q(n71969) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24558 ), .CK(Clk), .RN(n106379), .Q(n71371) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24557 ), .CK(Clk), .RN(Rst), .Q(n71666) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24563 ), .CK(Clk), .RN(n106482), .Q(n72415) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][29]  ( .D(n104140), 
        .CK(Clk), .RN(n106467), .Q(n69526) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24583 ), .CK(Clk), .RN(n106497), .Q(n70187) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][27]  ( .D(n104139), 
        .CK(Clk), .RN(n106471), .Q(n74033) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24572 ), .CK(Clk), .RN(Rst), .Q(n73023) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24580 ), .CK(Clk), .RN(n106471), .Q(n74174) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24578 ), .CK(Clk), .RN(Rst), .Q(n73750) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24585 ), .CK(Clk), .RN(Rst), .Q(n70473) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[15]  ( .D(n106589), .CK(Clk), .RN(Rst), 
        .Q(n69369), .QN(n107130) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[6]  ( .D(n106579), .CK(Clk), .RN(Rst), .Q(
        n69355), .QN(n107111) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[12]  ( .D(n106555), .CK(Clk), .RN(n106467), 
        .Q(\DLX_ControlUnit/cw2 [12]) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[8]  ( .D(n106568), .CK(Clk), .RN(Rst), .Q(
        n69357), .QN(n107112) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[2]  ( .D(n106593), .CK(Clk), .RN(Rst), .Q(
        n69351), .QN(n107110) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[7]  ( .D(n106573), .CK(Clk), .RN(n106467), 
        .Q(\DLX_ControlUnit/cw2 [7]) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][22]  ( .D(n104137), 
        .CK(Clk), .RN(Rst), .Q(n73454) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][20]  ( .D(n104136), 
        .CK(Clk), .RN(n106418), .Q(n73603) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24567 ), .CK(Clk), .RN(Rst), .Q(n70034) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][19]  ( .D(n104135), 
        .CK(Clk), .RN(Rst), .Q(n73165) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24564 ), .CK(Clk), .RN(Rst), .Q(n72705) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][15]  ( .D(n104134), 
        .CK(Clk), .RN(Rst), .Q(n70769) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][13]  ( .D(n104133), 
        .CK(Clk), .RN(n106411), .Q(n71073) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][10]  ( .D(n104132), 
        .CK(Clk), .RN(n106376), .Q(n71222) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24555 ), .CK(Clk), .RN(n106449), .Q(n69631) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][1]  ( .D(n104138), 
        .CK(Clk), .RN(n106417), .Q(n71522) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24586 ), .CK(Clk), .RN(n106501), .Q(n70331) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24569 ), .CK(Clk), .RN(n106384), .Q(n70928) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[72][6]  ( .D(n104131), 
        .CK(Clk), .RN(Rst), .Q(n72264) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24768 ), .CK(Clk), .RN(Rst), .Q(n73885) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25130 ), .CK(Clk), .RN(n106445), .Q(n70314) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25128 ), .CK(Clk), .RN(Rst), .Q(n69509) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][27]  ( .D(
        \DLX_Datapath/RegisterFile/N25126 ), .CK(Clk), .RN(Rst), .Q(n74016) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][25]  ( .D(
        \DLX_Datapath/RegisterFile/N25124 ), .CK(Clk), .RN(n106428), .Q(n74157) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][10]  ( .D(
        \DLX_Datapath/RegisterFile/N25109 ), .CK(Clk), .RN(n106377), .Q(n71205) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][8]  ( .D(
        \DLX_Datapath/RegisterFile/N25107 ), .CK(Clk), .RN(Rst), .Q(n72398) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][6]  ( .D(
        \DLX_Datapath/RegisterFile/N25105 ), .CK(Clk), .RN(n106478), .Q(n72247) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][4]  ( .D(
        \DLX_Datapath/RegisterFile/N25103 ), .CK(Clk), .RN(n106411), .Q(n71952) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][2]  ( .D(
        \DLX_Datapath/RegisterFile/N25101 ), .CK(Clk), .RN(n106427), .Q(n71649) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][1]  ( .D(
        \DLX_Datapath/RegisterFile/N25100 ), .CK(Clk), .RN(n106419), .Q(n71505) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25129 ), .CK(Clk), .RN(Rst), .Q(n70456) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][28]  ( .D(
        \DLX_Datapath/RegisterFile/N25127 ), .CK(Clk), .RN(Rst), .Q(n70170) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25125 ), .CK(Clk), .RN(n106437), .Q(n70603) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][24]  ( .D(
        \DLX_Datapath/RegisterFile/N25123 ), .CK(Clk), .RN(n106408), .Q(n74297) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][23]  ( .D(
        \DLX_Datapath/RegisterFile/N25122 ), .CK(Clk), .RN(Rst), .Q(n73733) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25108 ), .CK(Clk), .RN(n106483), .Q(n72688) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25104 ), .CK(Clk), .RN(Rst), .Q(n72096) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][3]  ( .D(
        \DLX_Datapath/RegisterFile/N25102 ), .CK(Clk), .RN(n106380), .Q(n71354) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][0]  ( .D(
        \DLX_Datapath/RegisterFile/N25099 ), .CK(Clk), .RN(Rst), .Q(n69614) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][7]  ( .D(
        \DLX_Datapath/RegisterFile/N25106 ), .CK(Clk), .RN(n106401), .Q(n71798) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][22]  ( .D(
        \DLX_Datapath/RegisterFile/N25121 ), .CK(Clk), .RN(Rst), .Q(n73437) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][21]  ( .D(
        \DLX_Datapath/RegisterFile/N25120 ), .CK(Clk), .RN(Rst), .Q(n73874) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][20]  ( .D(
        \DLX_Datapath/RegisterFile/N25119 ), .CK(Clk), .RN(Rst), .Q(n73586) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][19]  ( .D(
        \DLX_Datapath/RegisterFile/N25118 ), .CK(Clk), .RN(Rst), .Q(n73148) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][18]  ( .D(
        \DLX_Datapath/RegisterFile/N25117 ), .CK(Clk), .RN(Rst), .Q(n73290) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][17]  ( .D(
        \DLX_Datapath/RegisterFile/N25116 ), .CK(Clk), .RN(n106506), .Q(n73006) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][16]  ( .D(
        \DLX_Datapath/RegisterFile/N25115 ), .CK(Clk), .RN(n106502), .Q(n72856) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][15]  ( .D(
        \DLX_Datapath/RegisterFile/N25114 ), .CK(Clk), .RN(Rst), .Q(n70752) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][14]  ( .D(
        \DLX_Datapath/RegisterFile/N25113 ), .CK(Clk), .RN(n106385), .Q(n70911) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][13]  ( .D(
        \DLX_Datapath/RegisterFile/N25112 ), .CK(Clk), .RN(Rst), .Q(n71056) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][12]  ( .D(
        \DLX_Datapath/RegisterFile/N25111 ), .CK(Clk), .RN(n106432), .Q(n70017) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[55][11]  ( .D(
        \DLX_Datapath/RegisterFile/N25110 ), .CK(Clk), .RN(n106464), .Q(n72546) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24093 ), .CK(Clk), .RN(Rst), .Q(n73322) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24091 ), .CK(Clk), .RN(Rst), .Q(n72888) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24089 ), .CK(Clk), .RN(Rst), .Q(n70943) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24087 ), .CK(Clk), .RN(Rst), .Q(n70049) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24085 ), .CK(Clk), .RN(Rst), .Q(n71237) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24083 ), .CK(Clk), .RN(Rst), .Q(n72430) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24081 ), .CK(Clk), .RN(Rst), .Q(n72279) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24079 ), .CK(Clk), .RN(n106409), .Q(n71984) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24077 ), .CK(Clk), .RN(n106425), .Q(n71681) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24076 ), .CK(Clk), .RN(Rst), .Q(n71537) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24106 ), .CK(Clk), .RN(Rst), .Q(n70346) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24105 ), .CK(Clk), .RN(Rst), .Q(n70488) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24104 ), .CK(Clk), .RN(n106495), .Q(n69541) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24103 ), .CK(Clk), .RN(Rst), .Q(n70202) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24102 ), .CK(Clk), .RN(Rst), .Q(n74048) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24101 ), .CK(Clk), .RN(n106444), .Q(n70635) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24100 ), .CK(Clk), .RN(Rst), .Q(n74189) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24099 ), .CK(Clk), .RN(Rst), .Q(n74329) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24098 ), .CK(Clk), .RN(Rst), .Q(n73765) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24097 ), .CK(Clk), .RN(n106395), .Q(n73469) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24096 ), .CK(Clk), .RN(n106454), .Q(n73906) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24095 ), .CK(Clk), .RN(Rst), .Q(n73618) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24094 ), .CK(Clk), .RN(n106492), .Q(n73180) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24092 ), .CK(Clk), .RN(Rst), .Q(n73038) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24090 ), .CK(Clk), .RN(n106386), .Q(n70784) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24088 ), .CK(Clk), .RN(Rst), .Q(n71088) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24086 ), .CK(Clk), .RN(Rst), .Q(n72578) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24084 ), .CK(Clk), .RN(Rst), .Q(n72720) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24082 ), .CK(Clk), .RN(n106399), .Q(n71830) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24080 ), .CK(Clk), .RN(n106440), .Q(n72128) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24078 ), .CK(Clk), .RN(n106378), .Q(n71386) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[87][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24075 ), .CK(Clk), .RN(Rst), .Q(n69646) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23272 ), .CK(Clk), .RN(n106435), .Q(n69567), .QN(n107271) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][28]  ( .D(
        \DLX_Datapath/RegisterFile/N23271 ), .CK(Clk), .RN(Rst), .Q(n70228), 
        .QN(n107808) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23274 ), .CK(Clk), .RN(n106437), .Q(n70372), .QN(n107904) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[113][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23273 ), .CK(Clk), .RN(n106443), .Q(n70514), .QN(n108000) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][25]  ( .D(
        \DLX_Datapath/RegisterFile/N23172 ), .CK(Clk), .RN(Rst), .Q(n74218) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][10]  ( .D(
        \DLX_Datapath/RegisterFile/N23157 ), .CK(Clk), .RN(n106373), .Q(n71266) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24769 ), .CK(Clk), .RN(n106440), .Q(n73448) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24767 ), .CK(Clk), .RN(n106460), .Q(n73597) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24764 ), .CK(Clk), .RN(n106506), .Q(n73017) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][31]  ( .D(
        \DLX_Datapath/RegisterFile/N23146 ), .CK(Clk), .RN(n106438), .Q(n70376) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][30]  ( .D(
        \DLX_Datapath/RegisterFile/N23145 ), .CK(Clk), .RN(n106442), .Q(n70518) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[117][29]  ( .D(
        \DLX_Datapath/RegisterFile/N23144 ), .CK(Clk), .RN(Rst), .Q(n69571) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][19]  ( .D(n104186), 
        .CK(Clk), .RN(Rst), .Q(n73159) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23158 ), .CK(Clk), .RN(Rst), .Q(n72607) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[19]  ( .D(n59085), .CK(Clk), .RN(n106430), 
        .Q(n61540), .QN(n107416) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][27]  ( .D(
        \DLX_Datapath/RegisterFile/N23174 ), .CK(Clk), .RN(n106474), .Q(n74077) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[116][26]  ( .D(
        \DLX_Datapath/RegisterFile/N23173 ), .CK(Clk), .RN(n106374), .Q(n70664) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24770 ), .CK(Clk), .RN(n106444), .Q(n73744) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[66][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24765 ), .CK(Clk), .RN(n106495), .Q(n73301) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25322 ), .CK(Clk), .RN(n106446), .Q(n70308), .QN(n107867) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][30]  ( .D(
        \DLX_Datapath/RegisterFile/N25321 ), .CK(Clk), .RN(n106431), .Q(n70450), .QN(n107964) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[49][29]  ( .D(
        \DLX_Datapath/RegisterFile/N25320 ), .CK(Clk), .RN(Rst), .Q(n69503), 
        .QN(n107227) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24746 ), .CK(Clk), .RN(Rst), .Q(n70326) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24745 ), .CK(Clk), .RN(n106424), .Q(n70468) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24744 ), .CK(Clk), .RN(Rst), .Q(n69521) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24743 ), .CK(Clk), .RN(n106494), .Q(n70182) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24742 ), .CK(Clk), .RN(n106476), .Q(n74028) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24741 ), .CK(Clk), .RN(Rst), .Q(n70615) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24740 ), .CK(Clk), .RN(Rst), .Q(n74169) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24739 ), .CK(Clk), .RN(n106455), .Q(n74309) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24738 ), .CK(Clk), .RN(n106383), .Q(n73745) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24737 ), .CK(Clk), .RN(n106481), .Q(n73449) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24736 ), .CK(Clk), .RN(n106387), .Q(n73886) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24735 ), .CK(Clk), .RN(n106385), .Q(n73598) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24734 ), .CK(Clk), .RN(Rst), .Q(n73160) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24733 ), .CK(Clk), .RN(n106495), .Q(n73302) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24732 ), .CK(Clk), .RN(Rst), .Q(n73018) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24731 ), .CK(Clk), .RN(n106501), .Q(n72868) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][15]  ( .D(
        \DLX_Datapath/RegisterFile/N24730 ), .CK(Clk), .RN(Rst), .Q(n70764) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][14]  ( .D(
        \DLX_Datapath/RegisterFile/N24729 ), .CK(Clk), .RN(n106384), .Q(n70923) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][13]  ( .D(
        \DLX_Datapath/RegisterFile/N24728 ), .CK(Clk), .RN(n106409), .Q(n71068) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24727 ), .CK(Clk), .RN(n106466), .Q(n70029) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24726 ), .CK(Clk), .RN(n106430), .Q(n72558) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][10]  ( .D(
        \DLX_Datapath/RegisterFile/N24725 ), .CK(Clk), .RN(n106376), .Q(n71217) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24724 ), .CK(Clk), .RN(Rst), .Q(n72700) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24723 ), .CK(Clk), .RN(Rst), .Q(n72410) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24722 ), .CK(Clk), .RN(n106400), .Q(n71810) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][6]  ( .D(
        \DLX_Datapath/RegisterFile/N24721 ), .CK(Clk), .RN(Rst), .Q(n72259) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24720 ), .CK(Clk), .RN(n106422), .Q(n72108) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24719 ), .CK(Clk), .RN(n106410), .Q(n71964) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24718 ), .CK(Clk), .RN(n106379), .Q(n71366) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24717 ), .CK(Clk), .RN(Rst), .Q(n71661) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24715 ), .CK(Clk), .RN(Rst), .Q(n69626) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[67][1]  ( .D(
        \DLX_Datapath/RegisterFile/N24716 ), .CK(Clk), .RN(n106418), .Q(n71517) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][31]  ( .D(
        \DLX_Datapath/RegisterFile/N24234 ), .CK(Clk), .RN(Rst), .Q(n70342) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24233 ), .CK(Clk), .RN(Rst), .Q(n70484) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24230 ), .CK(Clk), .RN(n106434), .Q(n74044) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[83][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24229 ), .CK(Clk), .RN(Rst), .Q(n70631) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][7]  ( .D(n103989), 
        .CK(Clk), .RN(Rst), .Q(n71878), .QN(n109055) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26564 ), .CK(Clk), .RN(n106478), .Q(
        n110841) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26570 ), .CK(Clk), .RN(Rst), .Q(n107938)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26569 ), .CK(Clk), .RN(Rst), .Q(n108034)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26566 ), .CK(Clk), .RN(n106473), .Q(
        n110738) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26565 ), .CK(Clk), .RN(Rst), .Q(n108143)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26563 ), .CK(Clk), .RN(Rst), .Q(n110942)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26568 ), .CK(Clk), .RN(Rst), .Q(n107180)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[10][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26567 ), .CK(Clk), .RN(n106448), .Q(
        n107843) );
  DFFR_X2 \DLX_ControlUnit/RMLcw2_reg[0]  ( .D(n60376), .CK(Clk), .RN(Rst), 
        .Q(n69340), .QN(n106957) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][0]  ( .D(
        \DLX_Datapath/RegisterFile/N22699 ), .CK(Clk), .RN(Rst), .Q(n69689) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][31]  ( .D(
        \DLX_Datapath/RegisterFile/N22570 ), .CK(Clk), .RN(n106371), .Q(n70394), .QN(n107921) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][30]  ( .D(
        \DLX_Datapath/RegisterFile/N22569 ), .CK(Clk), .RN(n106441), .Q(n70536), .QN(n108017) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][29]  ( .D(
        \DLX_Datapath/RegisterFile/N22568 ), .CK(Clk), .RN(Rst), .Q(n69589), 
        .QN(n107287) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][28]  ( .D(
        \DLX_Datapath/RegisterFile/N22567 ), .CK(Clk), .RN(Rst), .Q(n70250), 
        .QN(n107825) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][27]  ( .D(
        \DLX_Datapath/RegisterFile/N22566 ), .CK(Clk), .RN(Rst), .Q(n74096), 
        .QN(n110721) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][26]  ( .D(
        \DLX_Datapath/RegisterFile/N22565 ), .CK(Clk), .RN(Rst), .Q(n70683), 
        .QN(n108125) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[135][25]  ( .D(
        \DLX_Datapath/RegisterFile/N22564 ), .CK(Clk), .RN(Rst), .Q(n74237), 
        .QN(n110824) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][3]  ( .D(
        \DLX_Datapath/RegisterFile/N22702 ), .CK(Clk), .RN(Rst), .Q(n71429) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][21]  ( .D(
        \DLX_Datapath/RegisterFile/N26432 ), .CK(Clk), .RN(Rst), .Q(n110636)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][19]  ( .D(
        \DLX_Datapath/RegisterFile/N26430 ), .CK(Clk), .RN(Rst), .Q(n110103)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][9]  ( .D(
        \DLX_Datapath/RegisterFile/N26420 ), .CK(Clk), .RN(n106502), .Q(
        n109745) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][8]  ( .D(
        \DLX_Datapath/RegisterFile/N26419 ), .CK(Clk), .RN(Rst), .Q(n109530)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][6]  ( .D(
        \DLX_Datapath/RegisterFile/N26417 ), .CK(Clk), .RN(Rst), .Q(n109415)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[130][5]  ( .D(
        \DLX_Datapath/RegisterFile/N22704 ), .CK(Clk), .RN(n106458), .Q(n72171) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][10]  ( .D(n104004), 
        .CK(Clk), .RN(n106373), .Q(n71262) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][9]  ( .D(
        \DLX_Datapath/RegisterFile/N23284 ), .CK(Clk), .RN(Rst), .Q(n72745) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[112][11]  ( .D(
        \DLX_Datapath/RegisterFile/N23286 ), .CK(Clk), .RN(n106453), .Q(n72603) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][29]  ( .D(
        \DLX_Datapath/RegisterFile/N24200 ), .CK(Clk), .RN(Rst), .Q(n69538) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[9]  ( .D(n103929), .CK(Clk), .RN(n106467), 
        .Q(\DLX_ControlUnit/cw2 [9]) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[25]  ( .D(n59098), .CK(Clk), .RN(Rst), .Q(
        n100767), .QN(n107421) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][20]  ( .D(
        \DLX_Datapath/RegisterFile/N26431 ), .CK(Clk), .RN(n106451), .Q(
        n110425) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][16]  ( .D(
        \DLX_Datapath/RegisterFile/N26427 ), .CK(Clk), .RN(Rst), .Q(n109878)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][22]  ( .D(
        \DLX_Datapath/RegisterFile/N26433 ), .CK(Clk), .RN(n106389), .Q(
        n110316) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][18]  ( .D(
        \DLX_Datapath/RegisterFile/N26429 ), .CK(Clk), .RN(n106398), .Q(
        n110210) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][14]  ( .D(
        \DLX_Datapath/RegisterFile/N26425 ), .CK(Clk), .RN(n106472), .Q(
        n108375) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][12]  ( .D(
        \DLX_Datapath/RegisterFile/N26423 ), .CK(Clk), .RN(Rst), .Q(n107723)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][1]  ( .D(
        \DLX_Datapath/RegisterFile/N26412 ), .CK(Clk), .RN(n106426), .Q(
        n108839) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][13]  ( .D(
        \DLX_Datapath/RegisterFile/N26424 ), .CK(Clk), .RN(Rst), .Q(n108486)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][10]  ( .D(
        \DLX_Datapath/RegisterFile/N26421 ), .CK(Clk), .RN(Rst), .Q(n108600)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][23]  ( .D(
        \DLX_Datapath/RegisterFile/N26434 ), .CK(Clk), .RN(Rst), .Q(n110531)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][17]  ( .D(
        \DLX_Datapath/RegisterFile/N26428 ), .CK(Clk), .RN(Rst), .Q(n109995)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][15]  ( .D(
        \DLX_Datapath/RegisterFile/N26426 ), .CK(Clk), .RN(Rst), .Q(n108252)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][11]  ( .D(
        \DLX_Datapath/RegisterFile/N26422 ), .CK(Clk), .RN(Rst), .Q(n109638)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][5]  ( .D(
        \DLX_Datapath/RegisterFile/N26416 ), .CK(Clk), .RN(n106428), .Q(
        n109296) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][4]  ( .D(
        \DLX_Datapath/RegisterFile/N26415 ), .CK(Clk), .RN(Rst), .Q(n109188)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][3]  ( .D(
        \DLX_Datapath/RegisterFile/N26414 ), .CK(Clk), .RN(n106421), .Q(
        n108723) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][2]  ( .D(
        \DLX_Datapath/RegisterFile/N26413 ), .CK(Clk), .RN(n106423), .Q(
        n108951) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][0]  ( .D(
        \DLX_Datapath/RegisterFile/N26411 ), .CK(Clk), .RN(Rst), .Q(n107189)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[14][7]  ( .D(
        \DLX_Datapath/RegisterFile/N26418 ), .CK(Clk), .RN(Rst), .Q(n109068)
         );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][22]  ( .D(
        \DLX_Datapath/RegisterFile/N24193 ), .CK(Clk), .RN(Rst), .Q(n73466) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][12]  ( .D(
        \DLX_Datapath/RegisterFile/N24183 ), .CK(Clk), .RN(Rst), .Q(n70046) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][9]  ( .D(
        \DLX_Datapath/RegisterFile/N24180 ), .CK(Clk), .RN(Rst), .Q(n72717) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][17]  ( .D(
        \DLX_Datapath/RegisterFile/N24188 ), .CK(Clk), .RN(n106493), .Q(n73035) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][25]  ( .D(
        \DLX_Datapath/RegisterFile/N24196 ), .CK(Clk), .RN(n106390), .Q(n74186) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][23]  ( .D(
        \DLX_Datapath/RegisterFile/N24194 ), .CK(Clk), .RN(Rst), .Q(n73762) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][6]  ( .D(n104098), 
        .CK(Clk), .RN(Rst), .Q(n72276) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][31]  ( .D(n104105), 
        .CK(Clk), .RN(Rst), .Q(n70343) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][14]  ( .D(n104099), 
        .CK(Clk), .RN(n106390), .Q(n70940) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][28]  ( .D(
        \DLX_Datapath/RegisterFile/N24199 ), .CK(Clk), .RN(Rst), .Q(n70199) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][15]  ( .D(n104108), 
        .CK(Clk), .RN(n106385), .Q(n70781) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][10]  ( .D(n104104), 
        .CK(Clk), .RN(Rst), .Q(n71234) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][20]  ( .D(
        \DLX_Datapath/RegisterFile/N24191 ), .CK(Clk), .RN(Rst), .Q(n73615) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][19]  ( .D(
        \DLX_Datapath/RegisterFile/N24190 ), .CK(Clk), .RN(n106492), .Q(n73177) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][27]  ( .D(
        \DLX_Datapath/RegisterFile/N24198 ), .CK(Clk), .RN(Rst), .Q(n74045) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][13]  ( .D(n104106), 
        .CK(Clk), .RN(Rst), .Q(n71085) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][0]  ( .D(
        \DLX_Datapath/RegisterFile/N24171 ), .CK(Clk), .RN(Rst), .Q(n69643) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][1]  ( .D(n104107), 
        .CK(Clk), .RN(Rst), .Q(n71534) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][30]  ( .D(
        \DLX_Datapath/RegisterFile/N26121 ), .CK(Clk), .RN(n106440), .Q(n70544) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][26]  ( .D(
        \DLX_Datapath/RegisterFile/N26117 ), .CK(Clk), .RN(Rst), .Q(n70691), 
        .QN(n108132) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][24]  ( .D(
        \DLX_Datapath/RegisterFile/N26115 ), .CK(Clk), .RN(n106423), .Q(n74385) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][29]  ( .D(
        \DLX_Datapath/RegisterFile/N26120 ), .CK(Clk), .RN(n106433), .Q(n69469) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][31]  ( .D(
        \DLX_Datapath/RegisterFile/N26122 ), .CK(Clk), .RN(Rst), .Q(n70402) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][28]  ( .D(
        \DLX_Datapath/RegisterFile/N26119 ), .CK(Clk), .RN(n106504), .Q(n70258), .QN(n107832) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][27]  ( .D(
        \DLX_Datapath/RegisterFile/N26118 ), .CK(Clk), .RN(Rst), .Q(n74104) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[24][25]  ( .D(
        \DLX_Datapath/RegisterFile/N26116 ), .CK(Clk), .RN(Rst), .Q(n74245) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[27]  ( .D(n103932), .CK(Clk), .RN(Rst), 
        .Q(n62198) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[25]  ( .D(n103948), .CK(Clk), .RN(Rst), 
        .Q(net2411291) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[26]  ( .D(n103953), .CK(Clk), .RN(Rst), 
        .Q(n66263) );
  DFFR_X2 \DLX_Datapath/TA_IFID_reg[24]  ( .D(n103943), .CK(Clk), .RN(Rst), 
        .Q(n62197) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][7]  ( .D(
        \DLX_Datapath/RegisterFile/N24178 ), .CK(Clk), .RN(Rst), .Q(n71827) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][3]  ( .D(
        \DLX_Datapath/RegisterFile/N24174 ), .CK(Clk), .RN(n106378), .Q(n71383) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][26]  ( .D(
        \DLX_Datapath/RegisterFile/N24197 ), .CK(Clk), .RN(n106444), .Q(n70632) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][21]  ( .D(
        \DLX_Datapath/RegisterFile/N24192 ), .CK(Clk), .RN(n106454), .Q(n73903) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][18]  ( .D(
        \DLX_Datapath/RegisterFile/N24189 ), .CK(Clk), .RN(Rst), .Q(n73319) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][16]  ( .D(
        \DLX_Datapath/RegisterFile/N24187 ), .CK(Clk), .RN(Rst), .Q(n72885) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][11]  ( .D(
        \DLX_Datapath/RegisterFile/N24182 ), .CK(Clk), .RN(Rst), .Q(n72575) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][8]  ( .D(
        \DLX_Datapath/RegisterFile/N24179 ), .CK(Clk), .RN(Rst), .Q(n72427) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][30]  ( .D(
        \DLX_Datapath/RegisterFile/N24201 ), .CK(Clk), .RN(n106424), .Q(n70485) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][5]  ( .D(
        \DLX_Datapath/RegisterFile/N24176 ), .CK(Clk), .RN(Rst), .Q(n72125) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][4]  ( .D(
        \DLX_Datapath/RegisterFile/N24175 ), .CK(Clk), .RN(n106409), .Q(n71981) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][2]  ( .D(
        \DLX_Datapath/RegisterFile/N24173 ), .CK(Clk), .RN(n106426), .Q(n71678) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[84][24]  ( .D(
        \DLX_Datapath/RegisterFile/N24195 ), .CK(Clk), .RN(Rst), .Q(n74326) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][31]  ( .D(
        \DLX_Datapath/RegisterFile/N25898 ), .CK(Clk), .RN(Rst), .Q(n70395) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][26]  ( .D(
        \DLX_Datapath/RegisterFile/N25893 ), .CK(Clk), .RN(Rst), .Q(n70684) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][9]  ( .D(
        \DLX_Datapath/RegisterFile/N25876 ), .CK(Clk), .RN(n106504), .Q(n72769) );
  DFFR_X2 \DLX_Datapath/RegisterFile/phy_regfile_reg[31][5]  ( .D(
        \DLX_Datapath/RegisterFile/N25872 ), .CK(Clk), .RN(n106455), .Q(n72177) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[22]  ( .D(n106574), .CK(Clk), .RN(Rst), .Q(
        n69765) );
  DFFR_X2 \DLX_Datapath/IR_IFID_reg[31]  ( .D(n106559), .CK(Clk), .RN(Rst), 
        .Q(n69381), .QN(n107149) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[6]  ( .D(n106581), .CK(Clk), .RN(n106468), 
        .Q(\DLX_ControlUnit/cw2 [6]) );
  DFFR_X2 \DLX_ControlUnit/cw2_reg[2]  ( .D(n106580), .CK(Clk), .RN(n106468), 
        .Q(\DLX_ControlUnit/cw2 [2]) );
  NAND2_X1 U90527 ( .A1(n69430), .A2(n105871), .ZN(n84077) );
  NAND2_X1 U90528 ( .A1(n71613), .A2(n83145), .ZN(n84039) );
  NAND2_X1 U90529 ( .A1(n83145), .A2(n71757), .ZN(n84010) );
  NAND2_X1 U90530 ( .A1(n71462), .A2(n83145), .ZN(n83981) );
  NAND2_X1 U90531 ( .A1(n72060), .A2(n83145), .ZN(n83952) );
  NAND2_X1 U90532 ( .A1(n72204), .A2(n83145), .ZN(n83923) );
  NAND2_X1 U90533 ( .A1(n71906), .A2(n83145), .ZN(n83865) );
  NAND2_X1 U90534 ( .A1(n72506), .A2(n83145), .ZN(n83836) );
  NAND2_X1 U90535 ( .A1(n83145), .A2(n72796), .ZN(n83807) );
  NAND2_X1 U90536 ( .A1(n72654), .A2(n83145), .ZN(n83748) );
  NAND2_X1 U90537 ( .A1(n70125), .A2(n105871), .ZN(n83719) );
  NAND2_X1 U90538 ( .A1(n71164), .A2(n105871), .ZN(n83690) );
  NAND2_X1 U90539 ( .A1(n71019), .A2(n105871), .ZN(n83661) );
  NAND2_X1 U90540 ( .A1(n70860), .A2(n105871), .ZN(n83632) );
  NAND2_X1 U90541 ( .A1(n72964), .A2(n105871), .ZN(n83603) );
  NAND2_X1 U90542 ( .A1(n73114), .A2(n105871), .ZN(n83574) );
  NAND2_X1 U90543 ( .A1(n73398), .A2(n105871), .ZN(n83545) );
  NAND2_X1 U90544 ( .A1(n73256), .A2(n105871), .ZN(n83516) );
  NAND2_X1 U90545 ( .A1(n73694), .A2(n105871), .ZN(n83487) );
  NAND2_X1 U90546 ( .A1(n73982), .A2(n105871), .ZN(n83458) );
  NAND2_X1 U90547 ( .A1(n73545), .A2(n105871), .ZN(n83429) );
  NAND2_X1 U90548 ( .A1(n73841), .A2(n105871), .ZN(n83400) );
  NAND2_X1 U90549 ( .A1(n74405), .A2(n105871), .ZN(n83371) );
  NAND2_X1 U90550 ( .A1(n74265), .A2(n105871), .ZN(n83342) );
  NAND2_X1 U90551 ( .A1(n70711), .A2(n105871), .ZN(n83313) );
  NAND2_X1 U90552 ( .A1(n74124), .A2(n105871), .ZN(n83283) );
  NAND2_X1 U90553 ( .A1(n70278), .A2(n105871), .ZN(n83251) );
  NAND2_X1 U90554 ( .A1(n69429), .A2(n105871), .ZN(n83219) );
  NAND2_X1 U90555 ( .A1(n70564), .A2(n105871), .ZN(n83190) );
  NAND2_X1 U90556 ( .A1(n70422), .A2(n105871), .ZN(n83144) );
  NAND2_X1 U90557 ( .A1(n71313), .A2(n83145), .ZN(n83778) );
  NAND2_X1 U90558 ( .A1(n83145), .A2(n72355), .ZN(n83894) );
  CLKBUF_X3 U90559 ( .A(n80041), .Z(n105151) );
  CLKBUF_X3 U90560 ( .A(n107022), .Z(n105199) );
  CLKBUF_X1 U90561 ( .A(n82142), .Z(n104893) );
  CLKBUF_X1 U90562 ( .A(n105013), .Z(n105155) );
  NAND2_X1 U90563 ( .A1(n99672), .A2(n99673), .ZN(n104377) );
  INV_X1 U90564 ( .A(n104377), .ZN(n99616) );
  NOR4_X1 U90565 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [3]), 
        .A2(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [2]), .A3(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [1]), .A4(n104913), 
        .ZN(n104378) );
  INV_X1 U90566 ( .A(n104378), .ZN(n104798) );
  NOR2_X1 U90567 ( .A1(n107128), .A2(n98369), .ZN(n94555) );
  NOR3_X1 U90568 ( .A1(n104923), .A2(n94848), .A3(n94553), .ZN(n94814) );
  NAND2_X1 U90569 ( .A1(n83162), .A2(n71144), .ZN(n104379) );
  INV_X1 U90570 ( .A(n104379), .ZN(n83671) );
  NAND2_X1 U90571 ( .A1(n99751), .A2(n99752), .ZN(n104380) );
  INV_X1 U90572 ( .A(n104380), .ZN(n99728) );
  OAI21_X1 U90573 ( .B1(n104783), .B2(n104913), .A(n82302), .ZN(n104804) );
  NOR4_X1 U90574 ( .A1(n105062), .A2(n104390), .A3(n104833), .A4(n62204), .ZN(
        n104381) );
  INV_X1 U90575 ( .A(n104381), .ZN(n105086) );
  NAND2_X1 U90576 ( .A1(n104785), .A2(n82287), .ZN(n104382) );
  INV_X1 U90577 ( .A(n104382), .ZN(n82027) );
  NOR2_X1 U90578 ( .A1(n96267), .A2(n106757), .ZN(n105426) );
  NAND2_X1 U90579 ( .A1(n83162), .A2(n70840), .ZN(n104383) );
  INV_X1 U90580 ( .A(n104383), .ZN(n83613) );
  NOR2_X1 U90581 ( .A1(n94661), .A2(n94553), .ZN(n105604) );
  NOR2_X1 U90582 ( .A1(n96416), .A2(n96417), .ZN(n105924) );
  NOR2_X1 U90583 ( .A1(n96293), .A2(n96294), .ZN(n105931) );
  NOR2_X1 U90584 ( .A1(n96166), .A2(n96167), .ZN(n105436) );
  NAND2_X1 U90585 ( .A1(n104743), .A2(n104494), .ZN(n104384) );
  INV_X1 U90586 ( .A(n104384), .ZN(n82324) );
  NAND2_X1 U90587 ( .A1(n100047), .A2(n100048), .ZN(n104385) );
  INV_X1 U90588 ( .A(n104385), .ZN(n100022) );
  AOI22_X1 U90589 ( .A1(n82260), .A2(n104918), .B1(n105153), .B2(n82329), .ZN(
        n82298) );
  NAND2_X1 U90590 ( .A1(n104729), .A2(n104785), .ZN(n104386) );
  INV_X1 U90591 ( .A(n104386), .ZN(n104919) );
  NOR2_X1 U90592 ( .A1(n96267), .A2(n106757), .ZN(n105427) );
  NAND2_X1 U90593 ( .A1(n83162), .A2(n73094), .ZN(n104387) );
  INV_X1 U90594 ( .A(n104387), .ZN(n83555) );
  NOR2_X1 U90595 ( .A1(n94661), .A2(n94553), .ZN(n105603) );
  NOR2_X1 U90596 ( .A1(n96293), .A2(n96354), .ZN(n105977) );
  NOR2_X1 U90597 ( .A1(n95169), .A2(n106748), .ZN(n105534) );
  NOR2_X1 U90598 ( .A1(n96416), .A2(n96486), .ZN(n105987) );
  NOR2_X1 U90599 ( .A1(n95725), .A2(n95726), .ZN(n105483) );
  NOR2_X1 U90600 ( .A1(n96166), .A2(n96231), .ZN(n105995) );
  AOI21_X1 U90601 ( .B1(n111159), .B2(net2465244), .A(n82075), .ZN(n82431) );
  NOR3_X1 U90602 ( .A1(n106697), .A2(n105056), .A3(n104582), .ZN(n81210) );
  NAND2_X1 U90603 ( .A1(n99811), .A2(n99812), .ZN(n104388) );
  INV_X1 U90604 ( .A(n104388), .ZN(n99747) );
  NAND2_X1 U90605 ( .A1(n99467), .A2(n99468), .ZN(n104389) );
  INV_X1 U90606 ( .A(n104389), .ZN(n99091) );
  NAND4_X2 U90607 ( .A1(n104831), .A2(n104832), .A3(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [0]), .A4(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [3]), .ZN(n104390) );
  INV_X1 U90608 ( .A(n104390), .ZN(n82465) );
  NAND2_X1 U90609 ( .A1(n99878), .A2(n99879), .ZN(n104391) );
  INV_X1 U90610 ( .A(n104391), .ZN(n99870) );
  NAND2_X1 U90611 ( .A1(n104918), .A2(n104804), .ZN(n104392) );
  INV_X1 U90612 ( .A(n104392), .ZN(n105018) );
  NOR2_X1 U90613 ( .A1(n96267), .A2(n106757), .ZN(n105428) );
  NAND2_X1 U90614 ( .A1(n83162), .A2(n73236), .ZN(n104393) );
  INV_X1 U90615 ( .A(n104393), .ZN(n83497) );
  NOR2_X1 U90616 ( .A1(n95448), .A2(n95449), .ZN(n104928) );
  NOR2_X1 U90617 ( .A1(n95488), .A2(n95516), .ZN(n104929) );
  AOI21_X1 U90618 ( .B1(n96010), .B2(n94554), .A(n96294), .ZN(n105934) );
  NOR2_X1 U90619 ( .A1(n94623), .A2(n94553), .ZN(n105613) );
  NOR2_X1 U90620 ( .A1(n95037), .A2(n106748), .ZN(n105555) );
  NOR2_X1 U90621 ( .A1(n96416), .A2(n96486), .ZN(n105988) );
  NOR2_X1 U90622 ( .A1(n96293), .A2(n96354), .ZN(n105978) );
  NOR2_X1 U90623 ( .A1(n96166), .A2(n96203), .ZN(n104975) );
  NOR2_X1 U90624 ( .A1(n95725), .A2(n95799), .ZN(n104936) );
  OAI21_X1 U90625 ( .B1(n62185), .B2(n104753), .A(n82170), .ZN(n82169) );
  AOI22_X1 U90626 ( .A1(n79809), .A2(\DLX_Datapath/ArithLogUnit/A_log [20]), 
        .B1(n104394), .B2(\DLX_Datapath/ArithLogUnit/B_log [20]), .ZN(n79808)
         );
  INV_X1 U90627 ( .A(n79811), .ZN(n104394) );
  NAND2_X1 U90628 ( .A1(n99626), .A2(n99627), .ZN(n104395) );
  INV_X1 U90629 ( .A(n104395), .ZN(n99583) );
  NOR2_X1 U90630 ( .A1(n82200), .A2(n105021), .ZN(n104896) );
  NOR3_X1 U90631 ( .A1(n62190), .A2(n105056), .A3(n106697), .ZN(n104396) );
  INV_X1 U90632 ( .A(n104396), .ZN(n81207) );
  OR2_X1 U90633 ( .A1(IR_in[11]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [3]), .ZN(n104414) );
  NAND2_X1 U90634 ( .A1(n82707), .A2(n82659), .ZN(n104894) );
  NOR4_X1 U90635 ( .A1(n95412), .A2(n111056), .A3(n94894), .A4(n94895), .ZN(
        n95170) );
  NAND2_X1 U90636 ( .A1(n99691), .A2(n99692), .ZN(n104397) );
  INV_X1 U90637 ( .A(n104397), .ZN(n99151) );
  NOR3_X1 U90638 ( .A1(n95911), .A2(n94848), .A3(n95517), .ZN(n95878) );
  AOI21_X1 U90639 ( .B1(n82271), .B2(n82272), .A(n105018), .ZN(n82297) );
  NOR2_X1 U90640 ( .A1(n105152), .A2(n104713), .ZN(n105050) );
  AOI21_X1 U90641 ( .B1(n96560), .B2(n94554), .A(n96800), .ZN(n106033) );
  NAND2_X1 U90642 ( .A1(n83162), .A2(n73962), .ZN(n104398) );
  INV_X1 U90643 ( .A(n104398), .ZN(n83439) );
  NAND2_X1 U90644 ( .A1(n100058), .A2(n100059), .ZN(n104399) );
  INV_X1 U90645 ( .A(n104399), .ZN(n99233) );
  NOR2_X1 U90646 ( .A1(n96127), .A2(n106757), .ZN(n105439) );
  NOR2_X1 U90647 ( .A1(n96204), .A2(n96231), .ZN(n105998) );
  NOR2_X1 U90648 ( .A1(n95448), .A2(n95516), .ZN(n105973) );
  NOR2_X1 U90649 ( .A1(n96331), .A2(n96354), .ZN(n105980) );
  NOR2_X1 U90650 ( .A1(n97710), .A2(n97780), .ZN(n106127) );
  NOR2_X1 U90651 ( .A1(n94770), .A2(n94553), .ZN(n105594) );
  NOR2_X1 U90652 ( .A1(n95169), .A2(n106748), .ZN(n105533) );
  NOR2_X1 U90653 ( .A1(n98004), .A2(n98005), .ZN(n105286) );
  NOR2_X1 U90654 ( .A1(n96933), .A2(n104697), .ZN(n104876) );
  NOR2_X1 U90655 ( .A1(n96454), .A2(n96486), .ZN(n105984) );
  NOR2_X1 U90656 ( .A1(n96416), .A2(n96453), .ZN(n104933) );
  AOI21_X1 U90657 ( .B1(n96010), .B2(n94771), .A(n96417), .ZN(n105926) );
  NOR2_X1 U90658 ( .A1(n96293), .A2(n96330), .ZN(n104960) );
  NOR2_X1 U90659 ( .A1(n96166), .A2(n96167), .ZN(n105434) );
  NOR2_X1 U90660 ( .A1(n95799), .A2(n95763), .ZN(n105476) );
  NOR2_X1 U90661 ( .A1(n95725), .A2(n95726), .ZN(n105481) );
  NOR2_X1 U90662 ( .A1(n97967), .A2(n98024), .ZN(n106087) );
  NOR3_X1 U90663 ( .A1(n104400), .A2(IR_in[2]), .A3(n81960), .ZN(n81958) );
  INV_X1 U90664 ( .A(n81998), .ZN(n104400) );
  NAND4_X2 U90665 ( .A1(n82185), .A2(n104868), .A3(n82183), .A4(n82184), .ZN(
        n60303) );
  AOI22_X1 U90666 ( .A1(n79842), .A2(\DLX_Datapath/ArithLogUnit/A_log [16]), 
        .B1(n104401), .B2(\DLX_Datapath/ArithLogUnit/B_log [16]), .ZN(n79841)
         );
  INV_X1 U90667 ( .A(n79844), .ZN(n104401) );
  NAND2_X1 U90668 ( .A1(n82412), .A2(n108275), .ZN(n104402) );
  INV_X1 U90669 ( .A(n104402), .ZN(n82320) );
  AOI22_X1 U90670 ( .A1(IR_in[10]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [2]), .B1(IR_in[9]), 
        .B2(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [1]), .ZN(n104403)
         );
  INV_X1 U90671 ( .A(n104403), .ZN(n104748) );
  NAND3_X2 U90672 ( .A1(n59435), .A2(n90271), .A3(n59443), .ZN(n90161) );
  NOR3_X1 U90673 ( .A1(n62190), .A2(n105055), .A3(n106697), .ZN(n104404) );
  INV_X1 U90674 ( .A(n104404), .ZN(n86190) );
  XOR2_X1 U90675 ( .A(n107027), .B(n95131), .Z(n86220) );
  NAND2_X1 U90676 ( .A1(n106771), .A2(n82281), .ZN(n82664) );
  NAND2_X1 U90677 ( .A1(n99931), .A2(n99932), .ZN(n104405) );
  INV_X1 U90678 ( .A(n104405), .ZN(n99907) );
  NAND2_X1 U90679 ( .A1(n99922), .A2(\DLX_Datapath/ArithLogUnit/B_mul [13]), 
        .ZN(n104406) );
  INV_X1 U90680 ( .A(n104406), .ZN(n99037) );
  AOI22_X1 U90681 ( .A1(n82302), .A2(n104913), .B1(n104407), .B2(n104408), 
        .ZN(n82260) );
  INV_X1 U90682 ( .A(n104773), .ZN(n104407) );
  INV_X1 U90683 ( .A(n104760), .ZN(n104408) );
  XOR2_X1 U90684 ( .A(n82217), .B(n105153), .Z(n82220) );
  AOI21_X1 U90685 ( .B1(n96560), .B2(n94554), .A(n96800), .ZN(n106034) );
  NAND2_X1 U90686 ( .A1(n86300), .A2(n81888), .ZN(n104409) );
  INV_X1 U90687 ( .A(n104409), .ZN(n86299) );
  NAND2_X1 U90688 ( .A1(n83162), .A2(n73525), .ZN(n104410) );
  INV_X1 U90689 ( .A(n104410), .ZN(n83410) );
  NAND2_X1 U90690 ( .A1(n100107), .A2(n100108), .ZN(n104411) );
  INV_X1 U90691 ( .A(n104411), .ZN(n99251) );
  NOR2_X1 U90692 ( .A1(n96527), .A2(n106757), .ZN(n105411) );
  NOR2_X1 U90693 ( .A1(n96088), .A2(n96013), .ZN(n104767) );
  NOR2_X1 U90694 ( .A1(n95762), .A2(n95763), .ZN(n104958) );
  NOR2_X1 U90695 ( .A1(n95448), .A2(n95516), .ZN(n105975) );
  NOR2_X1 U90696 ( .A1(n97967), .A2(n98004), .ZN(n105283) );
  NOR2_X1 U90697 ( .A1(n97710), .A2(n97711), .ZN(n105320) );
  NOR2_X1 U90698 ( .A1(n97574), .A2(n97673), .ZN(n105330) );
  NOR2_X1 U90699 ( .A1(n96969), .A2(n96970), .ZN(n105376) );
  NOR2_X1 U90700 ( .A1(n96910), .A2(n96837), .ZN(n105380) );
  NOR2_X1 U90701 ( .A1(n96454), .A2(n96453), .ZN(n105414) );
  NOR2_X1 U90702 ( .A1(n96331), .A2(n96330), .ZN(n105422) );
  NOR2_X1 U90703 ( .A1(n96293), .A2(n96294), .ZN(n105932) );
  NOR2_X1 U90704 ( .A1(n96204), .A2(n96203), .ZN(n105430) );
  NOR2_X1 U90705 ( .A1(n98005), .A2(n98024), .ZN(n106089) );
  NOR2_X1 U90706 ( .A1(n96933), .A2(n97031), .ZN(n104859) );
  NOR2_X1 U90707 ( .A1(n96416), .A2(n96417), .ZN(n105925) );
  NOR2_X1 U90708 ( .A1(n96166), .A2(n96231), .ZN(n105997) );
  NOR2_X1 U90709 ( .A1(n95725), .A2(n95799), .ZN(n104937) );
  NOR2_X1 U90710 ( .A1(n95410), .A2(n106748), .ZN(n104952) );
  NOR2_X1 U90711 ( .A1(n94770), .A2(n94553), .ZN(n105592) );
  OR2_X1 U90712 ( .A1(n105152), .A2(IR_in[4]), .ZN(n104422) );
  XOR2_X1 U90713 ( .A(n99012), .B(n81812), .Z(n81811) );
  AOI22_X1 U90714 ( .A1(n79908), .A2(\DLX_Datapath/ArithLogUnit/A_log [8]), 
        .B1(n104412), .B2(\DLX_Datapath/ArithLogUnit/B_log [8]), .ZN(n79907)
         );
  INV_X1 U90715 ( .A(n79910), .ZN(n104412) );
  OAI21_X1 U90716 ( .B1(net2465244), .B2(n104753), .A(n82040), .ZN(n82039) );
  NAND2_X1 U90717 ( .A1(n99766), .A2(n99767), .ZN(n104413) );
  INV_X1 U90718 ( .A(n104413), .ZN(n99707) );
  AOI21_X1 U90719 ( .B1(n69326), .B2(n59415), .A(\DLX_Datapath/IR_IDEX[29] ), 
        .ZN(n100338) );
  AOI21_X1 U90720 ( .B1(n105036), .B2(n105037), .A(n104774), .ZN(n105035) );
  NOR3_X1 U90721 ( .A1(n106697), .A2(n105058), .A3(n104582), .ZN(n85183) );
  OAI21_X1 U90722 ( .B1(n104752), .B2(n104750), .A(n104414), .ZN(n104743) );
  XOR2_X1 U90723 ( .A(n99973), .B(n99946), .Z(n99936) );
  NAND2_X1 U90724 ( .A1(n99886), .A2(n99887), .ZN(n104415) );
  INV_X1 U90725 ( .A(n104415), .ZN(n99860) );
  NAND3_X2 U90726 ( .A1(n107139), .A2(n59435), .A3(n90134), .ZN(n90153) );
  NOR3_X1 U90727 ( .A1(n62199), .A2(n62194), .A3(n104494), .ZN(n104832) );
  NAND2_X1 U90728 ( .A1(n99595), .A2(n99596), .ZN(n104416) );
  INV_X1 U90729 ( .A(n104416), .ZN(n99533) );
  NAND2_X1 U90730 ( .A1(n99375), .A2(n99376), .ZN(n104417) );
  INV_X1 U90731 ( .A(n104417), .ZN(n99051) );
  OAI21_X1 U90732 ( .B1(n57430), .B2(n105153), .A(n110963), .ZN(n105082) );
  OAI21_X1 U90733 ( .B1(n111130), .B2(n104920), .A(net113153), .ZN(n106345) );
  NAND2_X1 U90734 ( .A1(n104708), .A2(n105014), .ZN(n104418) );
  INV_X1 U90735 ( .A(n104418), .ZN(n82022) );
  NOR2_X1 U90736 ( .A1(n97449), .A2(n97547), .ZN(n105343) );
  NOR2_X1 U90737 ( .A1(n106328), .A2(n105204), .ZN(n81889) );
  NAND2_X1 U90738 ( .A1(n83114), .A2(n74206), .ZN(n104419) );
  INV_X1 U90739 ( .A(n104419), .ZN(n83325) );
  NOR3_X1 U90740 ( .A1(\dp_cluster_2/DLX_Datapath/RegisterFile/N27633 ), .A2(
        n86222), .A3(n86228), .ZN(n83259) );
  OAI21_X1 U90741 ( .B1(n104420), .B2(n99624), .A(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .ZN(n99279) );
  INV_X1 U90742 ( .A(n100146), .ZN(n104420) );
  NOR3_X1 U90743 ( .A1(n69800), .A2(n69330), .A3(n99001), .ZN(n104421) );
  INV_X1 U90744 ( .A(n104421), .ZN(n98980) );
  NOR2_X1 U90745 ( .A1(n97840), .A2(n97895), .ZN(n106118) );
  XOR2_X1 U90746 ( .A(n82487), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [2]), .Z(n106815) );
  NOR2_X1 U90747 ( .A1(n96204), .A2(n96231), .ZN(n106000) );
  NOR2_X1 U90748 ( .A1(n104847), .A2(n96052), .ZN(n104890) );
  NOR2_X1 U90749 ( .A1(n96050), .A2(n96013), .ZN(n105447) );
  NOR2_X1 U90750 ( .A1(n95725), .A2(n95762), .ZN(n104949) );
  NOR2_X1 U90751 ( .A1(n95488), .A2(n95489), .ZN(n104979) );
  NOR2_X1 U90752 ( .A1(n95448), .A2(n95449), .ZN(n104927) );
  NOR2_X1 U90753 ( .A1(n96837), .A2(n96874), .ZN(n105386) );
  NOR2_X1 U90754 ( .A1(n96527), .A2(n106757), .ZN(n105410) );
  NOR2_X1 U90755 ( .A1(n95989), .A2(n95555), .ZN(n105451) );
  NOR2_X1 U90756 ( .A1(n95912), .A2(n104822), .ZN(n105464) );
  AOI21_X1 U90757 ( .B1(n95450), .B2(n94554), .A(n95726), .ZN(n104970) );
  NOR2_X1 U90758 ( .A1(n98004), .A2(n98005), .ZN(n105287) );
  NOR2_X1 U90759 ( .A1(n97710), .A2(n97711), .ZN(n105321) );
  NOR2_X1 U90760 ( .A1(n97574), .A2(n97673), .ZN(n105331) );
  NOR2_X1 U90761 ( .A1(n96969), .A2(n96970), .ZN(n105375) );
  NOR2_X1 U90762 ( .A1(n96933), .A2(n104697), .ZN(n104877) );
  NOR2_X1 U90763 ( .A1(n96454), .A2(n96486), .ZN(n105986) );
  NOR2_X1 U90764 ( .A1(n96416), .A2(n96453), .ZN(n104934) );
  AOI21_X1 U90765 ( .B1(n96010), .B2(n94771), .A(n96417), .ZN(n105928) );
  NOR2_X1 U90766 ( .A1(n96331), .A2(n96354), .ZN(n105982) );
  NOR2_X1 U90767 ( .A1(n96293), .A2(n96330), .ZN(n104961) );
  NOR2_X1 U90768 ( .A1(n96166), .A2(n96203), .ZN(n104976) );
  NOR2_X1 U90769 ( .A1(n95799), .A2(n95763), .ZN(n105477) );
  NOR2_X1 U90770 ( .A1(n97967), .A2(n98060), .ZN(n105280) );
  NOR2_X1 U90771 ( .A1(n95300), .A2(n106748), .ZN(n104999) );
  NOR2_X1 U90772 ( .A1(n94770), .A2(n94553), .ZN(n105593) );
  NOR4_X1 U90773 ( .A1(n104422), .A2(n104423), .A3(IR_in[1]), .A4(n82636), 
        .ZN(n81980) );
  INV_X1 U90774 ( .A(n81998), .ZN(n104423) );
  XOR2_X1 U90775 ( .A(n99058), .B(n99388), .Z(n99387) );
  AOI22_X1 U90776 ( .A1(n79941), .A2(\DLX_Datapath/ArithLogUnit/A_log [4]), 
        .B1(n104424), .B2(\DLX_Datapath/ArithLogUnit/B_log [4]), .ZN(n79940)
         );
  INV_X1 U90777 ( .A(n79943), .ZN(n104424) );
  OAI21_X1 U90778 ( .B1(n57425), .B2(n104753), .A(n82145), .ZN(n82144) );
  NAND3_X2 U90779 ( .A1(n81221), .A2(n106280), .A3(n81232), .ZN(n81235) );
  NOR3_X1 U90780 ( .A1(n106697), .A2(n62190), .A3(n105058), .ZN(n85180) );
  XOR2_X1 U90781 ( .A(n99938), .B(n99901), .Z(n99891) );
  AOI21_X1 U90782 ( .B1(n64246), .B2(n64247), .A(n100278), .ZN(n100399) );
  AOI22_X1 U90783 ( .A1(n98944), .A2(n107129), .B1(n105036), .B2(n105037), 
        .ZN(n104814) );
  OAI21_X1 U90784 ( .B1(n104895), .B2(n104896), .A(n82302), .ZN(n104773) );
  OAI21_X1 U90785 ( .B1(n105041), .B2(n82290), .A(n82661), .ZN(n104465) );
  NAND3_X2 U90786 ( .A1(n59435), .A2(n107139), .A3(n90271), .ZN(n90171) );
  NAND2_X1 U90787 ( .A1(n99817), .A2(n99818), .ZN(n104425) );
  INV_X1 U90788 ( .A(n104425), .ZN(n99777) );
  NAND2_X1 U90789 ( .A1(n99966), .A2(n99967), .ZN(n104426) );
  INV_X1 U90790 ( .A(n104426), .ZN(n99952) );
  OAI21_X1 U90791 ( .B1(n100233), .B2(n104427), .A(n104428), .ZN(n104446) );
  INV_X1 U90792 ( .A(n100232), .ZN(n104428) );
  NAND2_X1 U90793 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0 [1]), 
        .A2(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_7/S_0 [0]), .ZN(n82329)
         );
  OAI21_X1 U90794 ( .B1(n82314), .B2(n105022), .A(n82306), .ZN(n104429) );
  INV_X1 U90795 ( .A(n104429), .ZN(n104791) );
  NAND2_X1 U90796 ( .A1(n99635), .A2(n99636), .ZN(n104430) );
  INV_X1 U90797 ( .A(n104430), .ZN(n99567) );
  NOR3_X1 U90798 ( .A1(n82468), .A2(n57425), .A3(n105062), .ZN(n82475) );
  NOR4_X1 U90799 ( .A1(n82444), .A2(net82027), .A3(n62183), .A4(n62202), .ZN(
        n104431) );
  INV_X1 U90800 ( .A(n104431), .ZN(n82452) );
  NOR2_X1 U90801 ( .A1(n105545), .A2(n95109), .ZN(n95077) );
  NOR2_X1 U90802 ( .A1(n104432), .A2(n94931), .ZN(n81683) );
  INV_X1 U90803 ( .A(n81680), .ZN(n104432) );
  NOR3_X1 U90804 ( .A1(IR_in[31]), .A2(n82774), .A3(n81993), .ZN(n82005) );
  NOR4_X1 U90805 ( .A1(n104755), .A2(n104433), .A3(IR_in[1]), .A4(IR_in[0]), 
        .ZN(n81989) );
  INV_X1 U90806 ( .A(n82014), .ZN(n104433) );
  OAI21_X1 U90807 ( .B1(n105152), .B2(n104713), .A(net113081), .ZN(n82026) );
  NOR2_X1 U90808 ( .A1(n95651), .A2(n95623), .ZN(n104990) );
  NAND2_X1 U90809 ( .A1(n104450), .A2(n104434), .ZN(n82856) );
  NAND2_X1 U90810 ( .A1(n83114), .A2(n70652), .ZN(n104435) );
  INV_X1 U90811 ( .A(n104435), .ZN(n83295) );
  NAND2_X1 U90812 ( .A1(n100159), .A2(n100160), .ZN(n104436) );
  INV_X1 U90813 ( .A(n104436), .ZN(n99280) );
  AOI21_X1 U90814 ( .B1(n98973), .B2(n98971), .A(n106956), .ZN(n104455) );
  NOR2_X1 U90815 ( .A1(n97748), .A2(n97780), .ZN(n106125) );
  NAND2_X1 U90816 ( .A1(n99411), .A2(n99412), .ZN(n104437) );
  INV_X1 U90817 ( .A(n104437), .ZN(n99068) );
  NOR2_X1 U90818 ( .A1(n98366), .A2(n98367), .ZN(n104880) );
  NOR2_X1 U90819 ( .A1(n97449), .A2(n97487), .ZN(n104870) );
  NOR2_X1 U90820 ( .A1(n98232), .A2(n98090), .ZN(n106214) );
  XOR2_X1 U90821 ( .A(n82490), .B(n59478), .Z(n82241) );
  NOR2_X1 U90822 ( .A1(n98801), .A2(n95131), .ZN(n106340) );
  NOR2_X1 U90823 ( .A1(n96837), .A2(n96838), .ZN(n105392) );
  NOR2_X1 U90824 ( .A1(n96050), .A2(n96013), .ZN(n105446) );
  NOR2_X1 U90825 ( .A1(n95488), .A2(n95489), .ZN(n104978) );
  NOR2_X1 U90826 ( .A1(n97967), .A2(n98004), .ZN(n105284) );
  NOR2_X1 U90827 ( .A1(n97574), .A2(n97637), .ZN(n106141) );
  NOR2_X1 U90828 ( .A1(n97356), .A2(n97428), .ZN(n105351) );
  NOR2_X1 U90829 ( .A1(n96454), .A2(n96453), .ZN(n105415) );
  NOR2_X1 U90830 ( .A1(n96331), .A2(n96330), .ZN(n105423) );
  NOR2_X1 U90831 ( .A1(n96204), .A2(n96203), .ZN(n105431) );
  NOR2_X1 U90832 ( .A1(n96127), .A2(n106757), .ZN(n105438) );
  NOR2_X1 U90833 ( .A1(n104847), .A2(n96052), .ZN(n104889) );
  NOR2_X1 U90834 ( .A1(n95989), .A2(n95555), .ZN(n105452) );
  NOR2_X1 U90835 ( .A1(n95948), .A2(n95517), .ZN(n105456) );
  NOR2_X1 U90836 ( .A1(n95912), .A2(n104822), .ZN(n105465) );
  NOR2_X1 U90837 ( .A1(n95762), .A2(n95763), .ZN(n104957) );
  AOI21_X1 U90838 ( .B1(n95450), .B2(n94554), .A(n95726), .ZN(n104971) );
  NOR2_X1 U90839 ( .A1(n98005), .A2(n98060), .ZN(n105278) );
  NOR2_X1 U90840 ( .A1(n97840), .A2(n97931), .ZN(n105299) );
  NOR2_X1 U90841 ( .A1(n97710), .A2(n97816), .ZN(n105311) );
  NOR2_X1 U90842 ( .A1(n97612), .A2(n97673), .ZN(n105329) );
  NOR2_X1 U90843 ( .A1(n97031), .A2(n96969), .ZN(n105372) );
  NOR2_X1 U90844 ( .A1(n96933), .A2(n96995), .ZN(n104850) );
  NOR2_X1 U90845 ( .A1(n96801), .A2(n96910), .ZN(n105384) );
  NOR2_X1 U90846 ( .A1(n96416), .A2(n96486), .ZN(n105989) );
  AOI21_X1 U90847 ( .B1(n96010), .B2(n94771), .A(n96417), .ZN(n105927) );
  NOR2_X1 U90848 ( .A1(n96293), .A2(n96354), .ZN(n105979) );
  NOR2_X1 U90849 ( .A1(n96166), .A2(n96231), .ZN(n105996) );
  NOR2_X1 U90850 ( .A1(n95725), .A2(n95799), .ZN(n104935) );
  NOR2_X1 U90851 ( .A1(n95448), .A2(n95516), .ZN(n105974) );
  NOR2_X1 U90852 ( .A1(n95169), .A2(n106748), .ZN(n105535) );
  NOR2_X1 U90853 ( .A1(n94661), .A2(n94553), .ZN(n105605) );
  NOR4_X1 U90854 ( .A1(n105150), .A2(IR_in[4]), .A3(n82000), .A4(n82636), .ZN(
        n81981) );
  NOR2_X1 U90855 ( .A1(n81916), .A2(n86222), .ZN(n81881) );
  XOR2_X1 U90856 ( .A(n81808), .B(n99031), .Z(n81807) );
  AOI22_X1 U90857 ( .A1(n79776), .A2(\DLX_Datapath/ArithLogUnit/A_log [24]), 
        .B1(n104438), .B2(\DLX_Datapath/ArithLogUnit/B_log [24]), .ZN(n79775)
         );
  INV_X1 U90858 ( .A(n79778), .ZN(n104438) );
  NOR2_X1 U90859 ( .A1(n104439), .A2(n82274), .ZN(n105069) );
  INV_X1 U90860 ( .A(n82283), .ZN(n104439) );
  NAND2_X1 U90861 ( .A1(n81255), .A2(n104475), .ZN(n104490) );
  NAND2_X1 U90862 ( .A1(n107106), .A2(n59454), .ZN(n105042) );
  AOI22_X1 U90863 ( .A1(n99664), .A2(n99661), .B1(n107482), .B2(n99628), .ZN(
        n99582) );
  OAI21_X1 U90864 ( .B1(n62662), .B2(n107104), .A(n62661), .ZN(n100250) );
  NAND3_X2 U90865 ( .A1(n84067), .A2(n106280), .A3(n84086), .ZN(n84078) );
  NOR3_X1 U90866 ( .A1(n62190), .A2(n105057), .A3(n106697), .ZN(n104440) );
  INV_X1 U90867 ( .A(n104440), .ZN(n84062) );
  AOI21_X1 U90868 ( .B1(n104441), .B2(\DLX_Datapath/CWP_IDEX[2] ), .A(n111028), 
        .ZN(n107108) );
  XOR2_X1 U90869 ( .A(n105054), .B(n100394), .Z(n90135) );
  NOR2_X1 U90870 ( .A1(n104442), .A2(n104443), .ZN(n100204) );
  XOR2_X1 U90871 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [8]), .B(
        \DLX_Datapath/ArithLogUnit/B_mul [7]), .Z(n104472) );
  NAND2_X1 U90872 ( .A1(\DLX_Datapath/ArithLogUnit/A_add [4]), .A2(
        \DLX_Datapath/ArithLogUnit/B_add [4]), .ZN(n104444) );
  INV_X1 U90873 ( .A(n104444), .ZN(n104370) );
  XOR2_X1 U90874 ( .A(n100035), .B(n100012), .Z(n100002) );
  NAND2_X1 U90875 ( .A1(n99502), .A2(n99503), .ZN(n104445) );
  INV_X1 U90876 ( .A(n104445), .ZN(n99473) );
  NOR4_X1 U90877 ( .A1(n104446), .A2(n106931), .A3(n100228), .A4(n100229), 
        .ZN(n100195) );
  NAND2_X1 U90878 ( .A1(n99351), .A2(n99352), .ZN(n104447) );
  INV_X1 U90879 ( .A(n104447), .ZN(n83106) );
  NAND2_X1 U90880 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [2]), 
        .A2(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [3]), .ZN(n82500)
         );
  NAND2_X1 U90881 ( .A1(n99829), .A2(n99830), .ZN(n104448) );
  INV_X1 U90882 ( .A(n104448), .ZN(n99786) );
  NAND2_X1 U90883 ( .A1(n104909), .A2(n94434), .ZN(n95074) );
  NOR2_X1 U90884 ( .A1(n104449), .A2(n82603), .ZN(n82537) );
  INV_X1 U90885 ( .A(n82611), .ZN(n104449) );
  OAI21_X1 U90886 ( .B1(n82200), .B2(n105019), .A(n82202), .ZN(n80128) );
  NOR2_X1 U90887 ( .A1(n97486), .A2(n97547), .ZN(n105340) );
  NOR2_X1 U90888 ( .A1(n95651), .A2(n95623), .ZN(n104991) );
  NAND2_X1 U90889 ( .A1(n104450), .A2(n111065), .ZN(n82857) );
  OAI21_X1 U90890 ( .B1(n82628), .B2(n82624), .A(n81991), .ZN(n104451) );
  INV_X1 U90891 ( .A(n104451), .ZN(n81985) );
  NAND2_X1 U90892 ( .A1(n83162), .A2(n73821), .ZN(n104452) );
  INV_X1 U90893 ( .A(n104452), .ZN(n83381) );
  NAND2_X1 U90894 ( .A1(n83114), .A2(n74065), .ZN(n104453) );
  INV_X1 U90895 ( .A(n104453), .ZN(n83266) );
  XOR2_X1 U90896 ( .A(n82475), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [1]), .Z(n106817) );
  XOR2_X1 U90897 ( .A(n99161), .B(n104483), .Z(n99735) );
  XOR2_X1 U90898 ( .A(n82465), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [1]), .Z(n106819) );
  NAND2_X1 U90899 ( .A1(n99540), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .ZN(n104454) );
  INV_X1 U90900 ( .A(n104454), .ZN(n100132) );
  AOI21_X1 U90901 ( .B1(n100295), .B2(n69339), .A(n104455), .ZN(n99003) );
  NOR2_X1 U90902 ( .A1(n96679), .A2(n96777), .ZN(n104873) );
  AOI21_X1 U90903 ( .B1(n82167), .B2(n57425), .A(n82164), .ZN(n82150) );
  NOR2_X1 U90904 ( .A1(n98366), .A2(n98471), .ZN(n104824) );
  NOR2_X1 U90905 ( .A1(n95948), .A2(n95517), .ZN(n105455) );
  OAI21_X1 U90906 ( .B1(n82766), .B2(n82629), .A(n80100), .ZN(n80069) );
  NOR2_X1 U90907 ( .A1(n98801), .A2(n95131), .ZN(n106339) );
  NOR2_X1 U90908 ( .A1(n98499), .A2(n98537), .ZN(n105256) );
  NOR2_X1 U90909 ( .A1(n98232), .A2(n98090), .ZN(n106215) );
  NOR2_X1 U90910 ( .A1(n97449), .A2(n104691), .ZN(n106064) );
  NOR2_X1 U90911 ( .A1(n96910), .A2(n96837), .ZN(n105379) );
  NOR2_X1 U90912 ( .A1(n95585), .A2(n95622), .ZN(n104973) );
  NOR2_X1 U90913 ( .A1(n98538), .A2(n98611), .ZN(n105248) );
  NOR2_X1 U90914 ( .A1(n98005), .A2(n98024), .ZN(n106090) );
  NOR2_X1 U90915 ( .A1(n97967), .A2(n98004), .ZN(n105285) );
  NOR2_X1 U90916 ( .A1(n97840), .A2(n97877), .ZN(n105303) );
  NOR2_X1 U90917 ( .A1(n97748), .A2(n97816), .ZN(n105309) );
  NOR2_X1 U90918 ( .A1(n97710), .A2(n97780), .ZN(n106126) );
  NOR2_X1 U90919 ( .A1(n97574), .A2(n97673), .ZN(n105332) );
  NOR2_X1 U90920 ( .A1(n97356), .A2(n97428), .ZN(n105350) );
  NOR2_X1 U90921 ( .A1(n97318), .A2(n97355), .ZN(n105361) );
  NOR2_X1 U90922 ( .A1(n96969), .A2(n96995), .ZN(n104866) );
  NOR2_X1 U90923 ( .A1(n96933), .A2(n96970), .ZN(n104860) );
  AOI21_X1 U90924 ( .B1(n96560), .B2(n94771), .A(n96932), .ZN(n106030) );
  NOR2_X1 U90925 ( .A1(n96801), .A2(n96874), .ZN(n105389) );
  NOR2_X1 U90926 ( .A1(n96741), .A2(n96717), .ZN(n106013) );
  NOR2_X1 U90927 ( .A1(n96527), .A2(n106757), .ZN(n105412) );
  NOR2_X1 U90928 ( .A1(n96454), .A2(n96486), .ZN(n105985) );
  NOR2_X1 U90929 ( .A1(n96416), .A2(n96453), .ZN(n104932) );
  NOR2_X1 U90930 ( .A1(n96331), .A2(n96354), .ZN(n105981) );
  NOR2_X1 U90931 ( .A1(n96293), .A2(n96330), .ZN(n104959) );
  AOI21_X1 U90932 ( .B1(n96010), .B2(n94554), .A(n96294), .ZN(n105933) );
  NOR2_X1 U90933 ( .A1(n96204), .A2(n96231), .ZN(n105999) );
  NOR2_X1 U90934 ( .A1(n96166), .A2(n96203), .ZN(n104974) );
  NOR2_X1 U90935 ( .A1(n96088), .A2(n96013), .ZN(n104768) );
  NOR2_X1 U90936 ( .A1(n95949), .A2(n95912), .ZN(n105459) );
  NOR2_X1 U90937 ( .A1(n95762), .A2(n95763), .ZN(n104956) );
  NOR2_X1 U90938 ( .A1(n95725), .A2(n95726), .ZN(n105482) );
  NOR2_X1 U90939 ( .A1(n95689), .A2(n95555), .ZN(n105487) );
  NOR2_X1 U90940 ( .A1(n95488), .A2(n95516), .ZN(n104931) );
  NOR2_X1 U90941 ( .A1(n95448), .A2(n95489), .ZN(n105498) );
  NOR2_X1 U90942 ( .A1(n95073), .A2(n105951), .ZN(n104953) );
  NOR2_X1 U90943 ( .A1(n95037), .A2(n106748), .ZN(n105556) );
  NOR2_X1 U90944 ( .A1(n94970), .A2(n105566), .ZN(n105560) );
  NOR2_X1 U90945 ( .A1(n94931), .A2(n105575), .ZN(n105568) );
  NOR2_X1 U90946 ( .A1(n94623), .A2(n94553), .ZN(n105612) );
  OAI21_X1 U90947 ( .B1(n82249), .B2(n82300), .A(n82271), .ZN(n82269) );
  NOR2_X1 U90948 ( .A1(n104805), .A2(n105151), .ZN(n105890) );
  XOR2_X1 U90949 ( .A(n99012), .B(n81816), .Z(n81815) );
  OAI21_X1 U90950 ( .B1(net113102), .B2(n57427), .A(n82214), .ZN(n82213) );
  AOI22_X1 U90951 ( .A1(n79741), .A2(\DLX_Datapath/ArithLogUnit/A_log [28]), 
        .B1(n104456), .B2(\DLX_Datapath/ArithLogUnit/B_log [28]), .ZN(n79740)
         );
  INV_X1 U90952 ( .A(n79743), .ZN(n104456) );
  NAND2_X1 U90953 ( .A1(n100496), .A2(n106958), .ZN(n104457) );
  INV_X1 U90954 ( .A(n104457), .ZN(\DLX_Datapath/RegisterFile/N46898 ) );
  OAI21_X1 U90955 ( .B1(n108852), .B2(n82024), .A(n82031), .ZN(n82028) );
  NAND2_X1 U90956 ( .A1(n99899), .A2(n99900), .ZN(n104458) );
  INV_X1 U90957 ( .A(n104458), .ZN(n99839) );
  XNOR2_X1 U90958 ( .A(n82686), .B(n82687), .ZN(n104848) );
  NOR3_X1 U90959 ( .A1(n107104), .A2(n64266), .A3(n104950), .ZN(n104459) );
  INV_X1 U90960 ( .A(n104459), .ZN(n104903) );
  NOR3_X1 U90961 ( .A1(n105057), .A2(n104582), .A3(n106697), .ZN(n104460) );
  INV_X1 U90962 ( .A(n104460), .ZN(n84066) );
  OAI21_X1 U90963 ( .B1(n99632), .B2(n99631), .A(n104461), .ZN(n104462) );
  INV_X1 U90964 ( .A(n99634), .ZN(n104461) );
  INV_X1 U90965 ( .A(n104462), .ZN(n99633) );
  OAI21_X1 U90966 ( .B1(n99814), .B2(n99813), .A(n104463), .ZN(n104464) );
  INV_X1 U90967 ( .A(n99816), .ZN(n104463) );
  INV_X1 U90968 ( .A(n104464), .ZN(n99815) );
  INV_X1 U90969 ( .A(n104465), .ZN(n104910) );
  NAND2_X1 U90970 ( .A1(n100396), .A2(n100397), .ZN(n104466) );
  INV_X1 U90971 ( .A(n104466), .ZN(n100391) );
  NOR4_X1 U90972 ( .A1(n81208), .A2(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] ), 
        .A3(n81238), .A4(n105058), .ZN(n85207) );
  NAND2_X1 U90973 ( .A1(\DLX_Datapath/ArithLogUnit/A_add [28]), .A2(
        \DLX_Datapath/ArithLogUnit/B_add [28]), .ZN(n104467) );
  INV_X1 U90974 ( .A(n104467), .ZN(n104369) );
  NAND2_X1 U90975 ( .A1(\DLX_Datapath/ArithLogUnit/A_add [24]), .A2(
        \DLX_Datapath/ArithLogUnit/B_add [24]), .ZN(n104468) );
  INV_X1 U90976 ( .A(n104468), .ZN(n104376) );
  NAND2_X1 U90977 ( .A1(\DLX_Datapath/ArithLogUnit/A_add [20]), .A2(
        \DLX_Datapath/ArithLogUnit/B_add [20]), .ZN(n104469) );
  INV_X1 U90978 ( .A(n104469), .ZN(n104375) );
  NAND2_X1 U90979 ( .A1(\DLX_Datapath/ArithLogUnit/A_add [16]), .A2(
        \DLX_Datapath/ArithLogUnit/B_add [16]), .ZN(n104470) );
  INV_X1 U90980 ( .A(n104470), .ZN(n104374) );
  NAND2_X1 U90981 ( .A1(\DLX_Datapath/ArithLogUnit/A_add [12]), .A2(
        \DLX_Datapath/ArithLogUnit/B_add [12]), .ZN(n104471) );
  INV_X1 U90982 ( .A(n104471), .ZN(n104373) );
  AOI22_X1 U90983 ( .A1(\DLX_Datapath/ArithLogUnit/B_mul [8]), .A2(n100086), 
        .B1(n104472), .B2(\DLX_Datapath/ArithLogUnit/B_mul [9]), .ZN(n100062)
         );
  NAND2_X1 U90984 ( .A1(\DLX_Datapath/ArithLogUnit/A_add [8]), .A2(
        \DLX_Datapath/ArithLogUnit/B_add [8]), .ZN(n104473) );
  INV_X1 U90985 ( .A(n104473), .ZN(n104372) );
  NOR2_X1 U90986 ( .A1(net2465244), .A2(net2465245), .ZN(n105032) );
  XOR2_X1 U90987 ( .A(n100004), .B(n99981), .Z(n99971) );
  NOR4_X1 U90988 ( .A1(n104474), .A2(n100273), .A3(n100274), .A4(n100275), 
        .ZN(n100199) );
  INV_X1 U90989 ( .A(n100268), .ZN(n104474) );
  OR2_X1 U90990 ( .A1(n95412), .A2(n104815), .ZN(n104878) );
  NAND2_X1 U90991 ( .A1(IR_in[7]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [3]), .ZN(n104475) );
  INV_X1 U90992 ( .A(n104475), .ZN(n104740) );
  XOR2_X1 U90993 ( .A(n104757), .B(\add_0_root_r2411/carry[7] ), .Z(n90136) );
  AOI21_X1 U90994 ( .B1(n105040), .B2(n105043), .A(n82200), .ZN(n104913) );
  OAI21_X1 U90995 ( .B1(n106936), .B2(n106845), .A(n82280), .ZN(n100318) );
  OAI21_X1 U90996 ( .B1(n99651), .B2(n99650), .A(n104476), .ZN(n104477) );
  INV_X1 U90997 ( .A(n99649), .ZN(n104476) );
  INV_X1 U90998 ( .A(n104477), .ZN(n99609) );
  XOR2_X1 U90999 ( .A(n100090), .B(n100078), .Z(n100067) );
  NOR3_X1 U91000 ( .A1(n109310), .A2(\DLX_Datapath/ArithLogUnit/B_mul [4]), 
        .A3(\DLX_Datapath/ArithLogUnit/B_mul [3]), .ZN(n99625) );
  NAND2_X1 U91001 ( .A1(n99421), .A2(n99422), .ZN(n104478) );
  INV_X1 U91002 ( .A(n104478), .ZN(n99392) );
  NOR3_X1 U91003 ( .A1(n83103), .A2(n83094), .A3(n83096), .ZN(n83097) );
  NOR3_X1 U91004 ( .A1(n106753), .A2(n94851), .A3(n94852), .ZN(n94732) );
  NOR2_X1 U91005 ( .A1(n105152), .A2(n104713), .ZN(n105889) );
  AOI22_X1 U91006 ( .A1(n82220), .A2(n57427), .B1(n104802), .B2(n104887), .ZN(
        n82219) );
  NOR2_X1 U91007 ( .A1(n95585), .A2(n95651), .ZN(n105965) );
  OAI21_X1 U91008 ( .B1(n104479), .B2(n82624), .A(n82645), .ZN(n111121) );
  INV_X1 U91009 ( .A(n80042), .ZN(n104479) );
  OAI21_X1 U91010 ( .B1(n105204), .B2(n106328), .A(n86230), .ZN(n81879) );
  NAND2_X1 U91011 ( .A1(n82852), .A2(DataIn_b[7]), .ZN(n104480) );
  INV_X1 U91012 ( .A(n104480), .ZN(n82821) );
  NOR3_X1 U91013 ( .A1(n111141), .A2(n80067), .A3(n80064), .ZN(n80086) );
  NAND2_X1 U91014 ( .A1(n83162), .A2(n74385), .ZN(n104481) );
  INV_X1 U91015 ( .A(n104481), .ZN(n83352) );
  NAND2_X1 U91016 ( .A1(n83114), .A2(n70363), .ZN(n104482) );
  INV_X1 U91017 ( .A(n104482), .ZN(n83113) );
  XOR2_X1 U91018 ( .A(n99101), .B(n99100), .Z(n99493) );
  NAND2_X1 U91019 ( .A1(n104794), .A2(n82311), .ZN(n104891) );
  NAND2_X1 U91020 ( .A1(n99736), .A2(n99737), .ZN(n104483) );
  INV_X1 U91021 ( .A(n104483), .ZN(n99158) );
  XOR2_X1 U91022 ( .A(n99181), .B(n99180), .Z(n99827) );
  NAND2_X1 U91023 ( .A1(n99428), .A2(
        \DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .ZN(n104484) );
  INV_X1 U91024 ( .A(n104484), .ZN(n100029) );
  XOR2_X1 U91025 ( .A(n99218), .B(n99217), .Z(n99995) );
  XOR2_X1 U91026 ( .A(n105063), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_3/S_0 [3]), .Z(n106820) );
  NOR2_X1 U91027 ( .A1(n97318), .A2(n97392), .ZN(n104864) );
  NOR2_X1 U91028 ( .A1(n98499), .A2(n98611), .ZN(n104826) );
  NOR2_X1 U91029 ( .A1(n98406), .A2(n98471), .ZN(n105260) );
  AOI21_X1 U91030 ( .B1(n96560), .B2(n94398), .A(n96680), .ZN(n106022) );
  NAND2_X1 U91031 ( .A1(n105129), .A2(n94331), .ZN(n106006) );
  NOR2_X1 U91032 ( .A1(n96050), .A2(n96013), .ZN(n105445) );
  NOR2_X1 U91033 ( .A1(n98801), .A2(n95131), .ZN(n106338) );
  NOR2_X1 U91034 ( .A1(n98538), .A2(n98537), .ZN(n104886) );
  NOR2_X1 U91035 ( .A1(n98366), .A2(n98367), .ZN(n104879) );
  NOR2_X1 U91036 ( .A1(n98232), .A2(n98090), .ZN(n106213) );
  NOR2_X1 U91037 ( .A1(n98089), .A2(n94999), .ZN(n106226) );
  NOR2_X1 U91038 ( .A1(n97967), .A2(n98024), .ZN(n106088) );
  NOR2_X1 U91039 ( .A1(n98004), .A2(n98005), .ZN(n105288) );
  NOR2_X1 U91040 ( .A1(n97840), .A2(n97895), .ZN(n106119) );
  NOR2_X1 U91041 ( .A1(n97877), .A2(n97878), .ZN(n105305) );
  NOR2_X1 U91042 ( .A1(n97747), .A2(n97748), .ZN(n105317) );
  NOR2_X1 U91043 ( .A1(n97710), .A2(n97711), .ZN(n105322) );
  NOR2_X1 U91044 ( .A1(n97574), .A2(n97637), .ZN(n106140) );
  NOR2_X1 U91045 ( .A1(n97611), .A2(n97612), .ZN(n105337) );
  NOR2_X1 U91046 ( .A1(n97449), .A2(n104695), .ZN(n104853) );
  NOR2_X1 U91047 ( .A1(n97486), .A2(n97487), .ZN(n105347) );
  NOR2_X1 U91048 ( .A1(n97356), .A2(n97355), .ZN(n105363) );
  NOR2_X1 U91049 ( .A1(n96969), .A2(n96970), .ZN(n105377) );
  NOR2_X1 U91050 ( .A1(n96933), .A2(n104697), .ZN(n104875) );
  NOR2_X1 U91051 ( .A1(n96910), .A2(n96837), .ZN(n105381) );
  NOR2_X1 U91052 ( .A1(n96801), .A2(n96838), .ZN(n105395) );
  NOR2_X1 U91053 ( .A1(n96717), .A2(n96777), .ZN(n105399) );
  NOR2_X1 U91054 ( .A1(n96679), .A2(n96741), .ZN(n104855) );
  NOR2_X1 U91055 ( .A1(n96454), .A2(n96453), .ZN(n105416) );
  NOR2_X1 U91056 ( .A1(n96416), .A2(n96417), .ZN(n105923) );
  NOR2_X1 U91057 ( .A1(n96331), .A2(n96330), .ZN(n105424) );
  NOR2_X1 U91058 ( .A1(n96293), .A2(n96294), .ZN(n105930) );
  NOR2_X1 U91059 ( .A1(n96204), .A2(n96203), .ZN(n105432) );
  NOR2_X1 U91060 ( .A1(n96166), .A2(n96167), .ZN(n105435) );
  NOR2_X1 U91061 ( .A1(n96127), .A2(n106757), .ZN(n105440) );
  NOR2_X1 U91062 ( .A1(n104847), .A2(n96052), .ZN(n104888) );
  NOR2_X1 U91063 ( .A1(n95989), .A2(n95555), .ZN(n105453) );
  NOR2_X1 U91064 ( .A1(n95948), .A2(n95517), .ZN(n105457) );
  NOR2_X1 U91065 ( .A1(n95912), .A2(n104822), .ZN(n105466) );
  NOR2_X1 U91066 ( .A1(n95799), .A2(n95763), .ZN(n105478) );
  NOR2_X1 U91067 ( .A1(n95725), .A2(n95762), .ZN(n104947) );
  AOI21_X1 U91068 ( .B1(n95450), .B2(n94554), .A(n95726), .ZN(n104969) );
  AOI21_X1 U91069 ( .B1(n95687), .B2(n105602), .A(n104703), .ZN(n104938) );
  NOR2_X1 U91070 ( .A1(n95623), .A2(n95622), .ZN(n105490) );
  NOR2_X1 U91071 ( .A1(n95488), .A2(n95489), .ZN(n104977) );
  NOR2_X1 U91072 ( .A1(n95448), .A2(n95449), .ZN(n104926) );
  NOR2_X1 U91073 ( .A1(n95109), .A2(n105951), .ZN(n105947) );
  NOR2_X1 U91074 ( .A1(n95073), .A2(n105545), .ZN(n105542) );
  NOR2_X1 U91075 ( .A1(n95037), .A2(n106748), .ZN(n105557) );
  NOR2_X1 U91076 ( .A1(n94931), .A2(n105566), .ZN(n105563) );
  AOI21_X1 U91077 ( .B1(n94932), .B2(n94258), .A(n105575), .ZN(n105572) );
  NOR2_X1 U91078 ( .A1(n94623), .A2(n94553), .ZN(n105614) );
  NAND2_X1 U91079 ( .A1(n82015), .A2(IR_in[4]), .ZN(n104485) );
  INV_X1 U91080 ( .A(n104485), .ZN(n82012) );
  NOR3_X1 U91081 ( .A1(n57430), .A2(n82490), .A3(n105068), .ZN(n104915) );
  XOR2_X1 U91082 ( .A(n105033), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [3]), .Z(n106818) );
  AOI22_X1 U91083 ( .A1(n81805), .A2(\DLX_Datapath/MUX_HDU_ALUInA [4]), .B1(
        n100153), .B2(n81804), .ZN(n104486) );
  INV_X1 U91084 ( .A(n104486), .ZN(\DLX_Datapath/ArithLogUnit/N117 ) );
  OAI21_X1 U91085 ( .B1(net113081), .B2(n104494), .A(n82107), .ZN(n82106) );
  AOI22_X1 U91086 ( .A1(n79875), .A2(\DLX_Datapath/ArithLogUnit/A_log [12]), 
        .B1(n104487), .B2(\DLX_Datapath/ArithLogUnit/B_log [12]), .ZN(n79874)
         );
  INV_X1 U91087 ( .A(n79877), .ZN(n104487) );
  OAI21_X1 U91088 ( .B1(n80100), .B2(n105151), .A(n81878), .ZN(n104488) );
  INV_X1 U91089 ( .A(n104488), .ZN(n81877) );
  OAI21_X1 U91090 ( .B1(n107418), .B2(n82024), .A(n82025), .ZN(n82017) );
  NAND2_X1 U91091 ( .A1(n69765), .A2(n106958), .ZN(n104489) );
  INV_X1 U91092 ( .A(n104489), .ZN(\DLX_Datapath/RegisterFile/N46899 ) );
  CLKBUF_X1 U91093 ( .A(n81478), .Z(n104766) );
  CLKBUF_X1 U91094 ( .A(n81478), .Z(n104765) );
  CLKBUF_X1 U91095 ( .A(n104735), .Z(n104737) );
  CLKBUF_X1 U91096 ( .A(n104735), .Z(n104736) );
  CLKBUF_X1 U91097 ( .A(n95840), .Z(n104818) );
  CLKBUF_X1 U91098 ( .A(n95840), .Z(n104817) );
  CLKBUF_X1 U91099 ( .A(n80001), .Z(net73629) );
  OR2_X1 U91100 ( .A1(n104490), .A2(n104739), .ZN(n104747) );
  INV_X1 U91101 ( .A(n82682), .ZN(n104900) );
  INV_X1 U91102 ( .A(net112469), .ZN(n104754) );
  INV_X1 U91103 ( .A(n82389), .ZN(n104796) );
  INV_X1 U91104 ( .A(n82388), .ZN(n104795) );
  INV_X1 U91105 ( .A(n82707), .ZN(n106807) );
  INV_X1 U91106 ( .A(n82286), .ZN(n104761) );
  INV_X1 U91107 ( .A(n82420), .ZN(net68723) );
  INV_X1 U91108 ( .A(n81255), .ZN(net68722) );
  INV_X1 U91109 ( .A(n104811), .ZN(n104728) );
  INV_X1 U91110 ( .A(n86230), .ZN(n111026) );
  CLKBUF_X1 U91111 ( .A(n82248), .Z(n105153) );
  INV_X1 U91112 ( .A(n82268), .ZN(n105027) );
  NAND2_X1 U91113 ( .A1(\DLX_Datapath/RegisterFile/N9337 ), .A2(n98940), .ZN(
        n104491) );
  CLKBUF_X3 U91114 ( .A(n96133), .Z(n104989) );
  CLKBUF_X1 U91115 ( .A(n82292), .Z(n105065) );
  CLKBUF_X1 U91116 ( .A(n98802), .Z(n104492) );
  CLKBUF_X1 U91117 ( .A(n94081), .Z(n104493) );
  CLKBUF_X1 U91118 ( .A(n94509), .Z(n104714) );
  INV_X1 U91119 ( .A(n59516), .ZN(n107096) );
  CLKBUF_X1 U91120 ( .A(n94509), .Z(n104715) );
  CLKBUF_X1 U91121 ( .A(n94509), .Z(n104716) );
  CLKBUF_X1 U91122 ( .A(n95520), .Z(n104845) );
  CLKBUF_X1 U91123 ( .A(n95520), .Z(n104846) );
  CLKBUF_X1 U91124 ( .A(n96357), .Z(n104837) );
  CLKBUF_X1 U91125 ( .A(n96357), .Z(n104838) );
  INV_X1 U91126 ( .A(n95074), .ZN(n105545) );
  INV_X1 U91127 ( .A(n94896), .ZN(n105575) );
  INV_X1 U91128 ( .A(n81688), .ZN(n105951) );
  CLKBUF_X1 U91129 ( .A(n95802), .Z(n104841) );
  CLKBUF_X1 U91130 ( .A(n95802), .Z(n104842) );
  NOR2_X1 U91131 ( .A1(\DLX_Datapath/CWP_IDEX[2] ), .A2(n104495), .ZN(n104500)
         );
  NAND2_X1 U91132 ( .A1(n94892), .A2(n105132), .ZN(n104503) );
  NAND2_X1 U91133 ( .A1(n94934), .A2(n105124), .ZN(n104504) );
  OR2_X1 U91134 ( .A1(n82317), .A2(n82315), .ZN(n104505) );
  XOR2_X1 U91135 ( .A(n82450), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [2]), .Z(n104507) );
  OR2_X1 U91136 ( .A1(n107126), .A2(n94895), .ZN(n104508) );
  XNOR2_X1 U91137 ( .A(n57429), .B(n105153), .ZN(n104509) );
  OR2_X1 U91138 ( .A1(IR_in[12]), .A2(n82318), .ZN(n104510) );
  OR2_X1 U91139 ( .A1(n100356), .A2(n100357), .ZN(n104511) );
  OR2_X1 U91140 ( .A1(n100365), .A2(n100366), .ZN(n104524) );
  INV_X1 U91141 ( .A(n94773), .ZN(n105591) );
  INV_X1 U91142 ( .A(n81967), .ZN(net112601) );
  NOR2_X1 U91158 ( .A1(n81336), .A2(n105092), .ZN(n104687) );
  CLKBUF_X2 U91159 ( .A(n81339), .Z(n106176) );
  CLKBUF_X3 U91160 ( .A(n94472), .Z(n104986) );
  CLKBUF_X3 U91161 ( .A(n94333), .Z(n104984) );
  NOR2_X1 U91162 ( .A1(n94970), .A2(n105954), .ZN(n104688) );
  NOR2_X1 U91163 ( .A1(n94970), .A2(n105954), .ZN(n104689) );
  CLKBUF_X3 U91164 ( .A(n81326), .Z(n104882) );
  CLKBUF_X3 U91165 ( .A(n96684), .Z(n105404) );
  NOR2_X1 U91166 ( .A1(n81564), .A2(n105090), .ZN(n104690) );
  CLKBUF_X1 U91167 ( .A(n81658), .Z(n105966) );
  NOR2_X1 U91168 ( .A1(n81459), .A2(n105092), .ZN(n104691) );
  CLKBUF_X1 U91169 ( .A(n81774), .Z(n105917) );
  NOR2_X1 U91170 ( .A1(n81443), .A2(n105092), .ZN(n104692) );
  CLKBUF_X2 U91171 ( .A(n81446), .Z(n106075) );
  OR2_X1 U91172 ( .A1(n107400), .A2(n105630), .ZN(n104693) );
  NAND2_X1 U91173 ( .A1(n104693), .A2(n94529), .ZN(
        \DLX_Datapath/RegisterFile/N26619 ) );
  NAND2_X1 U91174 ( .A1(n69346), .A2(\DLX_Datapath/IR_EXMEM[20] ), .ZN(n104995) );
  NOR2_X1 U91175 ( .A1(n81273), .A2(n105095), .ZN(n104694) );
  CLKBUF_X2 U91176 ( .A(n81276), .Z(n106249) );
  CLKBUF_X3 U91177 ( .A(n95415), .Z(n104982) );
  CLKBUF_X1 U91178 ( .A(n96839), .Z(n105390) );
  NOR2_X1 U91179 ( .A1(n81513), .A2(n105092), .ZN(n104695) );
  CLKBUF_X3 U91180 ( .A(n104503), .Z(n105413) );
  CLKBUF_X3 U91181 ( .A(n81690), .Z(n105946) );
  NAND2_X1 U91182 ( .A1(n100463), .A2(net113153), .ZN(n104696) );
  INV_X1 U91183 ( .A(n104696), .ZN(n80153) );
  CLKBUF_X3 U91184 ( .A(n80153), .Z(n106342) );
  INV_X1 U91185 ( .A(net113153), .ZN(net113157) );
  CLKBUF_X3 U91186 ( .A(n95041), .Z(n105548) );
  NOR2_X1 U91187 ( .A1(n81540), .A2(n105091), .ZN(n104697) );
  OR2_X1 U91188 ( .A1(n104811), .A2(n82280), .ZN(n104698) );
  NOR2_X1 U91189 ( .A1(n104810), .A2(n104698), .ZN(n104699) );
  INV_X1 U91190 ( .A(n104699), .ZN(n82024) );
  CLKBUF_X1 U91191 ( .A(n82688), .Z(n104700) );
  NOR2_X1 U91192 ( .A1(n95838), .A2(n105089), .ZN(n104701) );
  CLKBUF_X3 U91193 ( .A(n94899), .Z(n105569) );
  OR2_X1 U91194 ( .A1(n81281), .A2(n105470), .ZN(n104702) );
  NAND2_X1 U91195 ( .A1(n104702), .A2(n95859), .ZN(
        \DLX_Datapath/RegisterFile/N25464 ) );
  CLKBUF_X1 U91196 ( .A(n98166), .Z(n105273) );
  CLKBUF_X2 U91197 ( .A(n95133), .Z(n105536) );
  CLKBUF_X1 U91198 ( .A(n96802), .Z(n105396) );
  CLKBUF_X3 U91199 ( .A(n95077), .Z(n105539) );
  NOR2_X1 U91200 ( .A1(n95652), .A2(n105089), .ZN(n104703) );
  OR2_X1 U91201 ( .A1(n81629), .A2(n105269), .ZN(n104704) );
  NAND2_X1 U91202 ( .A1(n104704), .A2(n98311), .ZN(
        \DLX_Datapath/RegisterFile/N23075 ) );
  CLKBUF_X1 U91203 ( .A(n97512), .Z(n105344) );
  CLKBUF_X2 U91204 ( .A(n81476), .Z(n106059) );
  CLKBUF_X1 U91205 ( .A(n81493), .Z(n106058) );
  INV_X1 U91206 ( .A(n104751), .ZN(n104752) );
  CLKBUF_X1 U91207 ( .A(n107147), .Z(n104705) );
  NOR2_X1 U91208 ( .A1(n82330), .A2(n105151), .ZN(n104706) );
  AND2_X2 U91209 ( .A1(n104811), .A2(n104785), .ZN(n104708) );
  CLKBUF_X3 U91210 ( .A(n80041), .Z(n105152) );
  CLKBUF_X2 U91211 ( .A(n105030), .Z(n105045) );
  INV_X1 U91212 ( .A(net113152), .ZN(net113155) );
  INV_X1 U91213 ( .A(net113153), .ZN(net113159) );
  OR2_X1 U91214 ( .A1(n81383), .A2(n105421), .ZN(n104709) );
  NAND2_X1 U91215 ( .A1(n104709), .A2(n96368), .ZN(
        \DLX_Datapath/RegisterFile/N24992 ) );
  INV_X1 U91216 ( .A(n98940), .ZN(n104778) );
  CLKBUF_X3 U91217 ( .A(n94508), .Z(n105627) );
  OR2_X1 U91218 ( .A1(n82278), .A2(net73629), .ZN(n82608) );
  OR2_X1 U91219 ( .A1(n62247), .A2(net113091), .ZN(n104710) );
  NAND2_X1 U91220 ( .A1(n81877), .A2(n104710), .ZN(n62245) );
  OR2_X1 U91221 ( .A1(n81383), .A2(n106006), .ZN(n104711) );
  NAND2_X1 U91222 ( .A1(n104711), .A2(n96609), .ZN(
        \DLX_Datapath/RegisterFile/N24768 ) );
  CLKBUF_X3 U91223 ( .A(n105017), .Z(n105161) );
  CLKBUF_X3 U91224 ( .A(n105017), .Z(n105160) );
  OR2_X1 U91225 ( .A1(n81629), .A2(n105273), .ZN(n104712) );
  NAND2_X1 U91226 ( .A1(n98176), .A2(n104712), .ZN(
        \DLX_Datapath/RegisterFile/N23203 ) );
  NAND2_X1 U91227 ( .A1(n82280), .A2(n104761), .ZN(n104713) );
  INV_X1 U91228 ( .A(n82280), .ZN(n105014) );
  NOR2_X1 U91229 ( .A1(n104508), .A2(n94894), .ZN(n94893) );
  XNOR2_X1 U91230 ( .A(
        \add_0_root_sub_0_root_DLX_Datapath/RegisterFile/add_172/carry[6] ), 
        .B(\DLX_Datapath/RegisterFile/old_CWP2[2] ), .ZN(n104717) );
  CLKBUF_X1 U91231 ( .A(n81526), .Z(n106037) );
  CLKBUF_X3 U91232 ( .A(n98304), .Z(n105268) );
  NOR2_X1 U91233 ( .A1(n96012), .A2(n96013), .ZN(n104718) );
  NOR2_X1 U91234 ( .A1(n96012), .A2(n96013), .ZN(n104719) );
  CLKBUF_X3 U91235 ( .A(n81293), .Z(n106223) );
  CLKBUF_X2 U91236 ( .A(n97200), .Z(n105367) );
  OR2_X1 U91237 ( .A1(n107147), .A2(n104500), .ZN(n104721) );
  INV_X1 U91238 ( .A(n104787), .ZN(n104720) );
  OR2_X1 U91239 ( .A1(n104720), .A2(n104500), .ZN(n104994) );
  CLKBUF_X1 U91240 ( .A(n99340), .Z(n104722) );
  CLKBUF_X1 U91241 ( .A(n86284), .Z(n104723) );
  NOR2_X1 U91242 ( .A1(n81439), .A2(n105091), .ZN(n104724) );
  CLKBUF_X2 U91243 ( .A(n97137), .Z(n105368) );
  NOR2_X1 U91244 ( .A1(n81476), .A2(n105090), .ZN(n104725) );
  OR2_X1 U91245 ( .A1(n81378), .A2(n106059), .ZN(n104726) );
  NAND2_X1 U91246 ( .A1(n97174), .A2(n104726), .ZN(
        \DLX_Datapath/RegisterFile/N24200 ) );
  CLKBUF_X3 U91247 ( .A(n81264), .Z(n106265) );
  CLKBUF_X3 U91248 ( .A(n97395), .Z(n105353) );
  CLKBUF_X3 U91249 ( .A(n104504), .Z(n106229) );
  AND2_X2 U91250 ( .A1(n104727), .A2(n100377), .ZN(n82694) );
  NOR2_X1 U91251 ( .A1(n104500), .A2(n107147), .ZN(n104727) );
  NOR2_X1 U91252 ( .A1(n104728), .A2(n82280), .ZN(n104729) );
  AND2_X2 U91253 ( .A1(n105059), .A2(n105060), .ZN(n104730) );
  AND2_X2 U91254 ( .A1(n97235), .A2(n97296), .ZN(n104731) );
  CLKBUF_X3 U91255 ( .A(n96683), .Z(n105406) );
  CLKBUF_X1 U91256 ( .A(n80041), .Z(n105150) );
  CLKBUF_X3 U91257 ( .A(n97360), .Z(n105357) );
  CLKBUF_X1 U91258 ( .A(n104815), .Z(n104732) );
  AND2_X2 U91259 ( .A1(n96597), .A2(n96598), .ZN(n104733) );
  OR2_X1 U91260 ( .A1(n106345), .A2(n104920), .ZN(n104734) );
  OR2_X1 U91261 ( .A1(n106345), .A2(n104920), .ZN(n104735) );
  OR2_X1 U91262 ( .A1(n82277), .A2(net73629), .ZN(n82609) );
  CLKBUF_X3 U91263 ( .A(n81937), .Z(n105154) );
  NOR2_X1 U91264 ( .A1(n104739), .A2(n104740), .ZN(n104738) );
  INV_X1 U91265 ( .A(n104738), .ZN(n82091) );
  AND2_X2 U91266 ( .A1(n82422), .A2(n104756), .ZN(n104739) );
  INV_X1 U91267 ( .A(n104743), .ZN(net71745) );
  XNOR2_X1 U91268 ( .A(n104741), .B(n100252), .ZN(n100251) );
  CLKBUF_X2 U91269 ( .A(n106345), .Z(n106346) );
  INV_X1 U91270 ( .A(net113152), .ZN(net113154) );
  XOR2_X1 U91271 ( .A(n59454), .B(n59516), .Z(n94253) );
  CLKBUF_X1 U91272 ( .A(net2465244), .Z(n104912) );
  OAI21_X1 U91273 ( .B1(net113091), .B2(n104581), .A(n82095), .ZN(n82094) );
  NAND2_X1 U91274 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [1]), 
        .A2(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [2]), .ZN(net82027)
         );
  NOR2_X1 U91275 ( .A1(IR_in[9]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [1]), .ZN(n104744) );
  AOI21_X1 U91276 ( .B1(n104746), .B2(n104747), .A(n104748), .ZN(n104745) );
  NOR2_X1 U91277 ( .A1(IR_in[10]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [2]), .ZN(n104749) );
  NOR2_X1 U91278 ( .A1(n104745), .A2(n104749), .ZN(n104750) );
  NOR2_X1 U91279 ( .A1(n104744), .A2(n82420), .ZN(n104746) );
  NAND2_X1 U91280 ( .A1(IR_in[11]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_2/S_0 [3]), .ZN(n104751) );
  CLKBUF_X1 U91281 ( .A(net113102), .Z(n104753) );
  OR2_X1 U91282 ( .A1(IR_in[7]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [3]), .ZN(n104756) );
  INV_X1 U91283 ( .A(IR_in[6]), .ZN(n104755) );
  NAND2_X1 U91284 ( .A1(net113538), .A2(net112383), .ZN(n82424) );
  NAND2_X1 U91285 ( .A1(net113538), .A2(n104754), .ZN(n82423) );
  CLKBUF_X3 U91286 ( .A(n104922), .Z(n104757) );
  OR2_X1 U91287 ( .A1(n104913), .A2(n104783), .ZN(n104758) );
  XNOR2_X1 U91288 ( .A(n105081), .B(n57426), .ZN(n104759) );
  NAND2_X1 U91289 ( .A1(n105085), .A2(n82306), .ZN(n104760) );
  INV_X1 U91290 ( .A(n107128), .ZN(n104762) );
  INV_X1 U91291 ( .A(n104814), .ZN(n90137) );
  NOR2_X1 U91292 ( .A1(n105083), .A2(n104914), .ZN(n104763) );
  NOR2_X1 U91293 ( .A1(n97199), .A2(n97061), .ZN(n104764) );
  CLKBUF_X3 U91294 ( .A(n96056), .Z(n104769) );
  CLKBUF_X3 U91295 ( .A(n96056), .Z(n104770) );
  CLKBUF_X1 U91296 ( .A(net71745), .Z(net112358) );
  CLKBUF_X2 U91297 ( .A(n96623), .Z(n105408) );
  OR2_X1 U91298 ( .A1(n107406), .A2(n105629), .ZN(n104771) );
  NAND2_X1 U91299 ( .A1(n94533), .A2(n104771), .ZN(
        \DLX_Datapath/RegisterFile/N26616 ) );
  OR2_X1 U91300 ( .A1(n107412), .A2(n105629), .ZN(n104772) );
  NAND2_X1 U91301 ( .A1(n94537), .A2(n104772), .ZN(
        \DLX_Datapath/RegisterFile/N26613 ) );
  AND2_X2 U91302 ( .A1(n107129), .A2(n98944), .ZN(n104774) );
  OR2_X1 U91303 ( .A1(n111058), .A2(n105630), .ZN(n104775) );
  NAND2_X1 U91304 ( .A1(n94550), .A2(n104775), .ZN(
        \DLX_Datapath/RegisterFile/N26604 ) );
  OR2_X1 U91305 ( .A1(n107392), .A2(n105629), .ZN(n104776) );
  NAND2_X1 U91306 ( .A1(n104776), .A2(n94524), .ZN(
        \DLX_Datapath/RegisterFile/N26623 ) );
  AND2_X2 U91307 ( .A1(n97237), .A2(n97260), .ZN(n104777) );
  CLKBUF_X3 U91308 ( .A(n81554), .Z(n106028) );
  XNOR2_X1 U91309 ( .A(\DLX_Datapath/RegisterFile/N9337 ), .B(n104778), .ZN(
        n94895) );
  NOR2_X1 U91310 ( .A1(n81293), .A2(n105094), .ZN(n104779) );
  OR2_X1 U91311 ( .A1(n106223), .A2(n81394), .ZN(n104780) );
  NAND2_X1 U91312 ( .A1(n104780), .A2(n98223), .ZN(
        \DLX_Datapath/RegisterFile/N23155 ) );
  OAI21_X1 U91313 ( .B1(n80056), .B2(n111118), .A(n105165), .ZN(n104781) );
  INV_X1 U91314 ( .A(n104920), .ZN(n104788) );
  XNOR2_X1 U91315 ( .A(n104782), .B(n82380), .ZN(n82180) );
  XNOR2_X1 U91316 ( .A(n82381), .B(n62204), .ZN(n104782) );
  NOR2_X1 U91317 ( .A1(n104760), .A2(n104914), .ZN(n104783) );
  CLKBUF_X3 U91318 ( .A(n97062), .Z(n105128) );
  XNOR2_X1 U91319 ( .A(n105081), .B(n57426), .ZN(n104784) );
  AOI21_X1 U91320 ( .B1(n81921), .B2(n82280), .A(net113154), .ZN(n104785) );
  CLKBUF_X3 U91321 ( .A(n81338), .Z(n106178) );
  NOR2_X1 U91322 ( .A1(n104994), .A2(n104705), .ZN(n104786) );
  AOI21_X1 U91323 ( .B1(n104899), .B2(n104495), .A(n100278), .ZN(n104787) );
  CLKBUF_X3 U91324 ( .A(n81275), .Z(n106251) );
  AND2_X2 U91325 ( .A1(n104788), .A2(n104921), .ZN(n82435) );
  CLKBUF_X3 U91326 ( .A(n81441), .Z(n106085) );
  NOR2_X1 U91327 ( .A1(n96557), .A2(n96558), .ZN(n104789) );
  NOR2_X1 U91328 ( .A1(n96557), .A2(n96558), .ZN(n104790) );
  CLKBUF_X3 U91329 ( .A(n81390), .Z(n106121) );
  AND2_X2 U91330 ( .A1(n105085), .A2(n104791), .ZN(n105025) );
  CLKBUF_X3 U91331 ( .A(n97579), .Z(n105335) );
  CLKBUF_X3 U91332 ( .A(n81356), .Z(n106152) );
  CLKBUF_X3 U91333 ( .A(n98618), .Z(n105243) );
  CLKBUF_X3 U91334 ( .A(n81355), .Z(n106154) );
  CLKBUF_X3 U91335 ( .A(n81369), .Z(n106143) );
  CLKBUF_X3 U91336 ( .A(n96561), .Z(n105130) );
  CLKBUF_X1 U91337 ( .A(n81899), .Z(n105031) );
  CLKBUF_X3 U91338 ( .A(n97715), .Z(n105315) );
  OR2_X1 U91339 ( .A1(n82301), .A2(n105153), .ZN(n104792) );
  INV_X1 U91340 ( .A(n104792), .ZN(n104793) );
  CLKBUF_X3 U91341 ( .A(n97899), .Z(n105297) );
  XNOR2_X1 U91342 ( .A(n104892), .B(n82387), .ZN(n82385) );
  CLKBUF_X3 U91343 ( .A(n106595), .Z(n105165) );
  AOI21_X1 U91344 ( .B1(n82377), .B2(n104795), .A(n104796), .ZN(n104794) );
  OR2_X1 U91345 ( .A1(n104793), .A2(n82259), .ZN(n82256) );
  OR2_X1 U91346 ( .A1(n105025), .A2(n105024), .ZN(n104797) );
  NAND2_X1 U91347 ( .A1(n104804), .A2(n104792), .ZN(n104799) );
  XOR2_X1 U91348 ( .A(n111132), .B(n104801), .Z(n104800) );
  INV_X1 U91349 ( .A(n104800), .ZN(n80137) );
  XOR2_X1 U91350 ( .A(n104758), .B(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_6/S_0 [1]), .Z(n104801) );
  OAI21_X1 U91351 ( .B1(n104916), .B2(n82223), .A(n82224), .ZN(n104802) );
  OR2_X1 U91352 ( .A1(n62182), .A2(n111154), .ZN(n104803) );
  NAND2_X1 U91353 ( .A1(n104803), .A2(n82408), .ZN(n82142) );
  OR2_X1 U91354 ( .A1(n105014), .A2(n82286), .ZN(n104805) );
  AND2_X2 U91355 ( .A1(n59518), .A2(n104806), .ZN(n100278) );
  NAND2_X1 U91356 ( .A1(\DLX_Datapath/CWP_IDEX[1] ), .A2(n105044), .ZN(n104806) );
  XNOR2_X1 U91357 ( .A(n104995), .B(n69347), .ZN(n100368) );
  XOR2_X1 U91358 ( .A(n104759), .B(n105153), .Z(n104807) );
  AND2_X2 U91359 ( .A1(net2465400), .A2(n111158), .ZN(n104808) );
  INV_X1 U91360 ( .A(n104808), .ZN(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_1/RCA_1/add_38_2/carry[1] ) );
  NOR2_X1 U91361 ( .A1(n82000), .A2(n81960), .ZN(n104809) );
  OAI21_X1 U91362 ( .B1(n104920), .B2(n105014), .A(net113102), .ZN(n104810) );
  CLKBUF_X1 U91363 ( .A(n82281), .Z(n104811) );
  NOR2_X1 U91364 ( .A1(n94808), .A2(n94553), .ZN(n104812) );
  NOR2_X1 U91365 ( .A1(n94808), .A2(n94553), .ZN(n104813) );
  XNOR2_X1 U91366 ( .A(n98941), .B(n104717), .ZN(n104815) );
  NOR2_X1 U91367 ( .A1(n95874), .A2(n95517), .ZN(n104816) );
  NOR2_X1 U91368 ( .A1(n96012), .A2(n96013), .ZN(n104819) );
  NOR2_X1 U91369 ( .A1(n96012), .A2(n96013), .ZN(n104820) );
  CLKBUF_X1 U91370 ( .A(n104910), .Z(n104821) );
  CLKBUF_X2 U91371 ( .A(n81325), .Z(n106181) );
  CLKBUF_X3 U91372 ( .A(n81325), .Z(n106182) );
  NOR2_X1 U91373 ( .A1(n95875), .A2(n105094), .ZN(n104822) );
  CLKBUF_X3 U91374 ( .A(n95518), .Z(n105495) );
  CLKBUF_X3 U91375 ( .A(n98438), .Z(n104823) );
  CLKBUF_X3 U91376 ( .A(n98578), .Z(n104825) );
  CLKBUF_X3 U91377 ( .A(n81479), .Z(n104827) );
  CLKBUF_X2 U91378 ( .A(n81479), .Z(n104828) );
  CLKBUF_X3 U91379 ( .A(n98372), .Z(n104829) );
  CLKBUF_X2 U91380 ( .A(n98372), .Z(n104830) );
  NOR2_X1 U91381 ( .A1(n82452), .A2(n104499), .ZN(n104831) );
  NAND2_X1 U91382 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [1]), 
        .A2(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [2]), .ZN(n104833)
         );
  CLKBUF_X1 U91383 ( .A(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_0/S_0[1] ), 
        .Z(PC_out[1]) );
  NOR2_X1 U91384 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_0/S_0[1] ), 
        .A2(PC_out[0]), .ZN(n104835) );
  CLKBUF_X3 U91385 ( .A(n98373), .Z(n105263) );
  CLKBUF_X2 U91386 ( .A(n98373), .Z(n105264) );
  NOR2_X1 U91387 ( .A1(n96392), .A2(n106757), .ZN(n104836) );
  CLKBUF_X1 U91388 ( .A(n105065), .Z(n104839) );
  CLKBUF_X3 U91389 ( .A(n81264), .Z(n106264) );
  CLKBUF_X3 U91390 ( .A(n98439), .Z(n105259) );
  CLKBUF_X3 U91391 ( .A(n98579), .Z(n105247) );
  CLKBUF_X3 U91392 ( .A(n95374), .Z(n105504) );
  NOR2_X1 U91393 ( .A1(n95837), .A2(n95555), .ZN(n104840) );
  NOR2_X1 U91394 ( .A1(n96012), .A2(n96013), .ZN(n104843) );
  CLKBUF_X2 U91395 ( .A(n81296), .Z(n106217) );
  NOR2_X1 U91396 ( .A1(n95556), .A2(n95555), .ZN(n104844) );
  CLKBUF_X3 U91397 ( .A(n97783), .Z(n105310) );
  NOR2_X1 U91398 ( .A1(net2465244), .A2(n111160), .ZN(n105071) );
  INV_X1 U91399 ( .A(n59517), .ZN(n104898) );
  NOR2_X1 U91400 ( .A1(n96053), .A2(n105091), .ZN(n104847) );
  CLKBUF_X3 U91401 ( .A(n95878), .Z(n105463) );
  INV_X1 U91402 ( .A(n105611), .ZN(n105609) );
  INV_X1 U91403 ( .A(n94626), .ZN(n105611) );
  CLKBUF_X3 U91404 ( .A(n81610), .Z(n104849) );
  CLKBUF_X2 U91405 ( .A(n81610), .Z(n104851) );
  CLKBUF_X3 U91406 ( .A(n81515), .Z(n104852) );
  CLKBUF_X3 U91407 ( .A(n81582), .Z(n104854) );
  CLKBUF_X3 U91408 ( .A(n94854), .Z(n105578) );
  CLKBUF_X1 U91409 ( .A(n106749), .Z(n104856) );
  CLKBUF_X3 U91410 ( .A(n97784), .Z(n105308) );
  CLKBUF_X3 U91411 ( .A(n98027), .Z(n105279) );
  CLKBUF_X3 U91412 ( .A(n97844), .Z(n105304) );
  CLKBUF_X1 U91413 ( .A(n82075), .Z(n104857) );
  CLKBUF_X3 U91414 ( .A(n96015), .Z(n105450) );
  CLKBUF_X3 U91415 ( .A(n96998), .Z(n104858) );
  CLKBUF_X3 U91416 ( .A(n97578), .Z(n105336) );
  CLKBUF_X3 U91417 ( .A(n96936), .Z(n104861) );
  CLKBUF_X2 U91418 ( .A(n96936), .Z(n104862) );
  CLKBUF_X3 U91419 ( .A(n97359), .Z(n104863) );
  CLKBUF_X3 U91420 ( .A(n97845), .Z(n105302) );
  XNOR2_X1 U91421 ( .A(n105049), .B(n99340), .ZN(n82691) );
  CLKBUF_X3 U91422 ( .A(n81611), .Z(n104865) );
  CLKBUF_X2 U91423 ( .A(n81611), .Z(n104867) );
  OR2_X1 U91424 ( .A1(n62196), .A2(net113081), .ZN(n104868) );
  CLKBUF_X3 U91425 ( .A(n97935), .Z(n105290) );
  CLKBUF_X3 U91426 ( .A(n98028), .Z(n105277) );
  CLKBUF_X3 U91427 ( .A(n97453), .Z(n104869) );
  NOR2_X1 U91428 ( .A1(n105004), .A2(n104878), .ZN(n104871) );
  CLKBUF_X3 U91429 ( .A(n81445), .Z(n106076) );
  CLKBUF_X3 U91430 ( .A(n81445), .Z(n106077) );
  CLKBUF_X3 U91431 ( .A(n96744), .Z(n104872) );
  CLKBUF_X2 U91432 ( .A(n64266), .Z(n104874) );
  CLKBUF_X3 U91433 ( .A(n97898), .Z(n105298) );
  CLKBUF_X3 U91434 ( .A(n94665), .Z(n105600) );
  CLKBUF_X3 U91435 ( .A(n97579), .Z(n105334) );
  CLKBUF_X3 U91436 ( .A(n97714), .Z(n105316) );
  CLKBUF_X3 U91437 ( .A(n95264), .Z(n105514) );
  CLKBUF_X3 U91438 ( .A(n96877), .Z(n105382) );
  CLKBUF_X3 U91439 ( .A(n96877), .Z(n105383) );
  NAND2_X1 U91440 ( .A1(n82426), .A2(n82427), .ZN(net113538) );
  NOR2_X1 U91441 ( .A1(n105004), .A2(n104878), .ZN(n98091) );
  CLKBUF_X3 U91442 ( .A(n97360), .Z(n105356) );
  CLKBUF_X3 U91443 ( .A(n81556), .Z(n106026) );
  CLKBUF_X3 U91444 ( .A(n81461), .Z(n106066) );
  CLKBUF_X3 U91445 ( .A(n81461), .Z(n106065) );
  CLKBUF_X3 U91446 ( .A(n97395), .Z(n105352) );
  CLKBUF_X3 U91447 ( .A(n96683), .Z(n105405) );
  CLKBUF_X3 U91448 ( .A(n97715), .Z(n105314) );
  CLKBUF_X3 U91449 ( .A(n81390), .Z(n106120) );
  CLKBUF_X3 U91450 ( .A(n81462), .Z(n106063) );
  CLKBUF_X3 U91451 ( .A(n81446), .Z(n106074) );
  CLKBUF_X3 U91452 ( .A(n97899), .Z(n105296) );
  CLKBUF_X3 U91453 ( .A(n81355), .Z(n106153) );
  CLKBUF_X3 U91454 ( .A(n106749), .Z(n105177) );
  CLKBUF_X3 U91455 ( .A(n81369), .Z(n106142) );
  CLKBUF_X3 U91456 ( .A(n98543), .Z(n105251) );
  CLKBUF_X3 U91457 ( .A(n98543), .Z(n105252) );
  CLKBUF_X3 U91458 ( .A(n81326), .Z(n104881) );
  CLKBUF_X3 U91459 ( .A(n81543), .Z(n106029) );
  CLKBUF_X3 U91460 ( .A(n81543), .Z(n106031) );
  CLKBUF_X3 U91461 ( .A(n98505), .Z(n105255) );
  CLKBUF_X3 U91462 ( .A(n98542), .Z(n104883) );
  CLKBUF_X2 U91463 ( .A(n98542), .Z(n104884) );
  CLKBUF_X3 U91464 ( .A(n98504), .Z(n104885) );
  CLKBUF_X3 U91465 ( .A(n81338), .Z(n106177) );
  NOR2_X1 U91466 ( .A1(n111132), .A2(n57427), .ZN(n104887) );
  CLKBUF_X2 U91467 ( .A(n81566), .Z(n106023) );
  CLKBUF_X3 U91468 ( .A(n81566), .Z(n106024) );
  CLKBUF_X3 U91469 ( .A(n81356), .Z(n106151) );
  CLKBUF_X3 U91470 ( .A(n96804), .Z(n105394) );
  CLKBUF_X3 U91471 ( .A(n81276), .Z(n106248) );
  CLKBUF_X3 U91472 ( .A(n81309), .Z(n106202) );
  CLKBUF_X3 U91473 ( .A(n97514), .Z(n105342) );
  CLKBUF_X3 U91474 ( .A(n97935), .Z(n105291) );
  CLKBUF_X3 U91475 ( .A(n96841), .Z(n105388) );
  NAND2_X1 U91476 ( .A1(n82384), .A2(n104891), .ZN(n82187) );
  OAI21_X1 U91477 ( .B1(n106780), .B2(n82388), .A(n82389), .ZN(n104892) );
  CLKBUF_X3 U91478 ( .A(n97323), .Z(n105360) );
  CLKBUF_X3 U91479 ( .A(n97322), .Z(n105362) );
  INV_X1 U91480 ( .A(n104904), .ZN(n94295) );
  CLKBUF_X3 U91481 ( .A(n81516), .Z(n106040) );
  CLKBUF_X3 U91482 ( .A(n96805), .Z(n105393) );
  CLKBUF_X3 U91483 ( .A(n96999), .Z(n105371) );
  CLKBUF_X3 U91484 ( .A(n97515), .Z(n105341) );
  CLKBUF_X3 U91485 ( .A(n96842), .Z(n105387) );
  OR2_X1 U91486 ( .A1(n106770), .A2(n104894), .ZN(n82657) );
  CLKBUF_X3 U91487 ( .A(n81528), .Z(n106035) );
  CLKBUF_X3 U91488 ( .A(n81528), .Z(n106036) );
  CLKBUF_X3 U91489 ( .A(n97454), .Z(n105346) );
  CLKBUF_X3 U91490 ( .A(n96745), .Z(n105398) );
  CLKBUF_X3 U91491 ( .A(n97641), .Z(n105327) );
  CLKBUF_X3 U91492 ( .A(n97641), .Z(n105328) );
  CLKBUF_X3 U91493 ( .A(n106758), .Z(n105188) );
  CLKBUF_X2 U91494 ( .A(n106758), .Z(n105189) );
  CLKBUF_X3 U91495 ( .A(n97677), .Z(n105323) );
  CLKBUF_X3 U91496 ( .A(n97677), .Z(n105324) );
  CLKBUF_X2 U91497 ( .A(n97677), .Z(n105325) );
  CLKBUF_X3 U91498 ( .A(n96684), .Z(n105402) );
  CLKBUF_X3 U91499 ( .A(n96684), .Z(n105403) );
  CLKBUF_X3 U91500 ( .A(n81387), .Z(n106124) );
  CLKBUF_X2 U91501 ( .A(n81442), .Z(n106081) );
  CLKBUF_X3 U91502 ( .A(n81442), .Z(n106080) );
  CLKBUF_X3 U91503 ( .A(n81442), .Z(n106082) );
  NOR2_X1 U91504 ( .A1(n82316), .A2(n104897), .ZN(n104895) );
  NOR2_X1 U91505 ( .A1(n104895), .A2(n104896), .ZN(n104914) );
  OR2_X1 U91506 ( .A1(n104505), .A2(n82200), .ZN(n104897) );
  NOR2_X1 U91507 ( .A1(n104510), .A2(net71745), .ZN(n82316) );
  CLKBUF_X2 U91508 ( .A(n81760), .Z(n105919) );
  CLKBUF_X3 U91509 ( .A(n81760), .Z(n105920) );
  CLKBUF_X3 U91510 ( .A(n81583), .Z(n106014) );
  CLKBUF_X3 U91511 ( .A(n95803), .Z(n105472) );
  CLKBUF_X2 U91512 ( .A(n95803), .Z(n105473) );
  CLKBUF_X3 U91513 ( .A(n81291), .Z(n106225) );
  AND2_X2 U91514 ( .A1(n59516), .A2(n107106), .ZN(n100382) );
  CLKBUF_X3 U91515 ( .A(n81516), .Z(n106039) );
  AND2_X2 U91516 ( .A1(n105077), .A2(\DLX_Datapath/CWP_IDEX[2] ), .ZN(n104899)
         );
  INV_X1 U91517 ( .A(n104899), .ZN(n100276) );
  AND4_X4 U91518 ( .A1(n104901), .A2(n104900), .A3(n104848), .A4(n104902), 
        .ZN(n82681) );
  XNOR2_X1 U91519 ( .A(n82688), .B(n82689), .ZN(n104901) );
  XNOR2_X1 U91520 ( .A(n100419), .B(n59452), .ZN(n104902) );
  XOR2_X1 U91521 ( .A(n104903), .B(n104741), .Z(n100363) );
  CLKBUF_X3 U91522 ( .A(n95915), .Z(n105458) );
  CLKBUF_X3 U91523 ( .A(n96358), .Z(n105419) );
  CLKBUF_X3 U91524 ( .A(n95841), .Z(n105469) );
  CLKBUF_X3 U91525 ( .A(n95841), .Z(n105468) );
  CLKBUF_X3 U91526 ( .A(n105030), .Z(n105051) );
  CLKBUF_X3 U91527 ( .A(n81568), .Z(n106018) );
  CLKBUF_X3 U91528 ( .A(n81568), .Z(n106017) );
  OAI21_X1 U91529 ( .B1(n104757), .B2(n94893), .A(n69424), .ZN(n104904) );
  CLKBUF_X3 U91530 ( .A(n95521), .Z(n105494) );
  NAND2_X1 U91531 ( .A1(n104905), .A2(n104906), .ZN(n82458) );
  NOR2_X1 U91532 ( .A1(n82452), .A2(n104499), .ZN(n104905) );
  NOR2_X1 U91533 ( .A1(n62194), .A2(n104494), .ZN(n104906) );
  CLKBUF_X1 U91534 ( .A(n106769), .Z(n104907) );
  INV_X1 U91535 ( .A(net73629), .ZN(net113081) );
  INV_X1 U91536 ( .A(net113156), .ZN(net113091) );
  INV_X1 U91537 ( .A(net113154), .ZN(net113102) );
  INV_X1 U91538 ( .A(n80001), .ZN(net113152) );
  INV_X1 U91539 ( .A(n80001), .ZN(net113153) );
  INV_X1 U91540 ( .A(net113152), .ZN(net113156) );
  INV_X1 U91541 ( .A(n90137), .ZN(n107128) );
  AND2_X2 U91542 ( .A1(n105135), .A2(n94093), .ZN(n104908) );
  AND2_X2 U91543 ( .A1(n105135), .A2(n94093), .ZN(n104909) );
  INV_X1 U91544 ( .A(n104821), .ZN(n82613) );
  OR2_X1 U91545 ( .A1(n104802), .A2(n82218), .ZN(n104911) );
  NAND2_X1 U91546 ( .A1(n82219), .A2(n104911), .ZN(n80148) );
  XNOR2_X1 U91547 ( .A(n104915), .B(n57431), .ZN(n82284) );
  CLKBUF_X3 U91548 ( .A(n82021), .Z(n105897) );
  OR2_X1 U91549 ( .A1(n105025), .A2(n105024), .ZN(n104916) );
  INV_X1 U91550 ( .A(n104916), .ZN(n105020) );
  OR2_X1 U91551 ( .A1(n105025), .A2(n104917), .ZN(n105019) );
  NAND2_X1 U91552 ( .A1(n105040), .A2(n105043), .ZN(n104917) );
  OR2_X1 U91553 ( .A1(n82301), .A2(n105153), .ZN(n104918) );
  OR2_X1 U91554 ( .A1(n82654), .A2(n82653), .ZN(n104920) );
  OAI21_X1 U91555 ( .B1(n81922), .B2(net113157), .A(n80104), .ZN(n104921) );
  INV_X1 U91556 ( .A(n104921), .ZN(n105017) );
  XNOR2_X1 U91557 ( .A(n82256), .B(n104509), .ZN(n80150) );
  AND2_X2 U91558 ( .A1(n105035), .A2(n94081), .ZN(n104922) );
  INV_X1 U91559 ( .A(n104757), .ZN(n94093) );
  INV_X1 U91560 ( .A(n94895), .ZN(n105004) );
  NOR2_X1 U91561 ( .A1(n104763), .A2(n104798), .ZN(n82301) );
  CLKBUF_X3 U91562 ( .A(n98304), .Z(n105267) );
  CLKBUF_X3 U91563 ( .A(n97934), .Z(n105292) );
  CLKBUF_X2 U91564 ( .A(n97934), .Z(n105293) );
  AND2_X2 U91565 ( .A1(n105136), .A2(n94853), .ZN(n104923) );
  CLKBUF_X3 U91566 ( .A(n96234), .Z(n104924) );
  CLKBUF_X2 U91567 ( .A(n96234), .Z(n104925) );
  CLKBUF_X3 U91568 ( .A(n94856), .Z(n105577) );
  CLKBUF_X3 U91569 ( .A(n81296), .Z(n106216) );
  CLKBUF_X3 U91570 ( .A(n81649), .Z(n104930) );
  CLKBUF_X3 U91571 ( .A(n81596), .Z(n106003) );
  CLKBUF_X3 U91572 ( .A(n81596), .Z(n106004) );
  CLKBUF_X3 U91573 ( .A(n81596), .Z(n106005) );
  CLKBUF_X3 U91574 ( .A(n95655), .Z(n104939) );
  CLKBUF_X2 U91575 ( .A(n95655), .Z(n104940) );
  CLKBUF_X3 U91576 ( .A(n94668), .Z(n105003) );
  CLKBUF_X2 U91577 ( .A(n81597), .Z(n104941) );
  CLKBUF_X3 U91578 ( .A(n81597), .Z(n104942) );
  CLKBUF_X3 U91579 ( .A(n81597), .Z(n104943) );
  CLKBUF_X1 U91580 ( .A(n81597), .Z(n104944) );
  CLKBUF_X1 U91581 ( .A(n81597), .Z(n104945) );
  CLKBUF_X1 U91582 ( .A(n81597), .Z(n104946) );
  CLKBUF_X3 U91583 ( .A(n95729), .Z(n104948) );
  CLKBUF_X3 U91584 ( .A(n95376), .Z(n104951) );
  CLKBUF_X3 U91585 ( .A(n81691), .Z(n104954) );
  CLKBUF_X3 U91586 ( .A(n81691), .Z(n104955) );
  CLKBUF_X3 U91587 ( .A(n81339), .Z(n106175) );
  CLKBUF_X3 U91588 ( .A(n95455), .Z(n105497) );
  CLKBUF_X3 U91589 ( .A(n95455), .Z(n105496) );
  CLKBUF_X3 U91590 ( .A(n95589), .Z(n105489) );
  CLKBUF_X3 U91591 ( .A(n81291), .Z(n106224) );
  CLKBUF_X3 U91592 ( .A(n81683), .Z(n104962) );
  CLKBUF_X3 U91593 ( .A(n81683), .Z(n104963) );
  CLKBUF_X3 U91594 ( .A(n81683), .Z(n104964) );
  CLKBUF_X3 U91595 ( .A(n95955), .Z(n104965) );
  CLKBUF_X2 U91596 ( .A(n95955), .Z(n104966) );
  CLKBUF_X3 U91597 ( .A(n96493), .Z(n104967) );
  CLKBUF_X2 U91598 ( .A(n96493), .Z(n104968) );
  CLKBUF_X3 U91599 ( .A(n95590), .Z(n104972) );
  CLKBUF_X2 U91600 ( .A(n81735), .Z(n105935) );
  CLKBUF_X3 U91601 ( .A(n81660), .Z(n105964) );
  CLKBUF_X3 U91602 ( .A(n95415), .Z(n104980) );
  CLKBUF_X3 U91603 ( .A(n95415), .Z(n104981) );
  CLKBUF_X3 U91604 ( .A(n94333), .Z(n104983) );
  CLKBUF_X3 U91605 ( .A(n81275), .Z(n106250) );
  CLKBUF_X3 U91606 ( .A(n94472), .Z(n104985) );
  CLKBUF_X3 U91607 ( .A(n96133), .Z(n104987) );
  CLKBUF_X3 U91608 ( .A(n96133), .Z(n104988) );
  NAND2_X1 U91609 ( .A1(n104908), .A2(n94367), .ZN(n104992) );
  CLKBUF_X3 U91610 ( .A(n81777), .Z(n105915) );
  CLKBUF_X3 U91611 ( .A(n81777), .Z(n105916) );
  NAND2_X1 U91612 ( .A1(n104909), .A2(n94367), .ZN(n104993) );
  CLKBUF_X1 U91613 ( .A(n107104), .Z(n104996) );
  CLKBUF_X1 U91614 ( .A(n94257), .Z(n104997) );
  CLKBUF_X3 U91615 ( .A(n95266), .Z(n104998) );
  CLKBUF_X3 U91616 ( .A(n81776), .Z(n105000) );
  CLKBUF_X3 U91617 ( .A(n81776), .Z(n105001) );
  INV_X1 U91618 ( .A(n94506), .ZN(n105631) );
  CLKBUF_X3 U91619 ( .A(n94668), .Z(n105002) );
  AND2_X2 U91620 ( .A1(n105005), .A2(n105004), .ZN(n98654) );
  AND2_X2 U91621 ( .A1(n104815), .A2(n95412), .ZN(n105005) );
  CLKBUF_X3 U91622 ( .A(n81290), .Z(n106227) );
  CLKBUF_X3 U91623 ( .A(n81290), .Z(n106228) );
  CLKBUF_X3 U91624 ( .A(n82027), .Z(n105892) );
  CLKBUF_X3 U91625 ( .A(n82021), .Z(n105896) );
  OR2_X1 U91626 ( .A1(n111063), .A2(n105585), .ZN(n105006) );
  NAND2_X1 U91627 ( .A1(n94839), .A2(n105006), .ZN(
        \DLX_Datapath/RegisterFile/N26417 ) );
  OR2_X1 U91628 ( .A1(n107394), .A2(n105585), .ZN(n105007) );
  NAND2_X1 U91629 ( .A1(n94826), .A2(n105007), .ZN(
        \DLX_Datapath/RegisterFile/N26430 ) );
  OR2_X1 U91630 ( .A1(n107369), .A2(n105585), .ZN(n105008) );
  NAND2_X1 U91631 ( .A1(n94837), .A2(n105008), .ZN(
        \DLX_Datapath/RegisterFile/N26419 ) );
  OR2_X1 U91632 ( .A1(n107390), .A2(n105585), .ZN(n105009) );
  NAND2_X1 U91633 ( .A1(n94824), .A2(n105009), .ZN(
        \DLX_Datapath/RegisterFile/N26432 ) );
  CLKBUF_X3 U91634 ( .A(n81441), .Z(n106083) );
  CLKBUF_X3 U91635 ( .A(n81441), .Z(n106084) );
  OR2_X1 U91636 ( .A1(n107367), .A2(n105585), .ZN(n105010) );
  NAND2_X1 U91637 ( .A1(n94836), .A2(n105010), .ZN(
        \DLX_Datapath/RegisterFile/N26420 ) );
  INV_X1 U91638 ( .A(n94735), .ZN(n105011) );
  INV_X1 U91639 ( .A(n105011), .ZN(n105598) );
  CLKBUF_X3 U91640 ( .A(n96358), .Z(n105418) );
  INV_X2 U91641 ( .A(n105591), .ZN(n105590) );
  CLKBUF_X3 U91642 ( .A(n95076), .Z(n105540) );
  CLKBUF_X3 U91643 ( .A(n95076), .Z(n105541) );
  CLKBUF_X3 U91644 ( .A(n94937), .Z(n105561) );
  CLKBUF_X3 U91645 ( .A(n94937), .Z(n105562) );
  CLKBUF_X3 U91646 ( .A(n95040), .Z(n105549) );
  CLKBUF_X3 U91647 ( .A(n95040), .Z(n105550) );
  CLKBUF_X2 U91648 ( .A(n95040), .Z(n105551) );
  CLKBUF_X3 U91649 ( .A(n94899), .Z(n105567) );
  CLKBUF_X3 U91650 ( .A(n106750), .Z(n105178) );
  CLKBUF_X2 U91651 ( .A(n106750), .Z(n105179) );
  CLKBUF_X3 U91652 ( .A(n95521), .Z(n105493) );
  CLKBUF_X3 U91653 ( .A(n96017), .Z(n105448) );
  CLKBUF_X1 U91654 ( .A(n59517), .Z(n105012) );
  CLKBUF_X3 U91655 ( .A(n95077), .Z(n105537) );
  CLKBUF_X3 U91656 ( .A(n95077), .Z(n105538) );
  CLKBUF_X3 U91657 ( .A(n94938), .Z(n105558) );
  CLKBUF_X3 U91658 ( .A(n94938), .Z(n105559) );
  CLKBUF_X3 U91659 ( .A(n106756), .Z(n105187) );
  CLKBUF_X3 U91660 ( .A(n79979), .Z(n106351) );
  AND4_X4 U91661 ( .A1(n81981), .A2(IR_in[1]), .A3(net112601), .A4(net67007), 
        .ZN(n81996) );
  CLKBUF_X3 U91662 ( .A(n94814), .Z(n105581) );
  CLKBUF_X3 U91663 ( .A(n95654), .Z(n105485) );
  CLKBUF_X3 U91664 ( .A(n95654), .Z(n105486) );
  CLKBUF_X3 U91665 ( .A(n81690), .Z(n105948) );
  CLKBUF_X3 U91666 ( .A(n95878), .Z(n105461) );
  CLKBUF_X3 U91667 ( .A(n95878), .Z(n105462) );
  AND2_X2 U91668 ( .A1(n104785), .A2(n82276), .ZN(n105013) );
  INV_X1 U91669 ( .A(n105013), .ZN(n82019) );
  CLKBUF_X3 U91670 ( .A(n94898), .Z(n105570) );
  CLKBUF_X3 U91671 ( .A(n94898), .Z(n105571) );
  CLKBUF_X3 U91672 ( .A(n80152), .Z(n106343) );
  CLKBUF_X3 U91673 ( .A(n80152), .Z(n106344) );
  CLKBUF_X3 U91674 ( .A(n95041), .Z(n105546) );
  CLKBUF_X3 U91675 ( .A(n95041), .Z(n105547) );
  CLKBUF_X3 U91676 ( .A(n94856), .Z(n105576) );
  CLKBUF_X3 U91677 ( .A(n82027), .Z(n105891) );
  CLKBUF_X3 U91678 ( .A(n79970), .Z(n106354) );
  CLKBUF_X3 U91679 ( .A(n79979), .Z(n106350) );
  CLKBUF_X3 U91680 ( .A(n104699), .Z(n105159) );
  CLKBUF_X3 U91681 ( .A(n106755), .Z(n105184) );
  CLKBUF_X3 U91682 ( .A(n106755), .Z(n105185) );
  CLKBUF_X3 U91683 ( .A(n104699), .Z(n105158) );
  OR2_X1 U91684 ( .A1(n57431), .A2(net113081), .ZN(n105015) );
  NAND2_X1 U91685 ( .A1(n82275), .A2(n105015), .ZN(n82274) );
  AND2_X2 U91686 ( .A1(n105044), .A2(\DLX_Datapath/CWP_IDEX[1] ), .ZN(n105077)
         );
  CLKBUF_X3 U91687 ( .A(n105013), .Z(n105157) );
  CLKBUF_X3 U91688 ( .A(n104919), .Z(n105895) );
  OR2_X1 U91689 ( .A1(n107390), .A2(n104992), .ZN(n105016) );
  NAND2_X1 U91690 ( .A1(n105016), .A2(n95012), .ZN(
        \DLX_Datapath/RegisterFile/N26272 ) );
  CLKBUF_X3 U91691 ( .A(n79970), .Z(n106355) );
  CLKBUF_X3 U91692 ( .A(n82435), .Z(n105888) );
  CLKBUF_X3 U91693 ( .A(n106756), .Z(n105186) );
  CLKBUF_X3 U91694 ( .A(n106752), .Z(n105039) );
  CLKBUF_X3 U91695 ( .A(n106752), .Z(n105182) );
  CLKBUF_X3 U91696 ( .A(n106751), .Z(n105047) );
  CLKBUF_X3 U91697 ( .A(n106751), .Z(n105181) );
  NAND2_X1 U91698 ( .A1(net112383), .A2(IR_in[6]), .ZN(net112469) );
  CLKBUF_X3 U91699 ( .A(n94814), .Z(n105579) );
  CLKBUF_X3 U91700 ( .A(n94814), .Z(n105580) );
  CLKBUF_X3 U91701 ( .A(n105013), .Z(n105156) );
  CLKBUF_X3 U91702 ( .A(n104919), .Z(n105894) );
  NOR2_X1 U91703 ( .A1(n82316), .A2(n104505), .ZN(n82314) );
  NOR3_X1 U91704 ( .A1(n82311), .A2(n82313), .A3(n82312), .ZN(n105021) );
  INV_X1 U91705 ( .A(n105021), .ZN(n105022) );
  INV_X1 U91706 ( .A(n105043), .ZN(n105024) );
  NOR2_X1 U91707 ( .A1(n100367), .A2(n104524), .ZN(n100354) );
  CLKBUF_X3 U91708 ( .A(n82435), .Z(n105887) );
  INV_X1 U91709 ( .A(n104907), .ZN(n105023) );
  XNOR2_X1 U91710 ( .A(n104784), .B(n105153), .ZN(n80124) );
  XNOR2_X1 U91711 ( .A(n82269), .B(n105027), .ZN(n105026) );
  INV_X1 U91712 ( .A(n105026), .ZN(n80125) );
  INV_X1 U91713 ( .A(n105036), .ZN(n105028) );
  INV_X1 U91714 ( .A(n98942), .ZN(n105036) );
  AOI21_X1 U91715 ( .B1(n90137), .B2(n107131), .A(n104922), .ZN(n105029) );
  NOR2_X1 U91716 ( .A1(n104805), .A2(n105151), .ZN(n105030) );
  OR2_X1 U91717 ( .A1(IR_in[5]), .A2(
        \DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_1/S_0 [1]), .ZN(net112383) );
  NOR2_X1 U91718 ( .A1(n82468), .A2(n57425), .ZN(n105033) );
  CLKBUF_X1 U91719 ( .A(n62664), .Z(n105034) );
  CLKBUF_X1 U91720 ( .A(n106752), .Z(n105038) );
  OR2_X1 U91721 ( .A1(n59477), .A2(n82303), .ZN(n105040) );
  INV_X1 U91722 ( .A(net112358), .ZN(net112354) );
  INV_X1 U91723 ( .A(n82292), .ZN(n105041) );
  NOR3_X1 U91724 ( .A1(n104511), .A2(n100359), .A3(n100358), .ZN(n100355) );
  NAND2_X1 U91725 ( .A1(n105042), .A2(n100381), .ZN(n94257) );
  OR2_X1 U91726 ( .A1(n82304), .A2(n62191), .ZN(n105043) );
  CLKBUF_X1 U91727 ( .A(n106751), .Z(n105046) );
  NAND2_X1 U91728 ( .A1(n105048), .A2(n105059), .ZN(n98942) );
  NOR2_X1 U91729 ( .A1(n104721), .A2(n104720), .ZN(n105049) );
  NOR2_X1 U91730 ( .A1(n59517), .A2(n59516), .ZN(n105052) );
  CLKBUF_X1 U91731 ( .A(n106741), .Z(n105169) );
  CLKBUF_X1 U91732 ( .A(n81261), .Z(n106271) );
  CLKBUF_X1 U91733 ( .A(n107127), .Z(n105215) );
  CLKBUF_X1 U91734 ( .A(n107127), .Z(n105216) );
  CLKBUF_X1 U91735 ( .A(n107127), .Z(n105217) );
  CLKBUF_X1 U91736 ( .A(n107127), .Z(n105218) );
  CLKBUF_X1 U91737 ( .A(n107127), .Z(n105219) );
  CLKBUF_X1 U91738 ( .A(n107127), .Z(n105220) );
  CLKBUF_X1 U91739 ( .A(n107116), .Z(n105212) );
  CLKBUF_X1 U91740 ( .A(n107116), .Z(n105211) );
  CLKBUF_X1 U91741 ( .A(n107117), .Z(n105214) );
  CLKBUF_X1 U91742 ( .A(n107115), .Z(n105210) );
  CLKBUF_X1 U91743 ( .A(n107115), .Z(n105209) );
  CLKBUF_X1 U91744 ( .A(n107117), .Z(n105213) );
  CLKBUF_X1 U91745 ( .A(n81353), .Z(n106155) );
  CLKBUF_X2 U91746 ( .A(n95952), .Z(n105454) );
  CLKBUF_X1 U91747 ( .A(n106760), .Z(n105193) );
  CLKBUF_X1 U91748 ( .A(n106760), .Z(n105192) );
  CLKBUF_X1 U91749 ( .A(n106759), .Z(n105190) );
  CLKBUF_X1 U91750 ( .A(n81733), .Z(n105936) );
  CLKBUF_X1 U91751 ( .A(n96418), .Z(n105417) );
  CLKBUF_X1 U91752 ( .A(n95875), .Z(n105467) );
  CLKBUF_X1 U91753 ( .A(n95690), .Z(n105484) );
  CLKBUF_X1 U91754 ( .A(n81443), .Z(n106078) );
  CLKBUF_X1 U91755 ( .A(n97451), .Z(n105348) );
  CLKBUF_X1 U91756 ( .A(n81526), .Z(n106038) );
  CLKBUF_X1 U91757 ( .A(n96934), .Z(n105378) );
  CLKBUF_X1 U91758 ( .A(n98502), .Z(n105257) );
  CLKBUF_X1 U91759 ( .A(n97969), .Z(n105289) );
  CLKBUF_X1 U91760 ( .A(n97512), .Z(n105345) );
  CLKBUF_X1 U91761 ( .A(n96996), .Z(n105373) );
  CLKBUF_X1 U91762 ( .A(n98576), .Z(n105249) );
  CLKBUF_X1 U91763 ( .A(n98025), .Z(n105281) );
  CLKBUF_X1 U91764 ( .A(n81261), .Z(n106272) );
  CLKBUF_X1 U91765 ( .A(n81443), .Z(n106079) );
  CLKBUF_X1 U91766 ( .A(n97451), .Z(n105349) );
  CLKBUF_X1 U91767 ( .A(n81353), .Z(n106156) );
  CLKBUF_X1 U91768 ( .A(n98502), .Z(n105258) );
  CLKBUF_X1 U91769 ( .A(n96996), .Z(n105374) );
  CLKBUF_X1 U91770 ( .A(n98576), .Z(n105250) );
  CLKBUF_X1 U91771 ( .A(n98025), .Z(n105282) );
  CLKBUF_X1 U91772 ( .A(n96017), .Z(n105449) );
  CLKBUF_X1 U91773 ( .A(n106760), .Z(n105194) );
  CLKBUF_X1 U91774 ( .A(n106759), .Z(n105191) );
  INV_X1 U91775 ( .A(n105864), .ZN(n105863) );
  INV_X1 U91776 ( .A(n106279), .ZN(n106278) );
  CLKBUF_X1 U91777 ( .A(n84160), .Z(n105826) );
  CLKBUF_X1 U91778 ( .A(n85252), .Z(n105807) );
  CLKBUF_X1 U91779 ( .A(n83149), .Z(n105870) );
  CLKBUF_X1 U91780 ( .A(n85217), .Z(n105824) );
  CLKBUF_X1 U91781 ( .A(n106945), .Z(n105196) );
  CLKBUF_X1 U91782 ( .A(n84157), .Z(n105828) );
  CLKBUF_X1 U91783 ( .A(n85257), .Z(n105803) );
  CLKBUF_X1 U91784 ( .A(n80217), .Z(n106316) );
  CLKBUF_X1 U91785 ( .A(n80253), .Z(n106295) );
  CLKBUF_X1 U91786 ( .A(n84161), .Z(n105825) );
  CLKBUF_X1 U91787 ( .A(n85259), .Z(n105801) );
  CLKBUF_X1 U91788 ( .A(n84132), .Z(n105843) );
  CLKBUF_X1 U91789 ( .A(n84150), .Z(n105833) );
  CLKBUF_X1 U91790 ( .A(n83143), .Z(n105872) );
  CLKBUF_X1 U91791 ( .A(n106739), .Z(n105168) );
  CLKBUF_X1 U91792 ( .A(n84126), .Z(n105848) );
  CLKBUF_X1 U91793 ( .A(n80255), .Z(n106293) );
  CLKBUF_X1 U91794 ( .A(n84127), .Z(n105847) );
  CLKBUF_X1 U91795 ( .A(n84146), .Z(n105836) );
  INV_X1 U91796 ( .A(n83256), .ZN(n106741) );
  CLKBUF_X1 U91797 ( .A(n106738), .Z(n105167) );
  INV_X1 U91798 ( .A(n106012), .ZN(n106011) );
  INV_X1 U91799 ( .A(n106012), .ZN(n106010) );
  INV_X1 U91800 ( .A(n106012), .ZN(n106008) );
  INV_X1 U91801 ( .A(n105993), .ZN(n105992) );
  INV_X1 U91802 ( .A(n105993), .ZN(n105991) );
  INV_X1 U91803 ( .A(n105993), .ZN(n105990) );
  INV_X1 U91804 ( .A(n106258), .ZN(n106257) );
  INV_X1 U91805 ( .A(n106258), .ZN(n106256) );
  INV_X1 U91806 ( .A(n106258), .ZN(n106255) );
  INV_X1 U91807 ( .A(n106258), .ZN(n106254) );
  INV_X1 U91808 ( .A(n106207), .ZN(n106206) );
  INV_X1 U91809 ( .A(n106207), .ZN(n106205) );
  INV_X1 U91810 ( .A(n106207), .ZN(n106204) );
  INV_X1 U91811 ( .A(n106207), .ZN(n106203) );
  INV_X1 U91812 ( .A(n106102), .ZN(n106101) );
  INV_X1 U91813 ( .A(n106102), .ZN(n106100) );
  INV_X1 U91814 ( .A(n106102), .ZN(n106099) );
  INV_X1 U91815 ( .A(n106102), .ZN(n106098) );
  INV_X1 U91816 ( .A(n105972), .ZN(n105971) );
  INV_X1 U91817 ( .A(n105972), .ZN(n105970) );
  INV_X1 U91818 ( .A(n105972), .ZN(n105969) );
  INV_X1 U91819 ( .A(n105972), .ZN(n105968) );
  INV_X1 U91820 ( .A(n106150), .ZN(n106149) );
  INV_X1 U91821 ( .A(n106150), .ZN(n106148) );
  INV_X1 U91822 ( .A(n106150), .ZN(n106147) );
  INV_X1 U91823 ( .A(n106150), .ZN(n106146) );
  INV_X1 U91824 ( .A(n106212), .ZN(n106211) );
  INV_X1 U91825 ( .A(n106212), .ZN(n106210) );
  INV_X1 U91826 ( .A(n106212), .ZN(n106209) );
  INV_X1 U91827 ( .A(n106212), .ZN(n106208) );
  INV_X1 U91828 ( .A(n106139), .ZN(n106138) );
  INV_X1 U91829 ( .A(n106139), .ZN(n106137) );
  INV_X1 U91830 ( .A(n106139), .ZN(n106136) );
  INV_X1 U91831 ( .A(n106139), .ZN(n106135) );
  INV_X1 U91832 ( .A(n105554), .ZN(n105552) );
  INV_X1 U91833 ( .A(n105954), .ZN(n105953) );
  INV_X1 U91834 ( .A(n105954), .ZN(n105952) );
  INV_X1 U91835 ( .A(n105566), .ZN(n105565) );
  INV_X1 U91836 ( .A(n105545), .ZN(n105544) );
  INV_X1 U91837 ( .A(n105545), .ZN(n105543) );
  INV_X1 U91838 ( .A(n105566), .ZN(n105564) );
  INV_X1 U91839 ( .A(n105951), .ZN(n105950) );
  INV_X1 U91840 ( .A(n105951), .ZN(n105949) );
  INV_X1 U91841 ( .A(n105575), .ZN(n105574) );
  INV_X1 U91842 ( .A(n105575), .ZN(n105573) );
  INV_X1 U91843 ( .A(n105611), .ZN(n105610) );
  INV_X1 U91844 ( .A(n105631), .ZN(n105629) );
  INV_X1 U91845 ( .A(n105620), .ZN(n105618) );
  INV_X1 U91846 ( .A(n104923), .ZN(n105585) );
  INV_X1 U91847 ( .A(n105903), .ZN(n105901) );
  INV_X1 U91848 ( .A(n105903), .ZN(n105902) );
  INV_X1 U91849 ( .A(n105631), .ZN(n105630) );
  INV_X1 U91850 ( .A(n105011), .ZN(n105599) );
  INV_X1 U91851 ( .A(n105620), .ZN(n105619) );
  INV_X1 U91852 ( .A(n104923), .ZN(n105586) );
  CLKBUF_X1 U91853 ( .A(n105199), .Z(n105203) );
  CLKBUF_X1 U91854 ( .A(n105199), .Z(n105200) );
  CLKBUF_X1 U91855 ( .A(n105199), .Z(n105202) );
  CLKBUF_X1 U91856 ( .A(n105199), .Z(n105201) );
  CLKBUF_X1 U91857 ( .A(n94737), .Z(n105595) );
  CLKBUF_X1 U91858 ( .A(n94737), .Z(n105596) );
  CLKBUF_X1 U91859 ( .A(n105199), .Z(n105204) );
  CLKBUF_X1 U91860 ( .A(n81784), .Z(n105908) );
  CLKBUF_X1 U91861 ( .A(n81668), .Z(n105958) );
  CLKBUF_X1 U91862 ( .A(n94558), .Z(n105615) );
  CLKBUF_X1 U91863 ( .A(n94558), .Z(n105616) );
  CLKBUF_X1 U91864 ( .A(n94628), .Z(n105606) );
  CLKBUF_X1 U91865 ( .A(n94628), .Z(n105607) );
  CLKBUF_X1 U91866 ( .A(n94775), .Z(n105587) );
  CLKBUF_X1 U91867 ( .A(n94775), .Z(n105588) );
  CLKBUF_X1 U91868 ( .A(n94813), .Z(n105582) );
  CLKBUF_X1 U91869 ( .A(n94813), .Z(n105583) );
  CLKBUF_X1 U91870 ( .A(n95209), .Z(n105519) );
  CLKBUF_X1 U91871 ( .A(n95209), .Z(n105518) );
  CLKBUF_X1 U91872 ( .A(n81668), .Z(n105959) );
  CLKBUF_X1 U91873 ( .A(n81784), .Z(n105909) );
  CLKBUF_X1 U91874 ( .A(n95334), .Z(n105509) );
  CLKBUF_X1 U91875 ( .A(n95334), .Z(n105508) );
  CLKBUF_X1 U91876 ( .A(n81705), .Z(n105940) );
  CLKBUF_X1 U91877 ( .A(n81705), .Z(n105941) );
  CLKBUF_X1 U91878 ( .A(n95173), .Z(n105528) );
  CLKBUF_X1 U91879 ( .A(n95173), .Z(n105527) );
  CLKBUF_X1 U91880 ( .A(n81312), .Z(n106196) );
  CLKBUF_X1 U91881 ( .A(n81312), .Z(n106195) );
  CLKBUF_X1 U91882 ( .A(n96093), .Z(n105441) );
  CLKBUF_X1 U91883 ( .A(n80185), .Z(n106341) );
  CLKBUF_X1 U91884 ( .A(n81273), .Z(n106252) );
  CLKBUF_X1 U91885 ( .A(n107022), .Z(n105205) );
  CLKBUF_X1 U91886 ( .A(n81260), .Z(n106273) );
  CLKBUF_X1 U91887 ( .A(n81323), .Z(n106183) );
  CLKBUF_X1 U91888 ( .A(n81336), .Z(n106179) );
  CLKBUF_X1 U91889 ( .A(n81785), .Z(n105906) );
  CLKBUF_X1 U91890 ( .A(n81785), .Z(n105905) );
  CLKBUF_X1 U91891 ( .A(n95174), .Z(n105525) );
  CLKBUF_X1 U91892 ( .A(n95174), .Z(n105524) );
  CLKBUF_X1 U91893 ( .A(n81669), .Z(n105955) );
  CLKBUF_X1 U91894 ( .A(n81669), .Z(n105956) );
  CLKBUF_X1 U91895 ( .A(n81706), .Z(n105937) );
  CLKBUF_X1 U91896 ( .A(n81706), .Z(n105938) );
  CLKBUF_X1 U91897 ( .A(n95335), .Z(n105506) );
  CLKBUF_X1 U91898 ( .A(n95335), .Z(n105505) );
  CLKBUF_X1 U91899 ( .A(n95210), .Z(n105516) );
  CLKBUF_X1 U91900 ( .A(n95210), .Z(n105515) );
  CLKBUF_X1 U91901 ( .A(n81789), .Z(n105904) );
  CLKBUF_X1 U91902 ( .A(n106345), .Z(n106347) );
  CLKBUF_X1 U91903 ( .A(n107113), .Z(n105208) );
  CLKBUF_X1 U91904 ( .A(n107113), .Z(n105207) );
  CLKBUF_X1 U91905 ( .A(n81367), .Z(n106144) );
  CLKBUF_X2 U91906 ( .A(n96232), .Z(n105429) );
  CLKBUF_X2 U91907 ( .A(n95913), .Z(n105460) );
  CLKBUF_X1 U91908 ( .A(n94473), .Z(n105632) );
  CLKBUF_X1 U91909 ( .A(n94334), .Z(n105638) );
  CLKBUF_X1 U91910 ( .A(n98659), .Z(n105239) );
  CLKBUF_X1 U91911 ( .A(n98659), .Z(n105238) );
  CLKBUF_X1 U91912 ( .A(n81382), .Z(n106133) );
  CLKBUF_X1 U91913 ( .A(n98695), .Z(n105237) );
  CLKBUF_X1 U91914 ( .A(n98732), .Z(n105236) );
  CLKBUF_X1 U91915 ( .A(n98656), .Z(n105240) );
  CLKBUF_X1 U91916 ( .A(n98616), .Z(n105245) );
  CLKBUF_X1 U91917 ( .A(n94297), .Z(n105640) );
  CLKBUF_X1 U91918 ( .A(n94260), .Z(n105643) );
  CLKBUF_X1 U91919 ( .A(n94400), .Z(n105637) );
  CLKBUF_X1 U91920 ( .A(n94400), .Z(n105636) );
  CLKBUF_X1 U91921 ( .A(n94260), .Z(n105642) );
  CLKBUF_X1 U91922 ( .A(n81774), .Z(n105918) );
  CLKBUF_X1 U91923 ( .A(n96131), .Z(n105437) );
  CLKBUF_X1 U91924 ( .A(n95652), .Z(n105488) );
  CLKBUF_X1 U91925 ( .A(n97261), .Z(n105366) );
  CLKBUF_X1 U91926 ( .A(n81564), .Z(n106025) );
  CLKBUF_X1 U91927 ( .A(n96742), .Z(n105400) );
  CLKBUF_X1 U91928 ( .A(n98301), .Z(n105270) );
  CLKBUF_X1 U91929 ( .A(n97781), .Z(n105312) );
  CLKBUF_X1 U91930 ( .A(n98301), .Z(n105269) );
  CLKBUF_X1 U91931 ( .A(n96053), .Z(n105444) );
  CLKBUF_X1 U91932 ( .A(n81647), .Z(n105976) );
  CLKBUF_X1 U91933 ( .A(n81628), .Z(n105994) );
  CLKBUF_X1 U91934 ( .A(n81745), .Z(n105929) );
  CLKBUF_X1 U91935 ( .A(n81634), .Z(n105983) );
  CLKBUF_X1 U91936 ( .A(n95838), .Z(n105470) );
  CLKBUF_X1 U91937 ( .A(n97101), .Z(n105369) );
  CLKBUF_X1 U91938 ( .A(n81513), .Z(n106041) );
  CLKBUF_X1 U91939 ( .A(n81459), .Z(n106067) );
  CLKBUF_X1 U91940 ( .A(n97357), .Z(n105358) );
  CLKBUF_X1 U91941 ( .A(n81608), .Z(n106002) );
  CLKBUF_X1 U91942 ( .A(n96839), .Z(n105391) );
  CLKBUF_X1 U91943 ( .A(n81540), .Z(n106032) );
  CLKBUF_X1 U91944 ( .A(n81388), .Z(n106122) );
  CLKBUF_X1 U91945 ( .A(n81419), .Z(n106091) );
  CLKBUF_X1 U91946 ( .A(n98540), .Z(n105253) );
  CLKBUF_X1 U91947 ( .A(n97932), .Z(n105294) );
  CLKBUF_X1 U91948 ( .A(n81757), .Z(n105921) );
  CLKBUF_X1 U91949 ( .A(n81619), .Z(n106001) );
  CLKBUF_X1 U91950 ( .A(n81658), .Z(n105967) );
  CLKBUF_X1 U91951 ( .A(n81580), .Z(n106015) );
  CLKBUF_X1 U91952 ( .A(n98130), .Z(n105274) );
  CLKBUF_X1 U91953 ( .A(n96168), .Z(n105433) );
  CLKBUF_X1 U91954 ( .A(n95587), .Z(n105491) );
  CLKBUF_X1 U91955 ( .A(n95453), .Z(n105499) );
  CLKBUF_X1 U91956 ( .A(n97063), .Z(n105370) );
  CLKBUF_X1 U91957 ( .A(n98234), .Z(n105271) );
  CLKBUF_X1 U91958 ( .A(n98166), .Z(n105272) );
  CLKBUF_X1 U91959 ( .A(n97638), .Z(n105333) );
  CLKBUF_X1 U91960 ( .A(n96355), .Z(n105420) );
  CLKBUF_X1 U91961 ( .A(n96295), .Z(n105425) );
  CLKBUF_X1 U91962 ( .A(n95800), .Z(n105474) );
  CLKBUF_X1 U91963 ( .A(n95727), .Z(n105480) );
  CLKBUF_X1 U91964 ( .A(n96681), .Z(n105407) );
  CLKBUF_X1 U91965 ( .A(n96562), .Z(n105409) );
  CLKBUF_X1 U91966 ( .A(n97393), .Z(n105354) );
  CLKBUF_X1 U91967 ( .A(n97320), .Z(n105364) );
  CLKBUF_X1 U91968 ( .A(n98092), .Z(n105276) );
  CLKBUF_X1 U91969 ( .A(n97576), .Z(n105338) );
  CLKBUF_X1 U91970 ( .A(n98092), .Z(n105275) );
  CLKBUF_X1 U91971 ( .A(n81256), .Z(n106274) );
  CLKBUF_X1 U91972 ( .A(n94435), .Z(n105635) );
  CLKBUF_X1 U91973 ( .A(n94435), .Z(n105634) );
  CLKBUF_X1 U91974 ( .A(n96875), .Z(n105385) );
  CLKBUF_X1 U91975 ( .A(n96802), .Z(n105397) );
  CLKBUF_X1 U91976 ( .A(n97712), .Z(n105318) );
  CLKBUF_X1 U91977 ( .A(n98436), .Z(n105261) );
  CLKBUF_X1 U91978 ( .A(n98370), .Z(n105265) );
  CLKBUF_X1 U91979 ( .A(n97842), .Z(n105306) );
  CLKBUF_X1 U91980 ( .A(n97896), .Z(n105300) );
  CLKBUF_X1 U91981 ( .A(n81273), .Z(n106253) );
  CLKBUF_X1 U91982 ( .A(n94473), .Z(n105633) );
  CLKBUF_X1 U91983 ( .A(n94334), .Z(n105639) );
  CLKBUF_X1 U91984 ( .A(n98616), .Z(n105246) );
  CLKBUF_X1 U91985 ( .A(n96742), .Z(n105401) );
  CLKBUF_X1 U91986 ( .A(n97675), .Z(n105326) );
  CLKBUF_X1 U91987 ( .A(n97781), .Z(n105313) );
  CLKBUF_X1 U91988 ( .A(n95764), .Z(n105479) );
  CLKBUF_X1 U91989 ( .A(n95838), .Z(n105471) );
  CLKBUF_X1 U91990 ( .A(n81513), .Z(n106042) );
  CLKBUF_X1 U91991 ( .A(n97357), .Z(n105359) );
  CLKBUF_X1 U91992 ( .A(n81459), .Z(n106068) );
  CLKBUF_X1 U91993 ( .A(n81323), .Z(n106184) );
  CLKBUF_X1 U91994 ( .A(n98540), .Z(n105254) );
  CLKBUF_X1 U91995 ( .A(n81388), .Z(n106123) );
  CLKBUF_X1 U91996 ( .A(n81419), .Z(n106092) );
  CLKBUF_X1 U91997 ( .A(n97932), .Z(n105295) );
  CLKBUF_X1 U91998 ( .A(n81580), .Z(n106016) );
  CLKBUF_X1 U91999 ( .A(n81382), .Z(n106134) );
  CLKBUF_X1 U92000 ( .A(n95413), .Z(n105503) );
  CLKBUF_X1 U92001 ( .A(n81757), .Z(n105922) );
  CLKBUF_X1 U92002 ( .A(n81439), .Z(n106086) );
  CLKBUF_X1 U92003 ( .A(n81336), .Z(n106180) );
  CLKBUF_X1 U92004 ( .A(n81367), .Z(n106145) );
  CLKBUF_X1 U92005 ( .A(n95587), .Z(n105492) );
  CLKBUF_X1 U92006 ( .A(n97576), .Z(n105339) );
  CLKBUF_X1 U92007 ( .A(n97712), .Z(n105319) );
  CLKBUF_X1 U92008 ( .A(n96355), .Z(n105421) );
  CLKBUF_X1 U92009 ( .A(n95800), .Z(n105475) );
  CLKBUF_X1 U92010 ( .A(n97393), .Z(n105355) );
  CLKBUF_X1 U92011 ( .A(n97320), .Z(n105365) );
  CLKBUF_X1 U92012 ( .A(n98436), .Z(n105262) );
  CLKBUF_X1 U92013 ( .A(n98370), .Z(n105266) );
  CLKBUF_X1 U92014 ( .A(n97842), .Z(n105307) );
  CLKBUF_X1 U92015 ( .A(n97896), .Z(n105301) );
  CLKBUF_X1 U92016 ( .A(n94737), .Z(n105597) );
  CLKBUF_X1 U92017 ( .A(n81556), .Z(n106027) );
  CLKBUF_X1 U92018 ( .A(n94508), .Z(n105628) );
  CLKBUF_X1 U92019 ( .A(n94558), .Z(n105617) );
  CLKBUF_X1 U92020 ( .A(n94628), .Z(n105608) );
  CLKBUF_X1 U92021 ( .A(n94775), .Z(n105589) );
  CLKBUF_X1 U92022 ( .A(n95209), .Z(n105520) );
  CLKBUF_X1 U92023 ( .A(n94813), .Z(n105584) );
  CLKBUF_X1 U92024 ( .A(n95334), .Z(n105510) );
  CLKBUF_X1 U92025 ( .A(n81705), .Z(n105942) );
  CLKBUF_X1 U92026 ( .A(n95173), .Z(n105529) );
  CLKBUF_X1 U92027 ( .A(n81668), .Z(n105960) );
  CLKBUF_X1 U92028 ( .A(n81784), .Z(n105910) );
  CLKBUF_X1 U92029 ( .A(n81785), .Z(n105907) );
  CLKBUF_X1 U92030 ( .A(n95174), .Z(n105526) );
  CLKBUF_X1 U92031 ( .A(n81669), .Z(n105957) );
  CLKBUF_X1 U92032 ( .A(n81706), .Z(n105939) );
  CLKBUF_X1 U92033 ( .A(n95335), .Z(n105507) );
  CLKBUF_X1 U92034 ( .A(n95210), .Z(n105517) );
  CLKBUF_X1 U92035 ( .A(n94297), .Z(n105641) );
  CLKBUF_X1 U92036 ( .A(n95451), .Z(n105089) );
  INV_X1 U92037 ( .A(n94330), .ZN(n107116) );
  INV_X1 U92038 ( .A(n94433), .ZN(n107115) );
  INV_X1 U92039 ( .A(n94293), .ZN(n107117) );
  INV_X1 U92040 ( .A(n81798), .ZN(n106759) );
  INV_X1 U92041 ( .A(n98828), .ZN(n106760) );
  INV_X1 U92042 ( .A(n82609), .ZN(n106550) );
  INV_X1 U92043 ( .A(n81211), .ZN(n107024) );
  CLKBUF_X1 U92044 ( .A(n106361), .Z(n106363) );
  CLKBUF_X1 U92045 ( .A(n106361), .Z(n106366) );
  CLKBUF_X1 U92046 ( .A(n106361), .Z(n106364) );
  CLKBUF_X1 U92047 ( .A(n106361), .Z(n106365) );
  CLKBUF_X1 U92048 ( .A(n84106), .Z(n105853) );
  CLKBUF_X1 U92049 ( .A(n85272), .Z(n105791) );
  CLKBUF_X1 U92050 ( .A(n80257), .Z(n106291) );
  CLKBUF_X1 U92051 ( .A(n80214), .Z(n106319) );
  CLKBUF_X1 U92052 ( .A(n84156), .Z(n105829) );
  CLKBUF_X1 U92053 ( .A(n83154), .Z(n105866) );
  CLKBUF_X1 U92054 ( .A(n84152), .Z(n105832) );
  CLKBUF_X1 U92055 ( .A(n80216), .Z(n106317) );
  CLKBUF_X1 U92056 ( .A(n80236), .Z(n106306) );
  CLKBUF_X1 U92057 ( .A(n80210), .Z(n106321) );
  CLKBUF_X1 U92058 ( .A(n85256), .Z(n105804) );
  CLKBUF_X1 U92059 ( .A(n86485), .Z(n105693) );
  CLKBUF_X1 U92060 ( .A(n86495), .Z(n105687) );
  CLKBUF_X1 U92061 ( .A(n85266), .Z(n105797) );
  CLKBUF_X1 U92062 ( .A(n86353), .Z(n105765) );
  CLKBUF_X1 U92063 ( .A(n83137), .Z(n105874) );
  CLKBUF_X1 U92064 ( .A(n84134), .Z(n105842) );
  CLKBUF_X1 U92065 ( .A(n80252), .Z(n106296) );
  CLKBUF_X1 U92066 ( .A(n83131), .Z(n105878) );
  CLKBUF_X1 U92067 ( .A(n86543), .Z(n105669) );
  CLKBUF_X1 U92068 ( .A(n86347), .Z(n105769) );
  CLKBUF_X1 U92069 ( .A(n86335), .Z(n105777) );
  CLKBUF_X1 U92070 ( .A(n86369), .Z(n105757) );
  CLKBUF_X1 U92071 ( .A(n86361), .Z(n105763) );
  CLKBUF_X1 U92072 ( .A(n84140), .Z(n105838) );
  CLKBUF_X1 U92073 ( .A(n80254), .Z(n106294) );
  CLKBUF_X1 U92074 ( .A(n85244), .Z(n105810) );
  CLKBUF_X1 U92075 ( .A(n84148), .Z(n105835) );
  CLKBUF_X1 U92076 ( .A(n80246), .Z(n106300) );
  CLKBUF_X1 U92077 ( .A(n85226), .Z(n105822) );
  CLKBUF_X1 U92078 ( .A(n84130), .Z(n105845) );
  CLKBUF_X1 U92079 ( .A(n85236), .Z(n105816) );
  CLKBUF_X1 U92080 ( .A(n80228), .Z(n106309) );
  CLKBUF_X1 U92081 ( .A(n80220), .Z(n106315) );
  CLKBUF_X1 U92082 ( .A(n80240), .Z(n106304) );
  CLKBUF_X1 U92083 ( .A(n85230), .Z(n105820) );
  CLKBUF_X1 U92084 ( .A(n83160), .Z(n105861) );
  CLKBUF_X1 U92085 ( .A(n80242), .Z(n106302) );
  CLKBUF_X1 U92086 ( .A(n85232), .Z(n105818) );
  CLKBUF_X1 U92087 ( .A(n85268), .Z(n105795) );
  CLKBUF_X1 U92088 ( .A(n83151), .Z(n105868) );
  CLKBUF_X1 U92089 ( .A(n83126), .Z(n105882) );
  CLKBUF_X1 U92090 ( .A(n84110), .Z(n105851) );
  CLKBUF_X1 U92091 ( .A(n85270), .Z(n105793) );
  CLKBUF_X1 U92092 ( .A(n84154), .Z(n105830) );
  CLKBUF_X1 U92093 ( .A(n80208), .Z(n106322) );
  CLKBUF_X1 U92094 ( .A(n83129), .Z(n105879) );
  CLKBUF_X1 U92095 ( .A(n83159), .Z(n105862) );
  CLKBUF_X1 U92096 ( .A(n106737), .Z(n105166) );
  CLKBUF_X1 U92097 ( .A(n80229), .Z(n106308) );
  CLKBUF_X1 U92098 ( .A(n80215), .Z(n106318) );
  CLKBUF_X1 U92099 ( .A(n83136), .Z(n105875) );
  CLKBUF_X1 U92100 ( .A(n85237), .Z(n105815) );
  CLKBUF_X1 U92101 ( .A(n84131), .Z(n105844) );
  CLKBUF_X1 U92102 ( .A(n80247), .Z(n106299) );
  CLKBUF_X1 U92103 ( .A(n83150), .Z(n105869) );
  CLKBUF_X1 U92104 ( .A(n80237), .Z(n106305) );
  CLKBUF_X1 U92105 ( .A(n85233), .Z(n105817) );
  CLKBUF_X1 U92106 ( .A(n83166), .Z(n105854) );
  CLKBUF_X1 U92107 ( .A(n85231), .Z(n105819) );
  CLKBUF_X1 U92108 ( .A(n83123), .Z(n105883) );
  CLKBUF_X1 U92109 ( .A(n83161), .Z(n105860) );
  CLKBUF_X1 U92110 ( .A(n80221), .Z(n106314) );
  CLKBUF_X1 U92111 ( .A(n105173), .Z(n105174) );
  CLKBUF_X1 U92112 ( .A(n105173), .Z(n105175) );
  CLKBUF_X1 U92113 ( .A(n105805), .Z(n105806) );
  CLKBUF_X1 U92114 ( .A(n83132), .Z(n105877) );
  CLKBUF_X1 U92115 ( .A(n80211), .Z(n106320) );
  CLKBUF_X1 U92116 ( .A(n84149), .Z(n105834) );
  CLKBUF_X1 U92117 ( .A(n83138), .Z(n105873) );
  CLKBUF_X1 U92118 ( .A(n84107), .Z(n105852) );
  CLKBUF_X1 U92119 ( .A(n85273), .Z(n105790) );
  CLKBUF_X1 U92120 ( .A(n84135), .Z(n105841) );
  CLKBUF_X1 U92121 ( .A(n80258), .Z(n106290) );
  CLKBUF_X1 U92122 ( .A(n86510), .Z(n105680) );
  CLKBUF_X1 U92123 ( .A(n86410), .Z(n105734) );
  CLKBUF_X1 U92124 ( .A(n86438), .Z(n105718) );
  CLKBUF_X1 U92125 ( .A(n86434), .Z(n105720) );
  CLKBUF_X1 U92126 ( .A(n86352), .Z(n105766) );
  CLKBUF_X1 U92127 ( .A(n80223), .Z(n106312) );
  CLKBUF_X1 U92128 ( .A(n86376), .Z(n105752) );
  CLKBUF_X1 U92129 ( .A(n86544), .Z(n105668) );
  CLKBUF_X1 U92130 ( .A(n84141), .Z(n105837) );
  CLKBUF_X1 U92131 ( .A(n85243), .Z(n105811) );
  CLKBUF_X1 U92132 ( .A(n85267), .Z(n105796) );
  CLKBUF_X1 U92133 ( .A(n85269), .Z(n105794) );
  CLKBUF_X1 U92134 ( .A(n85227), .Z(n105821) );
  CLKBUF_X1 U92135 ( .A(n84153), .Z(n105831) );
  CLKBUF_X1 U92136 ( .A(n85263), .Z(n105798) );
  CLKBUF_X1 U92137 ( .A(n85239), .Z(n105813) );
  CLKBUF_X1 U92138 ( .A(n80249), .Z(n106297) );
  CLKBUF_X1 U92139 ( .A(n83152), .Z(n105867) );
  CLKBUF_X1 U92140 ( .A(n84124), .Z(n105849) );
  CLKBUF_X1 U92141 ( .A(n85224), .Z(n105823) );
  CLKBUF_X1 U92142 ( .A(n106946), .Z(n105197) );
  CLKBUF_X1 U92143 ( .A(n84128), .Z(n105846) );
  CLKBUF_X1 U92144 ( .A(n85250), .Z(n105808) );
  CLKBUF_X1 U92145 ( .A(n85260), .Z(n105800) );
  CLKBUF_X1 U92146 ( .A(\DLX_Datapath/ArithLogUnit/N112 ), .Z(n106368) );
  INV_X1 U92147 ( .A(n81209), .ZN(n106279) );
  CLKBUF_X1 U92148 ( .A(n86555), .Z(n105661) );
  CLKBUF_X1 U92149 ( .A(n86411), .Z(n105733) );
  CLKBUF_X1 U92150 ( .A(n86467), .Z(n105703) );
  CLKBUF_X1 U92151 ( .A(n85238), .Z(n105814) );
  CLKBUF_X1 U92152 ( .A(n80222), .Z(n106313) );
  CLKBUF_X1 U92153 ( .A(n80248), .Z(n106298) );
  CLKBUF_X1 U92154 ( .A(n85258), .Z(n105802) );
  CLKBUF_X1 U92155 ( .A(n85262), .Z(n105799) );
  CLKBUF_X1 U92156 ( .A(n98955), .Z(n105229) );
  CLKBUF_X1 U92157 ( .A(n83122), .Z(n105884) );
  CLKBUF_X1 U92158 ( .A(n83155), .Z(n105865) );
  CLKBUF_X1 U92159 ( .A(n83127), .Z(n105881) );
  CLKBUF_X1 U92160 ( .A(n86484), .Z(n105694) );
  CLKBUF_X1 U92161 ( .A(n86426), .Z(n105726) );
  CLKBUF_X1 U92162 ( .A(n80241), .Z(n106303) );
  CLKBUF_X1 U92163 ( .A(n84158), .Z(n105827) );
  CLKBUF_X1 U92164 ( .A(n81804), .Z(n105096) );
  CLKBUF_X1 U92165 ( .A(n81804), .Z(n105097) );
  INV_X1 U92166 ( .A(n83244), .ZN(n106738) );
  INV_X1 U92167 ( .A(n83239), .ZN(n106739) );
  CLKBUF_X1 U92168 ( .A(n83162), .Z(n105859) );
  INV_X1 U92169 ( .A(n81805), .ZN(n106945) );
  INV_X1 U92170 ( .A(n106132), .ZN(n106131) );
  INV_X1 U92171 ( .A(n106132), .ZN(n106129) );
  INV_X1 U92172 ( .A(n106132), .ZN(n106130) );
  INV_X1 U92173 ( .A(n106132), .ZN(n106128) );
  INV_X1 U92174 ( .A(n106334), .ZN(n106330) );
  INV_X1 U92175 ( .A(n106334), .ZN(n106331) );
  INV_X1 U92176 ( .A(n106334), .ZN(n106332) );
  INV_X1 U92177 ( .A(n106334), .ZN(n106333) );
  INV_X1 U92178 ( .A(n106189), .ZN(n106188) );
  INV_X1 U92179 ( .A(n106189), .ZN(n106187) );
  INV_X1 U92180 ( .A(n106189), .ZN(n106186) );
  INV_X1 U92181 ( .A(n106189), .ZN(n106185) );
  INV_X1 U92182 ( .A(n106194), .ZN(n106193) );
  INV_X1 U92183 ( .A(n106194), .ZN(n106192) );
  INV_X1 U92184 ( .A(n106194), .ZN(n106191) );
  INV_X1 U92185 ( .A(n106194), .ZN(n106190) );
  INV_X1 U92186 ( .A(n106107), .ZN(n106106) );
  INV_X1 U92187 ( .A(n106107), .ZN(n106105) );
  INV_X1 U92188 ( .A(n106107), .ZN(n106104) );
  INV_X1 U92189 ( .A(n106107), .ZN(n106103) );
  INV_X1 U92190 ( .A(n106166), .ZN(n106165) );
  INV_X1 U92191 ( .A(n106166), .ZN(n106164) );
  INV_X1 U92192 ( .A(n106166), .ZN(n106162) );
  INV_X1 U92193 ( .A(n106166), .ZN(n106163) );
  INV_X1 U92194 ( .A(n106222), .ZN(n106221) );
  INV_X1 U92195 ( .A(n106222), .ZN(n106220) );
  INV_X1 U92196 ( .A(n106222), .ZN(n106219) );
  INV_X1 U92197 ( .A(n106222), .ZN(n106218) );
  INV_X1 U92198 ( .A(n106112), .ZN(n106111) );
  INV_X1 U92199 ( .A(n106112), .ZN(n106110) );
  INV_X1 U92200 ( .A(n106112), .ZN(n106109) );
  INV_X1 U92201 ( .A(n106112), .ZN(n106108) );
  INV_X1 U92202 ( .A(n106161), .ZN(n106160) );
  INV_X1 U92203 ( .A(n106161), .ZN(n106159) );
  INV_X1 U92204 ( .A(n106161), .ZN(n106158) );
  INV_X1 U92205 ( .A(n106161), .ZN(n106157) );
  INV_X1 U92206 ( .A(n106201), .ZN(n106200) );
  INV_X1 U92207 ( .A(n106201), .ZN(n106199) );
  INV_X1 U92208 ( .A(n106201), .ZN(n106197) );
  INV_X1 U92209 ( .A(n106201), .ZN(n106198) );
  INV_X1 U92210 ( .A(n106117), .ZN(n106116) );
  INV_X1 U92211 ( .A(n106117), .ZN(n106115) );
  INV_X1 U92212 ( .A(n106117), .ZN(n106114) );
  INV_X1 U92213 ( .A(n106117), .ZN(n106113) );
  INV_X1 U92214 ( .A(n106263), .ZN(n106262) );
  INV_X1 U92215 ( .A(n106263), .ZN(n106261) );
  INV_X1 U92216 ( .A(n106263), .ZN(n106260) );
  INV_X1 U92217 ( .A(n106263), .ZN(n106259) );
  INV_X1 U92218 ( .A(n106047), .ZN(n106046) );
  INV_X1 U92219 ( .A(n106047), .ZN(n106045) );
  INV_X1 U92220 ( .A(n106047), .ZN(n106044) );
  INV_X1 U92221 ( .A(n106047), .ZN(n106043) );
  INV_X1 U92222 ( .A(n106052), .ZN(n106051) );
  INV_X1 U92223 ( .A(n106052), .ZN(n106050) );
  INV_X1 U92224 ( .A(n106052), .ZN(n106049) );
  INV_X1 U92225 ( .A(n106052), .ZN(n106048) );
  INV_X1 U92226 ( .A(n106057), .ZN(n106056) );
  INV_X1 U92227 ( .A(n106057), .ZN(n106055) );
  INV_X1 U92228 ( .A(n106057), .ZN(n106054) );
  INV_X1 U92229 ( .A(n106057), .ZN(n106053) );
  INV_X1 U92230 ( .A(n106097), .ZN(n106096) );
  INV_X1 U92231 ( .A(n106097), .ZN(n106095) );
  INV_X1 U92232 ( .A(n106097), .ZN(n106093) );
  INV_X1 U92233 ( .A(n106097), .ZN(n106094) );
  INV_X1 U92234 ( .A(n106247), .ZN(n106246) );
  INV_X1 U92235 ( .A(n106247), .ZN(n106245) );
  INV_X1 U92236 ( .A(n106247), .ZN(n106243) );
  INV_X1 U92237 ( .A(n106247), .ZN(n106244) );
  INV_X1 U92238 ( .A(n106239), .ZN(n106238) );
  INV_X1 U92239 ( .A(n106239), .ZN(n106237) );
  INV_X1 U92240 ( .A(n106239), .ZN(n106235) );
  INV_X1 U92241 ( .A(n106239), .ZN(n106236) );
  INV_X1 U92242 ( .A(n106174), .ZN(n106173) );
  INV_X1 U92243 ( .A(n106174), .ZN(n106172) );
  INV_X1 U92244 ( .A(n106174), .ZN(n106170) );
  INV_X1 U92245 ( .A(n106174), .ZN(n106171) );
  INV_X1 U92246 ( .A(n106234), .ZN(n106233) );
  INV_X1 U92247 ( .A(n106234), .ZN(n106232) );
  INV_X1 U92248 ( .A(n106234), .ZN(n106231) );
  INV_X1 U92249 ( .A(n106234), .ZN(n106230) );
  INV_X1 U92250 ( .A(n106073), .ZN(n106072) );
  INV_X1 U92251 ( .A(n106073), .ZN(n106071) );
  INV_X1 U92252 ( .A(n106073), .ZN(n106070) );
  INV_X1 U92253 ( .A(n106073), .ZN(n106069) );
  INV_X1 U92254 ( .A(n106270), .ZN(n106269) );
  INV_X1 U92255 ( .A(n106270), .ZN(n106268) );
  INV_X1 U92256 ( .A(n106270), .ZN(n106267) );
  INV_X1 U92257 ( .A(n106270), .ZN(n106266) );
  INV_X1 U92258 ( .A(n105513), .ZN(n105512) );
  INV_X1 U92259 ( .A(n105513), .ZN(n105511) );
  INV_X1 U92260 ( .A(n105963), .ZN(n105961) );
  INV_X1 U92261 ( .A(n105945), .ZN(n105943) );
  INV_X1 U92262 ( .A(n105945), .ZN(n105944) );
  INV_X1 U92263 ( .A(n105963), .ZN(n105962) );
  INV_X1 U92264 ( .A(n105532), .ZN(n105531) );
  INV_X1 U92265 ( .A(n105532), .ZN(n105530) );
  INV_X1 U92266 ( .A(n105914), .ZN(n105913) );
  INV_X1 U92267 ( .A(n105914), .ZN(n105912) );
  INV_X1 U92268 ( .A(n105523), .ZN(n105522) );
  INV_X1 U92269 ( .A(n105523), .ZN(n105521) );
  INV_X1 U92270 ( .A(n81795), .ZN(n105903) );
  CLKBUF_X1 U92271 ( .A(n98804), .Z(n105233) );
  CLKBUF_X1 U92272 ( .A(n98804), .Z(n105234) );
  CLKBUF_X1 U92273 ( .A(n106751), .Z(n105180) );
  CLKBUF_X1 U92274 ( .A(n106749), .Z(n105176) );
  INV_X1 U92275 ( .A(n95038), .ZN(n105554) );
  INV_X1 U92276 ( .A(n94935), .ZN(n105566) );
  INV_X1 U92277 ( .A(n98802), .ZN(n105235) );
  INV_X1 U92278 ( .A(n106007), .ZN(n106012) );
  INV_X1 U92279 ( .A(n94556), .ZN(n105620) );
  INV_X1 U92280 ( .A(n81680), .ZN(n105954) );
  CLKBUF_X2 U92281 ( .A(n97575), .Z(n105126) );
  CLKBUF_X2 U92282 ( .A(n82027), .Z(n105893) );
  CLKBUF_X1 U92283 ( .A(n106752), .Z(n105183) );
  INV_X1 U92284 ( .A(n95131), .ZN(n111023) );
  INV_X1 U92285 ( .A(n80097), .ZN(n106597) );
  CLKBUF_X1 U92286 ( .A(n95451), .Z(n105090) );
  CLKBUF_X1 U92287 ( .A(n95451), .Z(n105091) );
  CLKBUF_X1 U92288 ( .A(n95451), .Z(n105094) );
  CLKBUF_X1 U92289 ( .A(n105094), .Z(n105092) );
  CLKBUF_X1 U92290 ( .A(n105095), .Z(n105093) );
  CLKBUF_X1 U92291 ( .A(n105090), .Z(n105095) );
  INV_X1 U92292 ( .A(n94999), .ZN(n111025) );
  INV_X1 U92293 ( .A(n94397), .ZN(n106758) );
  INV_X1 U92294 ( .A(n96125), .ZN(n107127) );
  INV_X1 U92295 ( .A(n94468), .ZN(n107113) );
  INV_X1 U92296 ( .A(n81230), .ZN(n107026) );
  INV_X1 U92297 ( .A(n105858), .ZN(n105857) );
  INV_X1 U92298 ( .A(n105227), .ZN(n105226) );
  CLKBUF_X1 U92299 ( .A(n83145), .Z(n105871) );
  CLKBUF_X1 U92300 ( .A(n86509), .Z(n105681) );
  CLKBUF_X1 U92301 ( .A(n86553), .Z(n105663) );
  CLKBUF_X1 U92302 ( .A(n86541), .Z(n105671) );
  CLKBUF_X1 U92303 ( .A(n86469), .Z(n105701) );
  CLKBUF_X1 U92304 ( .A(n86449), .Z(n105715) );
  CLKBUF_X1 U92305 ( .A(n86451), .Z(n105713) );
  CLKBUF_X1 U92306 ( .A(n86497), .Z(n105685) );
  CLKBUF_X1 U92307 ( .A(n86489), .Z(n105691) );
  CLKBUF_X1 U92308 ( .A(n86491), .Z(n105689) );
  CLKBUF_X1 U92309 ( .A(n86483), .Z(n105695) );
  CLKBUF_X1 U92310 ( .A(n86477), .Z(n105699) );
  CLKBUF_X1 U92311 ( .A(n86409), .Z(n105735) );
  CLKBUF_X1 U92312 ( .A(n86399), .Z(n105741) );
  CLKBUF_X1 U92313 ( .A(n86391), .Z(n105747) );
  CLKBUF_X1 U92314 ( .A(n86393), .Z(n105745) );
  CLKBUF_X1 U92315 ( .A(n86437), .Z(n105719) );
  CLKBUF_X1 U92316 ( .A(n86439), .Z(n105717) );
  CLKBUF_X1 U92317 ( .A(n86431), .Z(n105723) );
  CLKBUF_X1 U92318 ( .A(n86433), .Z(n105721) );
  CLKBUF_X1 U92319 ( .A(n86425), .Z(n105727) );
  CLKBUF_X1 U92320 ( .A(n86419), .Z(n105731) );
  CLKBUF_X1 U92321 ( .A(n86421), .Z(n105729) );
  CLKBUF_X1 U92322 ( .A(n86351), .Z(n105767) );
  CLKBUF_X1 U92323 ( .A(n86345), .Z(n105771) );
  CLKBUF_X1 U92324 ( .A(n86457), .Z(n105709) );
  CLKBUF_X1 U92325 ( .A(n86397), .Z(n105743) );
  CLKBUF_X1 U92326 ( .A(n86479), .Z(n105697) );
  CLKBUF_X1 U92327 ( .A(n86427), .Z(n105725) );
  CLKBUF_X1 U92328 ( .A(n85242), .Z(n105812) );
  CLKBUF_X1 U92329 ( .A(n86463), .Z(n105705) );
  CLKBUF_X1 U92330 ( .A(n86535), .Z(n105675) );
  CLKBUF_X1 U92331 ( .A(n86525), .Z(n105676) );
  CLKBUF_X1 U92332 ( .A(n86513), .Z(n105679) );
  CLKBUF_X1 U92333 ( .A(n86507), .Z(n105683) );
  CLKBUF_X1 U92334 ( .A(n86547), .Z(n105667) );
  CLKBUF_X1 U92335 ( .A(n86537), .Z(n105673) );
  CLKBUF_X1 U92336 ( .A(n86341), .Z(n105773) );
  CLKBUF_X1 U92337 ( .A(n86333), .Z(n105779) );
  CLKBUF_X1 U92338 ( .A(n86379), .Z(n105751) );
  CLKBUF_X1 U92339 ( .A(n86381), .Z(n105749) );
  CLKBUF_X1 U92340 ( .A(n86373), .Z(n105755) );
  CLKBUF_X1 U92341 ( .A(n86375), .Z(n105753) );
  CLKBUF_X1 U92342 ( .A(n86367), .Z(n105759) );
  CLKBUF_X1 U92343 ( .A(n84138), .Z(n105840) );
  CLKBUF_X1 U92344 ( .A(n80226), .Z(n106311) );
  CLKBUF_X1 U92345 ( .A(n83135), .Z(n105876) );
  CLKBUF_X1 U92346 ( .A(n83128), .Z(n105880) );
  CLKBUF_X1 U92347 ( .A(n90519), .Z(n105645) );
  CLKBUF_X1 U92348 ( .A(n98953), .Z(n105231) );
  CLKBUF_X1 U92349 ( .A(n99022), .Z(n105225) );
  CLKBUF_X1 U92350 ( .A(n80260), .Z(n106283) );
  CLKBUF_X1 U92351 ( .A(n106285), .Z(n106284) );
  CLKBUF_X1 U92352 ( .A(n84139), .Z(n105839) );
  CLKBUF_X1 U92353 ( .A(n85245), .Z(n105809) );
  CLKBUF_X1 U92354 ( .A(n106282), .Z(n106285) );
  CLKBUF_X1 U92355 ( .A(n106745), .Z(n105171) );
  CLKBUF_X1 U92356 ( .A(n106745), .Z(n105172) );
  CLKBUF_X1 U92357 ( .A(n86508), .Z(n105682) );
  CLKBUF_X1 U92358 ( .A(n86514), .Z(n105678) );
  CLKBUF_X1 U92359 ( .A(n86556), .Z(n105660) );
  CLKBUF_X1 U92360 ( .A(n86462), .Z(n105706) );
  CLKBUF_X1 U92361 ( .A(n86458), .Z(n105708) );
  CLKBUF_X1 U92362 ( .A(n86452), .Z(n105712) );
  CLKBUF_X1 U92363 ( .A(n86496), .Z(n105686) );
  CLKBUF_X1 U92364 ( .A(n86498), .Z(n105684) );
  CLKBUF_X1 U92365 ( .A(n86492), .Z(n105688) );
  CLKBUF_X1 U92366 ( .A(n86478), .Z(n105698) );
  CLKBUF_X1 U92367 ( .A(n86480), .Z(n105696) );
  CLKBUF_X1 U92368 ( .A(n86404), .Z(n105738) );
  CLKBUF_X1 U92369 ( .A(n86398), .Z(n105742) );
  CLKBUF_X1 U92370 ( .A(n86392), .Z(n105746) );
  CLKBUF_X1 U92371 ( .A(n86394), .Z(n105744) );
  CLKBUF_X1 U92372 ( .A(n86432), .Z(n105722) );
  CLKBUF_X1 U92373 ( .A(n86422), .Z(n105728) );
  CLKBUF_X1 U92374 ( .A(n86342), .Z(n105772) );
  CLKBUF_X1 U92375 ( .A(n86406), .Z(n105736) );
  CLKBUF_X1 U92376 ( .A(n86440), .Z(n105716) );
  CLKBUF_X1 U92377 ( .A(n86464), .Z(n105704) );
  CLKBUF_X1 U92378 ( .A(n86456), .Z(n105710) );
  CLKBUF_X1 U92379 ( .A(n106949), .Z(n105198) );
  CLKBUF_X1 U92380 ( .A(n86554), .Z(n105662) );
  CLKBUF_X1 U92381 ( .A(n86548), .Z(n105666) );
  CLKBUF_X1 U92382 ( .A(n86550), .Z(n105664) );
  CLKBUF_X1 U92383 ( .A(n86536), .Z(n105674) );
  CLKBUF_X1 U92384 ( .A(n86538), .Z(n105672) );
  CLKBUF_X1 U92385 ( .A(n86468), .Z(n105702) );
  CLKBUF_X1 U92386 ( .A(n86348), .Z(n105768) );
  CLKBUF_X1 U92387 ( .A(n86340), .Z(n105774) );
  CLKBUF_X1 U92388 ( .A(n86334), .Z(n105778) );
  CLKBUF_X1 U92389 ( .A(n86336), .Z(n105776) );
  CLKBUF_X1 U92390 ( .A(n86380), .Z(n105750) );
  CLKBUF_X1 U92391 ( .A(n86374), .Z(n105754) );
  CLKBUF_X1 U92392 ( .A(n86370), .Z(n105756) );
  CLKBUF_X1 U92393 ( .A(n86362), .Z(n105762) );
  CLKBUF_X1 U92394 ( .A(n86382), .Z(n105748) );
  CLKBUF_X1 U92395 ( .A(n86364), .Z(n105760) );
  CLKBUF_X1 U92396 ( .A(n99027), .Z(n105223) );
  CLKBUF_X1 U92397 ( .A(n98954), .Z(n105230) );
  CLKBUF_X1 U92398 ( .A(n98956), .Z(n105228) );
  CLKBUF_X1 U92399 ( .A(n80243), .Z(n106301) );
  CLKBUF_X1 U92400 ( .A(n86318), .Z(n105782) );
  CLKBUF_X1 U92401 ( .A(n80234), .Z(n106307) );
  CLKBUF_X1 U92402 ( .A(n106934), .Z(n105195) );
  CLKBUF_X1 U92403 ( .A(n94109), .Z(n105143) );
  CLKBUF_X1 U92404 ( .A(n86403), .Z(n105739) );
  CLKBUF_X1 U92405 ( .A(n86549), .Z(n105665) );
  CLKBUF_X1 U92406 ( .A(n86363), .Z(n105761) );
  CLKBUF_X1 U92407 ( .A(n99026), .Z(n105224) );
  CLKBUF_X1 U92408 ( .A(n94127), .Z(n105142) );
  CLKBUF_X1 U92409 ( .A(n80227), .Z(n106310) );
  CLKBUF_X1 U92410 ( .A(n86516), .Z(n105677) );
  CLKBUF_X1 U92411 ( .A(n86450), .Z(n105714) );
  CLKBUF_X1 U92412 ( .A(n86490), .Z(n105690) );
  CLKBUF_X1 U92413 ( .A(n86428), .Z(n105724) );
  CLKBUF_X1 U92414 ( .A(n86368), .Z(n105758) );
  INV_X1 U92415 ( .A(n81232), .ZN(n106743) );
  INV_X1 U92416 ( .A(n81806), .ZN(n107481) );
  INV_X1 U92417 ( .A(n83114), .ZN(n106737) );
  INV_X1 U92418 ( .A(n94176), .ZN(n107095) );
  CLKBUF_X1 U92419 ( .A(n81804), .Z(n105098) );
  INV_X1 U92420 ( .A(n90189), .ZN(n107059) );
  INV_X1 U92421 ( .A(n99012), .ZN(n107480) );
  INV_X1 U92422 ( .A(\DLX_Datapath/ArithLogUnit/N177 ), .ZN(n106946) );
  INV_X1 U92423 ( .A(n84086), .ZN(n106740) );
  INV_X1 U92424 ( .A(n81977), .ZN(n111138) );
  INV_X1 U92425 ( .A(n99542), .ZN(n107482) );
  INV_X1 U92426 ( .A(n85180), .ZN(n106733) );
  INV_X1 U92427 ( .A(n99215), .ZN(n107519) );
  INV_X1 U92428 ( .A(n99505), .ZN(n107469) );
  CLKBUF_X1 U92429 ( .A(n106362), .Z(n106361) );
  INV_X1 U92430 ( .A(n86189), .ZN(n106699) );
  INV_X1 U92431 ( .A(n86210), .ZN(n106698) );
  INV_X1 U92432 ( .A(n85183), .ZN(n106734) );
  INV_X1 U92433 ( .A(n81210), .ZN(n106742) );
  INV_X1 U92434 ( .A(n99031), .ZN(n107479) );
  CLKBUF_X1 U92435 ( .A(n85253), .Z(n105805) );
  INV_X1 U92436 ( .A(n81242), .ZN(n106744) );
  INV_X1 U92437 ( .A(n85169), .ZN(n106736) );
  INV_X1 U92438 ( .A(n85185), .ZN(n106735) );
  INV_X1 U92439 ( .A(n99625), .ZN(n108744) );
  INV_X1 U92440 ( .A(n99488), .ZN(n109087) );
  INV_X1 U92441 ( .A(n79744), .ZN(n106948) );
  INV_X1 U92442 ( .A(n86222), .ZN(n106958) );
  CLKBUF_X1 U92443 ( .A(n82862), .Z(n105885) );
  INV_X1 U92444 ( .A(n94851), .ZN(n106763) );
  CLKBUF_X1 U92445 ( .A(n98619), .Z(n105242) );
  CLKBUF_X1 U92446 ( .A(n98619), .Z(n105241) );
  CLKBUF_X1 U92447 ( .A(n80189), .Z(n106335) );
  CLKBUF_X1 U92448 ( .A(n80189), .Z(n106336) );
  CLKBUF_X1 U92449 ( .A(n96091), .Z(n105443) );
  CLKBUF_X1 U92450 ( .A(n96091), .Z(n105442) );
  CLKBUF_X1 U92451 ( .A(n79971), .Z(n106352) );
  CLKBUF_X1 U92452 ( .A(n81925), .Z(n105898) );
  INV_X1 U92453 ( .A(n94848), .ZN(n111024) );
  INV_X1 U92454 ( .A(n95332), .ZN(n105513) );
  INV_X1 U92455 ( .A(n81666), .ZN(n105963) );
  INV_X1 U92456 ( .A(n81703), .ZN(n105945) );
  INV_X1 U92457 ( .A(n95171), .ZN(n105532) );
  INV_X1 U92458 ( .A(n81781), .ZN(n105914) );
  INV_X1 U92459 ( .A(n95207), .ZN(n105523) );
  INV_X1 U92460 ( .A(n81895), .ZN(n106696) );
  CLKBUF_X1 U92461 ( .A(n79971), .Z(n106353) );
  CLKBUF_X1 U92462 ( .A(n98618), .Z(n105244) );
  INV_X1 U92463 ( .A(n82885), .ZN(n111051) );
  INV_X1 U92464 ( .A(n95036), .ZN(n106748) );
  CLKBUF_X1 U92465 ( .A(n80189), .Z(n106337) );
  INV_X1 U92466 ( .A(n95412), .ZN(n107126) );
  INV_X1 U92467 ( .A(n82882), .ZN(n107159) );
  CLKBUF_X1 U92468 ( .A(n105502), .Z(n105500) );
  INV_X1 U92469 ( .A(n90119), .ZN(n107122) );
  INV_X1 U92470 ( .A(n82377), .ZN(n106780) );
  INV_X1 U92471 ( .A(n82990), .ZN(n108628) );
  INV_X1 U92472 ( .A(n83050), .ZN(n107163) );
  INV_X1 U92473 ( .A(n83014), .ZN(n107624) );
  INV_X1 U92474 ( .A(n82867), .ZN(n107628) );
  INV_X1 U92475 ( .A(n82614), .ZN(n106551) );
  INV_X1 U92476 ( .A(n82604), .ZN(n106552) );
  CLKBUF_X1 U92477 ( .A(n81588), .Z(n106007) );
  INV_X1 U92478 ( .A(n81903), .ZN(n106517) );
  INV_X1 U92479 ( .A(n82665), .ZN(n106771) );
  INV_X1 U92480 ( .A(n82289), .ZN(n106806) );
  INV_X1 U92481 ( .A(n82277), .ZN(n106844) );
  INV_X1 U92482 ( .A(n82594), .ZN(n106808) );
  INV_X1 U92483 ( .A(n95167), .ZN(n106751) );
  INV_X1 U92484 ( .A(n95034), .ZN(n106752) );
  INV_X1 U92485 ( .A(n95408), .ZN(n106749) );
  INV_X1 U92486 ( .A(n95298), .ZN(n106750) );
  INV_X1 U92487 ( .A(n90120), .ZN(n107114) );
  INV_X1 U92488 ( .A(n94366), .ZN(n107022) );
  INV_X1 U92489 ( .A(n82877), .ZN(n106829) );
  INV_X1 U92490 ( .A(n82962), .ZN(n108624) );
  INV_X1 U92491 ( .A(n82608), .ZN(n106553) );
  CLKBUF_X1 U92492 ( .A(n105502), .Z(n105501) );
  INV_X1 U92493 ( .A(n87266), .ZN(n107384) );
  INV_X1 U92494 ( .A(n87148), .ZN(n107382) );
  INV_X1 U92495 ( .A(n86912), .ZN(n107378) );
  INV_X1 U92496 ( .A(n89271), .ZN(n108974) );
  INV_X1 U92497 ( .A(n87030), .ZN(n107380) );
  INV_X1 U92498 ( .A(n86558), .ZN(n107373) );
  INV_X1 U92499 ( .A(n86303), .ZN(n107371) );
  INV_X1 U92500 ( .A(n86794), .ZN(n107376) );
  INV_X1 U92501 ( .A(n86676), .ZN(n106832) );
  INV_X1 U92502 ( .A(n100262), .ZN(n107148) );
  INV_X1 U92503 ( .A(n100146), .ZN(n108742) );
  INV_X1 U92504 ( .A(n100063), .ZN(n109088) );
  INV_X1 U92505 ( .A(n99186), .ZN(n106927) );
  INV_X1 U92506 ( .A(n99024), .ZN(n106929) );
  INV_X1 U92507 ( .A(n99404), .ZN(n108504) );
  INV_X1 U92508 ( .A(n99517), .ZN(n109085) );
  INV_X1 U92509 ( .A(n99665), .ZN(n108741) );
  INV_X1 U92510 ( .A(n81817), .ZN(n108272) );
  INV_X1 U92511 ( .A(n99383), .ZN(n107739) );
  INV_X1 U92512 ( .A(n99382), .ZN(n107737) );
  INV_X1 U92513 ( .A(n99850), .ZN(n107560) );
  INV_X1 U92514 ( .A(n106328), .ZN(n106326) );
  INV_X1 U92515 ( .A(n106328), .ZN(n106325) );
  INV_X1 U92516 ( .A(n106328), .ZN(n106324) );
  INV_X1 U92517 ( .A(n106328), .ZN(n106323) );
  INV_X1 U92518 ( .A(n82399), .ZN(n111134) );
  CLKBUF_X1 U92519 ( .A(\DLX_Datapath/ArithLogUnit/N178 ), .Z(n106369) );
  CLKBUF_X1 U92520 ( .A(n83165), .Z(n105855) );
  CLKBUF_X1 U92521 ( .A(n86405), .Z(n105737) );
  CLKBUF_X1 U92522 ( .A(n86339), .Z(n105775) );
  CLKBUF_X1 U92523 ( .A(n86461), .Z(n105707) );
  CLKBUF_X1 U92524 ( .A(n86455), .Z(n105711) );
  CLKBUF_X1 U92525 ( .A(n90511), .Z(n105650) );
  CLKBUF_X1 U92526 ( .A(n90513), .Z(n105648) );
  CLKBUF_X1 U92527 ( .A(n90507), .Z(n105651) );
  CLKBUF_X1 U92528 ( .A(n90309), .Z(n105654) );
  CLKBUF_X1 U92529 ( .A(n86319), .Z(n105781) );
  CLKBUF_X1 U92530 ( .A(n80259), .Z(n106287) );
  CLKBUF_X1 U92531 ( .A(n83164), .Z(n105856) );
  CLKBUF_X1 U92532 ( .A(n99625), .Z(n105109) );
  INV_X1 U92533 ( .A(n98972), .ZN(n108747) );
  CLKBUF_X1 U92534 ( .A(n106286), .Z(n106288) );
  CLKBUF_X1 U92535 ( .A(n106286), .Z(n106289) );
  CLKBUF_X1 U92536 ( .A(n85271), .Z(n105792) );
  CLKBUF_X1 U92537 ( .A(n86486), .Z(n105692) );
  CLKBUF_X1 U92538 ( .A(n86412), .Z(n105732) );
  CLKBUF_X1 U92539 ( .A(n86420), .Z(n105730) );
  CLKBUF_X1 U92540 ( .A(n86354), .Z(n105764) );
  CLKBUF_X1 U92541 ( .A(n86542), .Z(n105670) );
  CLKBUF_X1 U92542 ( .A(n86470), .Z(n105700) );
  CLKBUF_X1 U92543 ( .A(n90518), .Z(n105646) );
  CLKBUF_X1 U92544 ( .A(n90514), .Z(n105647) );
  CLKBUF_X1 U92545 ( .A(n90512), .Z(n105649) );
  CLKBUF_X1 U92546 ( .A(n90306), .Z(n105655) );
  CLKBUF_X1 U92547 ( .A(n86306), .Z(n105787) );
  CLKBUF_X1 U92548 ( .A(n86311), .Z(n105785) );
  CLKBUF_X1 U92549 ( .A(n90303), .Z(n105657) );
  CLKBUF_X1 U92550 ( .A(n60159), .Z(n106359) );
  CLKBUF_X1 U92551 ( .A(n99764), .Z(n105103) );
  INV_X1 U92552 ( .A(n82628), .ZN(n111145) );
  INV_X1 U92553 ( .A(n94245), .ZN(n107098) );
  INV_X1 U92554 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[16] ), .ZN(
        n107490) );
  INV_X1 U92555 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[17] ), .ZN(
        n107484) );
  CLKBUF_X1 U92556 ( .A(n99667), .Z(n105106) );
  CLKBUF_X1 U92557 ( .A(n99515), .Z(n105112) );
  CLKBUF_X1 U92558 ( .A(n99402), .Z(n105118) );
  CLKBUF_X1 U92559 ( .A(n81819), .Z(n105122) );
  INV_X1 U92560 ( .A(n79788), .ZN(n107586) );
  CLKBUF_X1 U92561 ( .A(n86234), .Z(n105788) );
  CLKBUF_X1 U92562 ( .A(n99624), .Z(n105107) );
  INV_X1 U92563 ( .A(n98996), .ZN(n105227) );
  INV_X1 U92564 ( .A(n86266), .ZN(n106934) );
  INV_X1 U92565 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[16] ), .ZN(
        n107558) );
  INV_X1 U92566 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/m_A[17] ), .ZN(
        n107556) );
  CLKBUF_X1 U92567 ( .A(n94129), .Z(n105140) );
  CLKBUF_X1 U92568 ( .A(n99718), .Z(n105105) );
  CLKBUF_X1 U92569 ( .A(n99623), .Z(n105108) );
  CLKBUF_X1 U92570 ( .A(n99541), .Z(n105111) );
  CLKBUF_X1 U92571 ( .A(n99429), .Z(n105117) );
  CLKBUF_X1 U92572 ( .A(n99015), .Z(n105121) );
  CLKBUF_X1 U92573 ( .A(n86400), .Z(n105740) );
  CLKBUF_X1 U92574 ( .A(n86346), .Z(n105770) );
  CLKBUF_X1 U92575 ( .A(n90520), .Z(n105644) );
  CLKBUF_X1 U92576 ( .A(n84113), .Z(n105850) );
  CLKBUF_X1 U92577 ( .A(n90298), .Z(n105659) );
  INV_X1 U92578 ( .A(n86215), .ZN(n106697) );
  CLKBUF_X1 U92579 ( .A(n60158), .Z(n106360) );
  CLKBUF_X1 U92580 ( .A(n99488), .Z(n105113) );
  CLKBUF_X1 U92581 ( .A(n106444), .Z(n106371) );
  CLKBUF_X1 U92582 ( .A(n106426), .Z(n106372) );
  INV_X1 U92583 ( .A(n83259), .ZN(n106761) );
  INV_X1 U92584 ( .A(n82387), .ZN(n111136) );
  INV_X1 U92585 ( .A(n90271), .ZN(n107100) );
  INV_X1 U92586 ( .A(n94066), .ZN(n107118) );
  CLKBUF_X1 U92587 ( .A(n105900), .Z(n105899) );
  CLKBUF_X1 U92588 ( .A(n99540), .Z(n105110) );
  CLKBUF_X1 U92589 ( .A(n99428), .Z(n105116) );
  CLKBUF_X1 U92590 ( .A(n99039), .Z(n105119) );
  CLKBUF_X1 U92591 ( .A(n99487), .Z(n105114) );
  INV_X1 U92592 ( .A(n94254), .ZN(n107097) );
  CLKBUF_X1 U92593 ( .A(n81199), .Z(n105100) );
  CLKBUF_X1 U92594 ( .A(n81199), .Z(n105099) );
  CLKBUF_X1 U92595 ( .A(n99719), .Z(n105104) );
  CLKBUF_X1 U92596 ( .A(n81199), .Z(n105101) );
  INV_X1 U92597 ( .A(n99321), .ZN(n106930) );
  INV_X1 U92598 ( .A(n80099), .ZN(n111118) );
  INV_X1 U92599 ( .A(n82617), .ZN(n106949) );
  CLKBUF_X1 U92600 ( .A(n99016), .Z(n105120) );
  INV_X1 U92601 ( .A(n99849), .ZN(n107570) );
  INV_X1 U92602 ( .A(n99058), .ZN(n107476) );
  INV_X1 U92603 ( .A(n90190), .ZN(n107093) );
  INV_X1 U92604 ( .A(n100192), .ZN(n106878) );
  INV_X1 U92605 ( .A(n86202), .ZN(n106700) );
  INV_X1 U92606 ( .A(n80100), .ZN(n111137) );
  INV_X1 U92607 ( .A(n86220), .ZN(n107025) );
  INV_X1 U92608 ( .A(n81909), .ZN(n106747) );
  INV_X1 U92609 ( .A(n99178), .ZN(n107492) );
  INV_X1 U92610 ( .A(n99098), .ZN(n107458) );
  INV_X1 U92611 ( .A(n99100), .ZN(n107454) );
  INV_X1 U92612 ( .A(n99678), .ZN(n107444) );
  INV_X1 U92613 ( .A(n99128), .ZN(n107437) );
  INV_X1 U92614 ( .A(n99138), .ZN(n107434) );
  INV_X1 U92615 ( .A(n99925), .ZN(n107517) );
  INV_X1 U92616 ( .A(n99119), .ZN(n107446) );
  INV_X1 U92617 ( .A(n99109), .ZN(n107453) );
  INV_X1 U92618 ( .A(n99738), .ZN(n107486) );
  INV_X1 U92619 ( .A(n99497), .ZN(n107461) );
  INV_X1 U92620 ( .A(n99078), .ZN(n107465) );
  INV_X1 U92621 ( .A(n99454), .ZN(n107472) );
  INV_X1 U92622 ( .A(n99415), .ZN(n107471) );
  INV_X1 U92623 ( .A(n90108), .ZN(n107136) );
  INV_X1 U92624 ( .A(n99319), .ZN(n106928) );
  INV_X1 U92625 ( .A(n100191), .ZN(n106879) );
  INV_X1 U92626 ( .A(n81976), .ZN(n111127) );
  INV_X1 U92627 ( .A(n79698), .ZN(n107584) );
  INV_X1 U92628 ( .A(n79699), .ZN(n107583) );
  INV_X1 U92629 ( .A(n79695), .ZN(n107580) );
  INV_X1 U92630 ( .A(n79696), .ZN(n107579) );
  INV_X1 U92631 ( .A(n79704), .ZN(n107589) );
  INV_X1 U92632 ( .A(n79705), .ZN(n107588) );
  INV_X1 U92633 ( .A(n79692), .ZN(n107602) );
  INV_X1 U92634 ( .A(n79693), .ZN(n107601) );
  INV_X1 U92635 ( .A(n79689), .ZN(n107607) );
  INV_X1 U92636 ( .A(n79690), .ZN(n107606) );
  INV_X1 U92637 ( .A(n79686), .ZN(n107613) );
  INV_X1 U92638 ( .A(n79687), .ZN(n107612) );
  INV_X1 U92639 ( .A(n79701), .ZN(n107594) );
  INV_X1 U92640 ( .A(n79702), .ZN(n107593) );
  CLKBUF_X1 U92641 ( .A(n80200), .Z(n106329) );
  CLKBUF_X1 U92642 ( .A(n80256), .Z(n106292) );
  CLKBUF_X1 U92643 ( .A(n86233), .Z(n105789) );
  INV_X1 U92644 ( .A(n82645), .ZN(n111122) );
  INV_X1 U92645 ( .A(n84054), .ZN(n106746) );
  CLKBUF_X1 U92646 ( .A(n58746), .Z(n106362) );
  INV_X1 U92647 ( .A(n82317), .ZN(n106823) );
  XNOR2_X1 U92648 ( .A(n82398), .B(n82394), .ZN(n82391) );
  INV_X1 U92649 ( .A(n100319), .ZN(n106846) );
  INV_X1 U92650 ( .A(n100232), .ZN(n106848) );
  INV_X1 U92651 ( .A(n82323), .ZN(n110442) );
  INV_X1 U92652 ( .A(n80119), .ZN(n106775) );
  INV_X1 U92653 ( .A(n80143), .ZN(n106790) );
  INV_X1 U92654 ( .A(n80115), .ZN(n106789) );
  INV_X1 U92655 ( .A(n80117), .ZN(n106788) );
  INV_X1 U92656 ( .A(n80129), .ZN(n106774) );
  INV_X1 U92657 ( .A(n80101), .ZN(n106792) );
  INV_X1 U92658 ( .A(n80131), .ZN(n106795) );
  INV_X1 U92659 ( .A(n80141), .ZN(n106794) );
  INV_X1 U92660 ( .A(n80139), .ZN(n106799) );
  INV_X1 U92661 ( .A(n80107), .ZN(n106798) );
  INV_X1 U92662 ( .A(n80109), .ZN(n106797) );
  INV_X1 U92663 ( .A(n80111), .ZN(n106796) );
  INV_X1 U92664 ( .A(n80113), .ZN(n106793) );
  CLKBUF_X1 U92665 ( .A(n82806), .Z(n105886) );
  CLKBUF_X1 U92666 ( .A(n98831), .Z(n105232) );
  XNOR2_X1 U92667 ( .A(n99334), .B(n82687), .ZN(n100314) );
  CLKBUF_X1 U92668 ( .A(n81280), .Z(n106240) );
  CLKBUF_X1 U92669 ( .A(n81342), .Z(n106167) );
  CLKBUF_X1 U92670 ( .A(n81472), .Z(n106060) );
  CLKBUF_X1 U92671 ( .A(n81567), .Z(n106019) );
  CLKBUF_X1 U92672 ( .A(n94536), .Z(n105626) );
  CLKBUF_X1 U92673 ( .A(n94544), .Z(n105623) );
  CLKBUF_X1 U92674 ( .A(n94546), .Z(n105622) );
  CLKBUF_X1 U92675 ( .A(n81783), .Z(n105911) );
  CLKBUF_X1 U92676 ( .A(n94548), .Z(n105621) );
  CLKBUF_X1 U92677 ( .A(n81472), .Z(n106061) );
  CLKBUF_X1 U92678 ( .A(n81567), .Z(n106020) );
  CLKBUF_X1 U92679 ( .A(n81280), .Z(n106241) );
  CLKBUF_X1 U92680 ( .A(n81342), .Z(n106168) );
  CLKBUF_X1 U92681 ( .A(n79980), .Z(n106348) );
  CLKBUF_X1 U92682 ( .A(n94544), .Z(n105624) );
  INV_X1 U92683 ( .A(n94852), .ZN(n107028) );
  INV_X1 U92684 ( .A(n82853), .ZN(n111052) );
  INV_X1 U92685 ( .A(n99323), .ZN(n106935) );
  INV_X1 U92686 ( .A(n90127), .ZN(n107123) );
  INV_X1 U92687 ( .A(n96130), .ZN(n106757) );
  INV_X1 U92688 ( .A(n82971), .ZN(n108625) );
  INV_X1 U92689 ( .A(n82886), .ZN(n111049) );
  INV_X1 U92690 ( .A(n82174), .ZN(n106782) );
  INV_X1 U92691 ( .A(n80146), .ZN(n106776) );
  INV_X1 U92692 ( .A(n80134), .ZN(n106791) );
  INV_X1 U92693 ( .A(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 [3]), .ZN(
        n106801) );
  INV_X1 U92694 ( .A(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 [2]), .ZN(
        n106802) );
  INV_X1 U92695 ( .A(\DLX_Datapath/TA_adder/P4_SumGen/CSel_i_0/S_0 [1]), .ZN(
        n106803) );
  INV_X1 U92696 ( .A(n104893), .ZN(n106777) );
  CLKBUF_X1 U92697 ( .A(n79980), .Z(n106349) );
  INV_X1 U92698 ( .A(n80122), .ZN(n106773) );
  INV_X1 U92699 ( .A(n82193), .ZN(n106781) );
  INV_X1 U92700 ( .A(n82187), .ZN(n106778) );
  INV_X1 U92701 ( .A(n82180), .ZN(n106779) );
  CLKBUF_X1 U92702 ( .A(n82805), .Z(n105144) );
  INV_X1 U92703 ( .A(n82056), .ZN(n106800) );
  CLKBUF_X1 U92704 ( .A(n81280), .Z(n106242) );
  CLKBUF_X1 U92705 ( .A(n81342), .Z(n106169) );
  CLKBUF_X1 U92706 ( .A(n81472), .Z(n106062) );
  CLKBUF_X1 U92707 ( .A(n81567), .Z(n106021) );
  CLKBUF_X1 U92708 ( .A(n94544), .Z(n105625) );
  INV_X1 U92709 ( .A(n99349), .ZN(n107061) );
  INV_X1 U92710 ( .A(n94068), .ZN(n107147) );
  INV_X1 U92711 ( .A(n82659), .ZN(n106805) );
  INV_X1 U92712 ( .A(n94081), .ZN(n107131) );
  INV_X1 U92713 ( .A(n90110), .ZN(n107140) );
  INV_X1 U92714 ( .A(n82405), .ZN(n107746) );
  INV_X1 U92715 ( .A(n95451), .ZN(n105502) );
  INV_X1 U92716 ( .A(n82278), .ZN(n106843) );
  INV_X1 U92717 ( .A(n82789), .ZN(n107160) );
  INV_X1 U92718 ( .A(n94732), .ZN(n106754) );
  INV_X1 U92719 ( .A(n82876), .ZN(n106831) );
  INV_X1 U92720 ( .A(n82318), .ZN(n108275) );
  INV_X1 U92721 ( .A(n82164), .ZN(n107745) );
  INV_X1 U92722 ( .A(n82328), .ZN(n110441) );
  INV_X1 U92723 ( .A(n100394), .ZN(n107060) );
  INV_X1 U92724 ( .A(n82597), .ZN(n106810) );
  INV_X1 U92725 ( .A(n82616), .ZN(n106811) );
  INV_X1 U92726 ( .A(n82600), .ZN(n106804) );
  INV_X1 U92727 ( .A(n83095), .ZN(n107062) );
  INV_X1 U92728 ( .A(n89977), .ZN(n111058) );
  INV_X1 U92729 ( .A(n104722), .ZN(n107103) );
  INV_X1 U92730 ( .A(n94730), .ZN(n106756) );
  INV_X1 U92731 ( .A(n94888), .ZN(n106755) );
  INV_X1 U92732 ( .A(n87620), .ZN(n107390) );
  INV_X1 U92733 ( .A(n87384), .ZN(n107386) );
  INV_X1 U92734 ( .A(n87738), .ZN(n107392) );
  INV_X1 U92735 ( .A(n87502), .ZN(n107388) );
  INV_X1 U92736 ( .A(n87974), .ZN(n107396) );
  INV_X1 U92737 ( .A(n87856), .ZN(n107394) );
  INV_X1 U92738 ( .A(n88092), .ZN(n107398) );
  INV_X1 U92739 ( .A(n88210), .ZN(n107400) );
  INV_X1 U92740 ( .A(n81794), .ZN(n107367) );
  INV_X1 U92741 ( .A(n88800), .ZN(n107410) );
  INV_X1 U92742 ( .A(n89153), .ZN(n107369) );
  INV_X1 U92743 ( .A(n81792), .ZN(n111063) );
  INV_X1 U92744 ( .A(n89506), .ZN(n111062) );
  INV_X1 U92745 ( .A(n89624), .ZN(n111061) );
  INV_X1 U92746 ( .A(n81790), .ZN(n111059) );
  INV_X1 U92747 ( .A(n89742), .ZN(n111060) );
  INV_X1 U92748 ( .A(n88918), .ZN(n107412) );
  INV_X1 U92749 ( .A(n88564), .ZN(n107406) );
  INV_X1 U92750 ( .A(n88446), .ZN(n107404) );
  INV_X1 U92751 ( .A(n88328), .ZN(n107402) );
  INV_X1 U92752 ( .A(n88682), .ZN(n107408) );
  INV_X1 U92753 ( .A(n90096), .ZN(n111057) );
  INV_X1 U92754 ( .A(n81968), .ZN(n111120) );
  INV_X1 U92755 ( .A(n83102), .ZN(n106880) );
  INV_X1 U92756 ( .A(n100324), .ZN(n106845) );
  INV_X1 U92757 ( .A(n82457), .ZN(n106821) );
  INV_X1 U92758 ( .A(n82484), .ZN(n106816) );
  INV_X1 U92759 ( .A(n82023), .ZN(n106772) );
  INV_X1 U92760 ( .A(n80072), .ZN(n106572) );
  INV_X1 U92761 ( .A(n82266), .ZN(n105080) );
  INV_X1 U92762 ( .A(
        \add_1_root_DLX_Datapath/TA_adder/P4_SumGen/CSel_i_4/RCA_1/add_38_2/carry[2] ), .ZN(n109782) );
  INV_X1 U92763 ( .A(n94483), .ZN(n106980) );
  INV_X1 U92764 ( .A(n94481), .ZN(n106982) );
  INV_X1 U92765 ( .A(n94484), .ZN(n106979) );
  INV_X1 U92766 ( .A(n94482), .ZN(n106981) );
  INV_X1 U92767 ( .A(n94486), .ZN(n106977) );
  INV_X1 U92768 ( .A(n94485), .ZN(n106978) );
  INV_X1 U92769 ( .A(n94487), .ZN(n106976) );
  INV_X1 U92770 ( .A(n94488), .ZN(n106975) );
  INV_X1 U92771 ( .A(n94495), .ZN(n106968) );
  INV_X1 U92772 ( .A(n94493), .ZN(n106970) );
  INV_X1 U92773 ( .A(n94496), .ZN(n106967) );
  INV_X1 U92774 ( .A(n94498), .ZN(n106965) );
  INV_X1 U92775 ( .A(n94499), .ZN(n106964) );
  INV_X1 U92776 ( .A(n94500), .ZN(n106963) );
  INV_X1 U92777 ( .A(n94502), .ZN(n106961) );
  INV_X1 U92778 ( .A(n94501), .ZN(n106962) );
  INV_X1 U92779 ( .A(n94494), .ZN(n106969) );
  INV_X1 U92780 ( .A(n94491), .ZN(n106972) );
  INV_X1 U92781 ( .A(n94490), .ZN(n106973) );
  INV_X1 U92782 ( .A(n94489), .ZN(n106974) );
  INV_X1 U92783 ( .A(n94492), .ZN(n106971) );
  INV_X1 U92784 ( .A(n94504), .ZN(n106959) );
  INV_X1 U92785 ( .A(n94344), .ZN(n107011) );
  INV_X1 U92786 ( .A(n94342), .ZN(n107013) );
  INV_X1 U92787 ( .A(n94345), .ZN(n107010) );
  INV_X1 U92788 ( .A(n94343), .ZN(n107012) );
  INV_X1 U92789 ( .A(n94347), .ZN(n107008) );
  INV_X1 U92790 ( .A(n94346), .ZN(n107009) );
  INV_X1 U92791 ( .A(n94348), .ZN(n107007) );
  INV_X1 U92792 ( .A(n94349), .ZN(n107006) );
  INV_X1 U92793 ( .A(n94356), .ZN(n106999) );
  INV_X1 U92794 ( .A(n94354), .ZN(n107001) );
  INV_X1 U92795 ( .A(n94357), .ZN(n106998) );
  INV_X1 U92796 ( .A(n94359), .ZN(n106996) );
  INV_X1 U92797 ( .A(n94360), .ZN(n106995) );
  INV_X1 U92798 ( .A(n94361), .ZN(n106994) );
  INV_X1 U92799 ( .A(n94363), .ZN(n106992) );
  INV_X1 U92800 ( .A(n94362), .ZN(n106993) );
  INV_X1 U92801 ( .A(n94355), .ZN(n107000) );
  INV_X1 U92802 ( .A(n94352), .ZN(n107003) );
  INV_X1 U92803 ( .A(n94351), .ZN(n107004) );
  INV_X1 U92804 ( .A(n94350), .ZN(n107005) );
  INV_X1 U92805 ( .A(n94353), .ZN(n107002) );
  INV_X1 U92806 ( .A(n94365), .ZN(n106990) );
  INV_X1 U92807 ( .A(n94503), .ZN(n106960) );
  INV_X1 U92808 ( .A(n94364), .ZN(n106991) );
  INV_X1 U92809 ( .A(n94497), .ZN(n106966) );
  INV_X1 U92810 ( .A(n94358), .ZN(n106997) );
  INV_X1 U92811 ( .A(n94480), .ZN(n106983) );
  INV_X1 U92812 ( .A(n94479), .ZN(n106984) );
  INV_X1 U92813 ( .A(n94477), .ZN(n106986) );
  INV_X1 U92814 ( .A(n94478), .ZN(n106985) );
  INV_X1 U92815 ( .A(n94474), .ZN(n106988) );
  INV_X1 U92816 ( .A(n94471), .ZN(n106989) );
  INV_X1 U92817 ( .A(n94476), .ZN(n106987) );
  INV_X1 U92818 ( .A(n94475), .ZN(n106833) );
  INV_X1 U92819 ( .A(n94341), .ZN(n107014) );
  INV_X1 U92820 ( .A(n94340), .ZN(n107015) );
  INV_X1 U92821 ( .A(n94338), .ZN(n107017) );
  INV_X1 U92822 ( .A(n94339), .ZN(n107016) );
  INV_X1 U92823 ( .A(n94335), .ZN(n107019) );
  INV_X1 U92824 ( .A(n94332), .ZN(n107020) );
  INV_X1 U92825 ( .A(n94337), .ZN(n107018) );
  INV_X1 U92826 ( .A(n94336), .ZN(n106834) );
  INV_X1 U92827 ( .A(n80088), .ZN(n106558) );
  OAI21_X1 U92828 ( .B1(n104807), .B2(n104734), .A(n80123), .ZN(n105053) );
  INV_X1 U92829 ( .A(n94083), .ZN(n107119) );
  INV_X1 U92830 ( .A(n90118), .ZN(n107121) );
  INV_X1 U92831 ( .A(n90115), .ZN(n107124) );
  INV_X1 U92832 ( .A(n99729), .ZN(n107440) );
  NOR2_X1 U92833 ( .A1(n90290), .A2(n90291), .ZN(n105054) );
  INV_X1 U92834 ( .A(n99808), .ZN(n107507) );
  INV_X1 U92835 ( .A(n99982), .ZN(n107537) );
  INV_X1 U92836 ( .A(n100013), .ZN(n107542) );
  INV_X1 U92837 ( .A(n99947), .ZN(n107533) );
  INV_X1 U92838 ( .A(n100045), .ZN(n107530) );
  INV_X1 U92839 ( .A(n99724), .ZN(n107452) );
  INV_X1 U92840 ( .A(n100100), .ZN(n107539) );
  INV_X1 U92841 ( .A(n99584), .ZN(n107463) );
  INV_X1 U92842 ( .A(n99577), .ZN(n107457) );
  INV_X1 U92843 ( .A(n99465), .ZN(n107460) );
  INV_X1 U92844 ( .A(n99558), .ZN(n107456) );
  INV_X1 U92845 ( .A(n99821), .ZN(n107495) );
  INV_X1 U92846 ( .A(n99748), .ZN(n107488) );
  INV_X1 U92847 ( .A(n99639), .ZN(n107443) );
  INV_X1 U92848 ( .A(n99420), .ZN(n107475) );
  INV_X1 U92849 ( .A(n99374), .ZN(n107478) );
  INV_X1 U92850 ( .A(\DLX_Datapath/ArithLogUnit/N179 ), .ZN(n106952) );
  INV_X1 U92851 ( .A(n99695), .ZN(n107433) );
  INV_X1 U92852 ( .A(n100113), .ZN(n107555) );
  INV_X1 U92853 ( .A(n99902), .ZN(n107526) );
  INV_X1 U92854 ( .A(n99770), .ZN(n107489) );
  INV_X1 U92855 ( .A(n99909), .ZN(n107509) );
  INV_X1 U92856 ( .A(n99862), .ZN(n107499) );
  INV_X1 U92857 ( .A(n99954), .ZN(n107512) );
  INV_X1 U92858 ( .A(n99989), .ZN(n107518) );
  INV_X1 U92859 ( .A(n99708), .ZN(n107445) );
  INV_X1 U92860 ( .A(n99608), .ZN(n107438) );
  INV_X1 U92861 ( .A(n90117), .ZN(n107125) );
  INV_X1 U92862 ( .A(n99520), .ZN(n107455) );
  INV_X1 U92863 ( .A(n99522), .ZN(n107521) );
  INV_X1 U92864 ( .A(n99439), .ZN(n107466) );
  INV_X1 U92865 ( .A(n99552), .ZN(n107462) );
  INV_X1 U92866 ( .A(n99670), .ZN(n107450) );
  INV_X1 U92867 ( .A(n99683), .ZN(n107540) );
  INV_X1 U92868 ( .A(n99682), .ZN(n107439) );
  INV_X1 U92869 ( .A(n99479), .ZN(n107473) );
  INV_X1 U92870 ( .A(n99569), .ZN(n107442) );
  INV_X1 U92871 ( .A(n99381), .ZN(n107559) );
  INV_X1 U92872 ( .A(n99882), .ZN(n107508) );
  INV_X1 U92873 ( .A(n99833), .ZN(n107498) );
  INV_X1 U92874 ( .A(n99038), .ZN(n107557) );
  INV_X1 U92875 ( .A(n99498), .ZN(n107464) );
  INV_X1 U92876 ( .A(n99676), .ZN(n107451) );
  INV_X1 U92877 ( .A(n100051), .ZN(n107528) );
  INV_X1 U92878 ( .A(n99599), .ZN(n107448) );
  INV_X1 U92879 ( .A(n99474), .ZN(n107467) );
  INV_X1 U92880 ( .A(n99871), .ZN(n107497) );
  INV_X1 U92881 ( .A(n99393), .ZN(n107474) );
  INV_X1 U92882 ( .A(n100023), .ZN(n107524) );
  INV_X1 U92883 ( .A(n99755), .ZN(n107496) );
  INV_X1 U92884 ( .A(n99534), .ZN(n107447) );
  INV_X1 U92885 ( .A(n99787), .ZN(n107493) );
  INV_X1 U92886 ( .A(n99935), .ZN(n107520) );
  INV_X1 U92887 ( .A(n99970), .ZN(n107525) );
  INV_X1 U92888 ( .A(n99890), .ZN(n107513) );
  INV_X1 U92889 ( .A(n100001), .ZN(n107529) );
  INV_X1 U92890 ( .A(n100066), .ZN(n107538) );
  INV_X1 U92891 ( .A(n99413), .ZN(n107506) );
  INV_X1 U92892 ( .A(n98978), .ZN(n106951) );
  INV_X1 U92893 ( .A(n99547), .ZN(n107468) );
  INV_X1 U92894 ( .A(n86272), .ZN(n107101) );
  INV_X1 U92895 ( .A(n99794), .ZN(n107494) );
  INV_X1 U92896 ( .A(n99702), .ZN(n107435) );
  INV_X1 U92897 ( .A(n99618), .ZN(n107449) );
  INV_X1 U92898 ( .A(n99841), .ZN(n107500) );
  INV_X1 U92899 ( .A(n99776), .ZN(n107487) );
  INV_X1 U92900 ( .A(n99739), .ZN(n107545) );
  INV_X1 U92901 ( .A(n99660), .ZN(n107483) );
  INV_X1 U92902 ( .A(n99856), .ZN(n107501) );
  INV_X1 U92903 ( .A(n106277), .ZN(n106275) );
  INV_X1 U92904 ( .A(n106277), .ZN(n106276) );
  INV_X1 U92905 ( .A(n99851), .ZN(n107569) );
  INV_X1 U92906 ( .A(n82006), .ZN(n111126) );
  XNOR2_X1 U92907 ( .A(n86297), .B(n100220), .ZN(n100273) );
  INV_X1 U92908 ( .A(n100170), .ZN(n108740) );
  INV_X1 U92909 ( .A(n100111), .ZN(n109086) );
  INV_X1 U92910 ( .A(n100020), .ZN(n108503) );
  INV_X1 U92911 ( .A(n99868), .ZN(n108271) );
  CLKBUF_X1 U92912 ( .A(n90305), .Z(n105656) );
  CLKBUF_X1 U92913 ( .A(n86317), .Z(n105783) );
  CLKBUF_X1 U92914 ( .A(n90302), .Z(n105658) );
  CLKBUF_X1 U92915 ( .A(n86310), .Z(n105786) );
  CLKBUF_X1 U92916 ( .A(n79716), .Z(n106356) );
  CLKBUF_X1 U92917 ( .A(n79714), .Z(n106357) );
  INV_X1 U92918 ( .A(n82400), .ZN(n111135) );
  CLKBUF_X1 U92919 ( .A(n90312), .Z(n105652) );
  CLKBUF_X1 U92920 ( .A(n90310), .Z(n105653) );
  CLKBUF_X1 U92921 ( .A(n86320), .Z(n105780) );
  CLKBUF_X1 U92922 ( .A(n86314), .Z(n105784) );
  CLKBUF_X1 U92923 ( .A(n99849), .Z(n105102) );
  XOR2_X1 U92924 ( .A(\DLX_Datapath/RegisterFile/N27074 ), .B(n104328), .Z(
        n105055) );
  XOR2_X1 U92925 ( .A(\DLX_Datapath/RegisterFile/N27074 ), .B(n104328), .Z(
        n105056) );
  XOR2_X1 U92926 ( .A(\DLX_Datapath/RegisterFile/N27074 ), .B(n104328), .Z(
        n105057) );
  INV_X1 U92927 ( .A(n81974), .ZN(n111124) );
  INV_X1 U92928 ( .A(n80064), .ZN(n111147) );
  XOR2_X1 U92929 ( .A(\DLX_Datapath/RegisterFile/N27074 ), .B(n104328), .Z(
        n105058) );
  INV_X1 U92930 ( .A(n82624), .ZN(n111128) );
  INV_X1 U92931 ( .A(n79821), .ZN(n107582) );
  INV_X1 U92932 ( .A(n79920), .ZN(n107615) );
  INV_X1 U92933 ( .A(n79887), .ZN(n107609) );
  INV_X1 U92934 ( .A(n99235), .ZN(n107428) );
  INV_X1 U92935 ( .A(n99270), .ZN(n107430) );
  INV_X1 U92936 ( .A(n99281), .ZN(n107549) );
  INV_X1 U92937 ( .A(n99198), .ZN(n107511) );
  INV_X1 U92938 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [25]), .ZN(n106872) );
  INV_X1 U92939 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [24]), .ZN(n106871) );
  INV_X1 U92940 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [27]), .ZN(n106874) );
  INV_X1 U92941 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [21]), .ZN(n106868) );
  INV_X1 U92942 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [23]), .ZN(n106870) );
  INV_X1 U92943 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [20]), .ZN(n106867) );
  INV_X1 U92944 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [22]), .ZN(n106869) );
  INV_X1 U92945 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [18]), .ZN(n106865) );
  INV_X1 U92946 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [19]), .ZN(n106866) );
  INV_X1 U92947 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [17]), .ZN(n106864) );
  INV_X1 U92948 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [16]), .ZN(n106863) );
  INV_X1 U92949 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [15]), .ZN(n106862) );
  INV_X1 U92950 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [26]), .ZN(n106873) );
  INV_X1 U92951 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [14]), .ZN(n106861) );
  INV_X1 U92952 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [13]), .ZN(n106860) );
  INV_X1 U92953 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [12]), .ZN(n106859) );
  INV_X1 U92954 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [10]), .ZN(n106857) );
  INV_X1 U92955 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [9]), .ZN(n106856) );
  INV_X1 U92956 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [8]), .ZN(n106855) );
  INV_X1 U92957 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [6]), .ZN(n106853) );
  INV_X1 U92958 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [5]), .ZN(n106852) );
  INV_X1 U92959 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [7]), .ZN(n106854) );
  INV_X1 U92960 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [11]), .ZN(n106858) );
  INV_X1 U92961 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [28]), .ZN(n106875) );
  CLKBUF_X1 U92962 ( .A(n99449), .Z(n105115) );
  INV_X1 U92963 ( .A(n79854), .ZN(n107604) );
  INV_X1 U92964 ( .A(n79720), .ZN(n107591) );
  INV_X1 U92965 ( .A(n99253), .ZN(n107429) );
  INV_X1 U92966 ( .A(n99090), .ZN(n107459) );
  INV_X1 U92967 ( .A(n99130), .ZN(n107441) );
  INV_X1 U92968 ( .A(n99120), .ZN(n107535) );
  INV_X1 U92969 ( .A(n99110), .ZN(n107532) );
  INV_X1 U92970 ( .A(n99169), .ZN(n107485) );
  INV_X1 U92971 ( .A(n99160), .ZN(n107431) );
  INV_X1 U92972 ( .A(n99150), .ZN(n107432) );
  INV_X1 U92973 ( .A(n99050), .ZN(n107477) );
  INV_X1 U92974 ( .A(n99070), .ZN(n107470) );
  INV_X1 U92975 ( .A(n81812), .ZN(n107491) );
  INV_X1 U92976 ( .A(n79755), .ZN(n107596) );
  INV_X1 U92977 ( .A(n99140), .ZN(n107436) );
  INV_X1 U92978 ( .A(n99060), .ZN(n107505) );
  CLKBUF_X1 U92979 ( .A(n94111), .Z(n105139) );
  CLKBUF_X1 U92980 ( .A(n94114), .Z(n105138) );
  CLKBUF_X1 U92981 ( .A(n94112), .Z(n105141) );
  INV_X1 U92982 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [2]), .ZN(n106850) );
  INV_X1 U92983 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [1]), .ZN(n106849) );
  INV_X1 U92984 ( .A(\DLX_Datapath/MUX_HDU_ALUInA [3]), .ZN(n106851) );
  INV_X1 U92985 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [0]), .ZN(n106768) );
  INV_X1 U92986 ( .A(n81804), .ZN(n105900) );
  INV_X1 U92987 ( .A(n81975), .ZN(n111148) );
  INV_X1 U92988 ( .A(n82407), .ZN(n111131) );
  INV_X1 U92989 ( .A(n85154), .ZN(n106701) );
  INV_X1 U92990 ( .A(n85121), .ZN(n106702) );
  INV_X1 U92991 ( .A(n85088), .ZN(n106703) );
  INV_X1 U92992 ( .A(n85055), .ZN(n106704) );
  INV_X1 U92993 ( .A(n85022), .ZN(n106705) );
  INV_X1 U92994 ( .A(n84989), .ZN(n106706) );
  INV_X1 U92995 ( .A(n84956), .ZN(n106707) );
  INV_X1 U92996 ( .A(n84923), .ZN(n106708) );
  INV_X1 U92997 ( .A(n84890), .ZN(n106709) );
  INV_X1 U92998 ( .A(n84857), .ZN(n106710) );
  INV_X1 U92999 ( .A(n84824), .ZN(n106711) );
  INV_X1 U93000 ( .A(n84791), .ZN(n106712) );
  INV_X1 U93001 ( .A(n84758), .ZN(n106713) );
  INV_X1 U93002 ( .A(n84725), .ZN(n106714) );
  INV_X1 U93003 ( .A(n84692), .ZN(n106715) );
  INV_X1 U93004 ( .A(n84659), .ZN(n106716) );
  INV_X1 U93005 ( .A(n84626), .ZN(n106717) );
  INV_X1 U93006 ( .A(n84593), .ZN(n106718) );
  INV_X1 U93007 ( .A(n84560), .ZN(n106719) );
  INV_X1 U93008 ( .A(n84527), .ZN(n106720) );
  INV_X1 U93009 ( .A(n84494), .ZN(n106721) );
  INV_X1 U93010 ( .A(n84461), .ZN(n106722) );
  INV_X1 U93011 ( .A(n84428), .ZN(n106723) );
  INV_X1 U93012 ( .A(n84395), .ZN(n106724) );
  INV_X1 U93013 ( .A(n84362), .ZN(n106725) );
  INV_X1 U93014 ( .A(n84329), .ZN(n106726) );
  INV_X1 U93015 ( .A(n84296), .ZN(n106727) );
  INV_X1 U93016 ( .A(n84263), .ZN(n106728) );
  INV_X1 U93017 ( .A(n84230), .ZN(n106729) );
  INV_X1 U93018 ( .A(n84197), .ZN(n106730) );
  INV_X1 U93019 ( .A(n84164), .ZN(n106731) );
  INV_X1 U93020 ( .A(n84097), .ZN(n106732) );
  INV_X1 U93021 ( .A(n99344), .ZN(n107102) );
  INV_X1 U93022 ( .A(n98977), .ZN(n110957) );
  INV_X1 U93023 ( .A(n82636), .ZN(n111139) );
  INV_X1 U93024 ( .A(n105064), .ZN(
        \add_0_root_add_0_root_DLX_Datapath/RegisterFile/add_243_3/carry[6] )
         );
  INV_X1 U93025 ( .A(n82303), .ZN(n111133) );
  INV_X1 U93026 ( .A(n79797), .ZN(n106911) );
  INV_X1 U93027 ( .A(n79789), .ZN(n106913) );
  INV_X1 U93028 ( .A(n79780), .ZN(n106915) );
  INV_X1 U93029 ( .A(n79830), .ZN(n106905) );
  INV_X1 U93030 ( .A(n79822), .ZN(n106907) );
  INV_X1 U93031 ( .A(n79813), .ZN(n106909) );
  INV_X1 U93032 ( .A(n79896), .ZN(n106893) );
  INV_X1 U93033 ( .A(n79929), .ZN(n106887) );
  INV_X1 U93034 ( .A(n79921), .ZN(n106889) );
  INV_X1 U93035 ( .A(n79912), .ZN(n106891) );
  INV_X1 U93036 ( .A(n79953), .ZN(n106883) );
  INV_X1 U93037 ( .A(n79961), .ZN(n106881) );
  INV_X1 U93038 ( .A(n79945), .ZN(n106885) );
  INV_X1 U93039 ( .A(n79888), .ZN(n106895) );
  INV_X1 U93040 ( .A(n79879), .ZN(n106897) );
  INV_X1 U93041 ( .A(n79863), .ZN(n106899) );
  INV_X1 U93042 ( .A(n79855), .ZN(n106901) );
  INV_X1 U93043 ( .A(n79846), .ZN(n106903) );
  INV_X1 U93044 ( .A(n79764), .ZN(n106917) );
  INV_X1 U93045 ( .A(n79756), .ZN(n106919) );
  INV_X1 U93046 ( .A(n79747), .ZN(n106921) );
  INV_X1 U93047 ( .A(n79721), .ZN(n106923) );
  INV_X1 U93048 ( .A(n79706), .ZN(n106925) );
  INV_X1 U93049 ( .A(n79729), .ZN(n106839) );
  INV_X1 U93050 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [2]), .ZN(n106884) );
  INV_X1 U93051 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [1]), .ZN(n106882) );
  INV_X1 U93052 ( .A(n100231), .ZN(n106931) );
  INV_X1 U93053 ( .A(n98971), .ZN(n106950) );
  INV_X1 U93054 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [31]), .ZN(n106926) );
  INV_X1 U93055 ( .A(n94065), .ZN(n107146) );
  INV_X1 U93056 ( .A(n90109), .ZN(n107120) );
  INV_X1 U93057 ( .A(n80091), .ZN(n111119) );
  INV_X1 U93058 ( .A(n82770), .ZN(n111129) );
  INV_X1 U93059 ( .A(n99326), .ZN(n106938) );
  INV_X1 U93060 ( .A(n100061), .ZN(n109090) );
  INV_X1 U93061 ( .A(n99924), .ZN(n107738) );
  INV_X1 U93062 ( .A(n98973), .ZN(n106947) );
  INV_X1 U93063 ( .A(n100144), .ZN(n108743) );
  INV_X1 U93064 ( .A(n99901), .ZN(n107516) );
  INV_X1 U93065 ( .A(n100012), .ZN(n107534) );
  INV_X1 U93066 ( .A(n99946), .ZN(n107523) );
  INV_X1 U93067 ( .A(n99981), .ZN(n107527) );
  INV_X1 U93068 ( .A(n99217), .ZN(n107427) );
  INV_X1 U93069 ( .A(n100078), .ZN(n107543) );
  INV_X1 U93070 ( .A(n99180), .ZN(n107425) );
  INV_X1 U93071 ( .A(n99753), .ZN(n107522) );
  INV_X1 U93072 ( .A(n99668), .ZN(n107510) );
  INV_X1 U93073 ( .A(n99933), .ZN(n107541) );
  INV_X1 U93074 ( .A(n99999), .ZN(n107546) );
  INV_X1 U93075 ( .A(n100064), .ZN(n107554) );
  INV_X1 U93076 ( .A(n99968), .ZN(n107544) );
  INV_X1 U93077 ( .A(n99888), .ZN(n107536) );
  INV_X1 U93078 ( .A(n99987), .ZN(n107550) );
  INV_X1 U93079 ( .A(n100079), .ZN(n107547) );
  INV_X1 U93080 ( .A(n99807), .ZN(n107515) );
  INV_X1 U93081 ( .A(n100112), .ZN(n107548) );
  INV_X1 U93082 ( .A(n99927), .ZN(n107553) );
  INV_X1 U93083 ( .A(n99080), .ZN(n107514) );
  INV_X1 U93084 ( .A(n99170), .ZN(n107552) );
  INV_X1 U93085 ( .A(n99199), .ZN(n107426) );
  INV_X1 U93086 ( .A(n105123), .ZN(n106954) );
  INV_X1 U93087 ( .A(n99504), .ZN(n107504) );
  INV_X1 U93088 ( .A(n99452), .ZN(n107503) );
  INV_X1 U93089 ( .A(n81962), .ZN(n111161) );
  INV_X1 U93090 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [3]), .ZN(n106886) );
  INV_X1 U93091 ( .A(n79697), .ZN(n107585) );
  INV_X1 U93092 ( .A(n79694), .ZN(n107581) );
  INV_X1 U93093 ( .A(n79703), .ZN(n107590) );
  INV_X1 U93094 ( .A(n79691), .ZN(n107603) );
  INV_X1 U93095 ( .A(n79688), .ZN(n107608) );
  INV_X1 U93096 ( .A(n79685), .ZN(n107614) );
  INV_X1 U93097 ( .A(n79700), .ZN(n107595) );
  INV_X1 U93098 ( .A(n79684), .ZN(n107577) );
  INV_X1 U93099 ( .A(n79683), .ZN(n107576) );
  INV_X1 U93100 ( .A(n79682), .ZN(n107575) );
  INV_X1 U93101 ( .A(n82332), .ZN(n111130) );
  INV_X1 U93102 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [9]), .ZN(n106894) );
  INV_X1 U93103 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [5]), .ZN(n106888) );
  INV_X1 U93104 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [6]), .ZN(n106890) );
  INV_X1 U93105 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [7]), .ZN(n106892) );
  INV_X1 U93106 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [10]), .ZN(n106896) );
  INV_X1 U93107 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [11]), .ZN(n106898) );
  INV_X1 U93108 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [13]), .ZN(n106900) );
  INV_X1 U93109 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [14]), .ZN(n106902) );
  INV_X1 U93110 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [15]), .ZN(n106904) );
  INV_X1 U93111 ( .A(n81966), .ZN(n111157) );
  INV_X1 U93112 ( .A(n84095), .ZN(n106745) );
  INV_X1 U93113 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [21]), .ZN(n106912) );
  INV_X1 U93114 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [22]), .ZN(n106914) );
  INV_X1 U93115 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [23]), .ZN(n106916) );
  INV_X1 U93116 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [17]), .ZN(n106906) );
  INV_X1 U93117 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [18]), .ZN(n106908) );
  INV_X1 U93118 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [19]), .ZN(n106910) );
  INV_X1 U93119 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [25]), .ZN(n106918) );
  INV_X1 U93120 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [26]), .ZN(n106920) );
  INV_X1 U93121 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [27]), .ZN(n106922) );
  INV_X1 U93122 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [30]), .ZN(n106924) );
  INV_X1 U93123 ( .A(\DLX_Datapath/MUX_HDU_ALUInB [29]), .ZN(n106840) );
  INV_X1 U93124 ( .A(n99271), .ZN(n107551) );
  INV_X1 U93125 ( .A(n81809), .ZN(n106877) );
  INV_X1 U93126 ( .A(n81802), .ZN(n106841) );
  INV_X1 U93127 ( .A(n81813), .ZN(n106876) );
  INV_X1 U93128 ( .A(n87619), .ZN(n107049) );
  INV_X1 U93129 ( .A(n91602), .ZN(n107083) );
  INV_X1 U93130 ( .A(n87383), .ZN(n107051) );
  INV_X1 U93131 ( .A(n91368), .ZN(n107085) );
  INV_X1 U93132 ( .A(n87737), .ZN(n107048) );
  INV_X1 U93133 ( .A(n91719), .ZN(n107082) );
  INV_X1 U93134 ( .A(n87501), .ZN(n107050) );
  INV_X1 U93135 ( .A(n91485), .ZN(n107084) );
  INV_X1 U93136 ( .A(n87973), .ZN(n107046) );
  INV_X1 U93137 ( .A(n91953), .ZN(n107080) );
  INV_X1 U93138 ( .A(n87855), .ZN(n107047) );
  INV_X1 U93139 ( .A(n91836), .ZN(n107081) );
  INV_X1 U93140 ( .A(n88091), .ZN(n107045) );
  INV_X1 U93141 ( .A(n92070), .ZN(n107079) );
  INV_X1 U93142 ( .A(n88209), .ZN(n107044) );
  INV_X1 U93143 ( .A(n92187), .ZN(n107078) );
  INV_X1 U93144 ( .A(n88917), .ZN(n107038) );
  INV_X1 U93145 ( .A(n89035), .ZN(n107037) );
  INV_X1 U93146 ( .A(n93006), .ZN(n107071) );
  INV_X1 U93147 ( .A(n88799), .ZN(n107039) );
  INV_X1 U93148 ( .A(n92772), .ZN(n107073) );
  INV_X1 U93149 ( .A(n89152), .ZN(n107036) );
  INV_X1 U93150 ( .A(n93123), .ZN(n107070) );
  INV_X1 U93151 ( .A(n89388), .ZN(n107034) );
  INV_X1 U93152 ( .A(n93357), .ZN(n107068) );
  INV_X1 U93153 ( .A(n89505), .ZN(n107033) );
  INV_X1 U93154 ( .A(n93474), .ZN(n107067) );
  INV_X1 U93155 ( .A(n89623), .ZN(n107032) );
  INV_X1 U93156 ( .A(n93591), .ZN(n107066) );
  INV_X1 U93157 ( .A(n89859), .ZN(n107030) );
  INV_X1 U93158 ( .A(n93825), .ZN(n107064) );
  INV_X1 U93159 ( .A(n89741), .ZN(n107031) );
  INV_X1 U93160 ( .A(n93708), .ZN(n107065) );
  INV_X1 U93161 ( .A(n92889), .ZN(n107072) );
  INV_X1 U93162 ( .A(n88563), .ZN(n107041) );
  INV_X1 U93163 ( .A(n92538), .ZN(n107075) );
  INV_X1 U93164 ( .A(n88445), .ZN(n107042) );
  INV_X1 U93165 ( .A(n92421), .ZN(n107076) );
  INV_X1 U93166 ( .A(n88327), .ZN(n107043) );
  INV_X1 U93167 ( .A(n92304), .ZN(n107077) );
  INV_X1 U93168 ( .A(n88681), .ZN(n107040) );
  INV_X1 U93169 ( .A(n92655), .ZN(n107074) );
  INV_X1 U93170 ( .A(n89976), .ZN(n107029) );
  INV_X1 U93171 ( .A(n93942), .ZN(n107063) );
  INV_X1 U93172 ( .A(n87265), .ZN(n107052) );
  INV_X1 U93173 ( .A(n91251), .ZN(n107086) );
  INV_X1 U93174 ( .A(n87147), .ZN(n107053) );
  INV_X1 U93175 ( .A(n91134), .ZN(n107087) );
  INV_X1 U93176 ( .A(n86911), .ZN(n107055) );
  INV_X1 U93177 ( .A(n90900), .ZN(n107089) );
  INV_X1 U93178 ( .A(n89270), .ZN(n107035) );
  INV_X1 U93179 ( .A(n93240), .ZN(n107069) );
  INV_X1 U93180 ( .A(n87029), .ZN(n107054) );
  INV_X1 U93181 ( .A(n91017), .ZN(n107088) );
  INV_X1 U93182 ( .A(n86557), .ZN(n107057) );
  INV_X1 U93183 ( .A(n90549), .ZN(n107091) );
  INV_X1 U93184 ( .A(n86301), .ZN(n107058) );
  INV_X1 U93185 ( .A(n90294), .ZN(n107092) );
  INV_X1 U93186 ( .A(n86793), .ZN(n107056) );
  INV_X1 U93187 ( .A(n90783), .ZN(n107090) );
  INV_X1 U93188 ( .A(n90666), .ZN(n106835) );
  INV_X1 U93189 ( .A(n86675), .ZN(n106836) );
  AND2_X2 U93190 ( .A1(n105059), .A2(n105060), .ZN(n98944) );
  INV_X1 U93191 ( .A(n80016), .ZN(n106673) );
  INV_X1 U93192 ( .A(n80017), .ZN(n106672) );
  INV_X1 U93193 ( .A(n80020), .ZN(n106669) );
  INV_X1 U93194 ( .A(n80021), .ZN(n106668) );
  INV_X1 U93195 ( .A(n80022), .ZN(n106667) );
  INV_X1 U93196 ( .A(n80023), .ZN(n106666) );
  INV_X1 U93197 ( .A(n80025), .ZN(n106664) );
  INV_X1 U93198 ( .A(n80024), .ZN(n106665) );
  INV_X1 U93199 ( .A(n80018), .ZN(n106671) );
  INV_X1 U93200 ( .A(n80019), .ZN(n106670) );
  INV_X1 U93201 ( .A(n80007), .ZN(n106682) );
  INV_X1 U93202 ( .A(n80006), .ZN(n106683) );
  INV_X1 U93203 ( .A(n80004), .ZN(n106685) );
  INV_X1 U93204 ( .A(n80010), .ZN(n106679) );
  INV_X1 U93205 ( .A(n80008), .ZN(n106681) );
  INV_X1 U93206 ( .A(n80011), .ZN(n106678) );
  INV_X1 U93207 ( .A(n80009), .ZN(n106680) );
  INV_X1 U93208 ( .A(n80012), .ZN(n106677) );
  INV_X1 U93209 ( .A(n80013), .ZN(n106676) );
  INV_X1 U93210 ( .A(n80014), .ZN(n106675) );
  INV_X1 U93211 ( .A(n80005), .ZN(n106684) );
  INV_X1 U93212 ( .A(n80015), .ZN(n106674) );
  INV_X1 U93213 ( .A(n80026), .ZN(n106663) );
  INV_X1 U93214 ( .A(n80003), .ZN(n106686) );
  INV_X1 U93215 ( .A(n79983), .ZN(n106659) );
  INV_X1 U93216 ( .A(n79987), .ZN(n106655) );
  INV_X1 U93217 ( .A(n79988), .ZN(n106654) );
  INV_X1 U93218 ( .A(n79986), .ZN(n106656) );
  INV_X1 U93219 ( .A(n79985), .ZN(n106657) );
  INV_X1 U93220 ( .A(n79982), .ZN(n106660) );
  INV_X1 U93221 ( .A(n79984), .ZN(n106658) );
  INV_X1 U93222 ( .A(n79981), .ZN(n106661) );
  INV_X1 U93223 ( .A(n79978), .ZN(n106662) );
  INV_X1 U93224 ( .A(n100347), .ZN(n106932) );
  INV_X1 U93225 ( .A(n79969), .ZN(n106694) );
  INV_X1 U93226 ( .A(n79975), .ZN(n106690) );
  INV_X1 U93227 ( .A(n79974), .ZN(n106691) );
  INV_X1 U93228 ( .A(n79976), .ZN(n106689) );
  INV_X1 U93229 ( .A(n79973), .ZN(n106692) );
  INV_X1 U93230 ( .A(n79972), .ZN(n106693) );
  INV_X1 U93231 ( .A(n79977), .ZN(n106688) );
  INV_X1 U93232 ( .A(n80002), .ZN(n106687) );
  INV_X1 U93233 ( .A(n82496), .ZN(n106814) );
  INV_X1 U93234 ( .A(n82788), .ZN(n107155) );
  INV_X1 U93235 ( .A(n82961), .ZN(n108626) );
  INV_X1 U93236 ( .A(n82991), .ZN(n108630) );
  INV_X1 U93237 ( .A(n82868), .ZN(n107630) );
  INV_X1 U93238 ( .A(n100362), .ZN(n107141) );
  XOR2_X1 U93239 ( .A(\DLX_Datapath/HazardDetUnit/N111 ), .B(n105061), .Z(
        n100385) );
  CLKBUF_X1 U93240 ( .A(n62189), .Z(n106358) );
  CLKBUF_X1 U93241 ( .A(n100414), .Z(n105222) );
  INV_X1 U93242 ( .A(n82977), .ZN(n108623) );
  CLKBUF_X1 U93243 ( .A(n100417), .Z(n105221) );
  INV_X1 U93244 ( .A(n105031), .ZN(n107099) );
  INV_X1 U93245 ( .A(n80150), .ZN(n106784) );
  INV_X1 U93246 ( .A(n82904), .ZN(n107158) );
  INV_X1 U93247 ( .A(n81887), .ZN(n111140) );
  INV_X1 U93248 ( .A(n80148), .ZN(n106787) );
  INV_X1 U93249 ( .A(n80128), .ZN(n106785) );
  INV_X1 U93250 ( .A(n80106), .ZN(n106786) );
  INV_X1 U93251 ( .A(n100228), .ZN(n106933) );
  INV_X1 U93252 ( .A(n80038), .ZN(n106598) );
  INV_X1 U93253 ( .A(n82627), .ZN(n106596) );
  INV_X1 U93254 ( .A(n100310), .ZN(n106762) );
  NAND2_X1 U93255 ( .A1(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_5/S_0 [0]), 
        .A2(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_4/S_0 [3]), .ZN(n105062)
         );
  CLKBUF_X1 U93256 ( .A(net2465245), .Z(n105075) );
  INV_X1 U93257 ( .A(n100256), .ZN(n106939) );
  NOR2_X1 U93258 ( .A1(n82458), .A2(n62199), .ZN(n105063) );
  INV_X1 U93259 ( .A(n83076), .ZN(n107157) );
  INV_X1 U93260 ( .A(n83051), .ZN(n107165) );
  INV_X1 U93261 ( .A(n83015), .ZN(n107626) );
  INV_X1 U93262 ( .A(n82914), .ZN(n107629) );
  INV_X1 U93263 ( .A(n82915), .ZN(n107627) );
  INV_X1 U93264 ( .A(n83043), .ZN(n107164) );
  INV_X1 U93265 ( .A(n83042), .ZN(n107162) );
  INV_X1 U93266 ( .A(n83029), .ZN(n107625) );
  INV_X1 U93267 ( .A(n83030), .ZN(n107623) );
  INV_X1 U93268 ( .A(n82938), .ZN(n108629) );
  INV_X1 U93269 ( .A(n82937), .ZN(n108627) );
  INV_X1 U93270 ( .A(n80068), .ZN(n106574) );
  INV_X1 U93271 ( .A(n80087), .ZN(n106559) );
  INV_X1 U93272 ( .A(n80062), .ZN(n106576) );
  INV_X1 U93273 ( .A(n80070), .ZN(n106573) );
  INV_X1 U93274 ( .A(n80055), .ZN(n106582) );
  INV_X1 U93275 ( .A(n80054), .ZN(n106583) );
  INV_X1 U93276 ( .A(n80053), .ZN(n106584) );
  INV_X1 U93277 ( .A(n80063), .ZN(n106575) );
  INV_X1 U93278 ( .A(n80052), .ZN(n106585) );
  INV_X1 U93279 ( .A(n80081), .ZN(n106564) );
  INV_X1 U93280 ( .A(n80051), .ZN(n106586) );
  INV_X1 U93281 ( .A(n80050), .ZN(n106587) );
  INV_X1 U93282 ( .A(n80049), .ZN(n106588) );
  INV_X1 U93283 ( .A(n80048), .ZN(n106589) );
  INV_X1 U93284 ( .A(n80047), .ZN(n106590) );
  INV_X1 U93285 ( .A(n80079), .ZN(n106566) );
  INV_X1 U93286 ( .A(n80046), .ZN(n106591) );
  INV_X1 U93287 ( .A(n80061), .ZN(n106577) );
  INV_X1 U93288 ( .A(n80078), .ZN(n106567) );
  INV_X1 U93289 ( .A(n80077), .ZN(n106568) );
  INV_X1 U93290 ( .A(n80060), .ZN(n106578) );
  INV_X1 U93291 ( .A(n80059), .ZN(n106579) );
  INV_X1 U93292 ( .A(n80076), .ZN(n106569) );
  INV_X1 U93293 ( .A(n80075), .ZN(n106570) );
  INV_X1 U93294 ( .A(n80045), .ZN(n106592) );
  INV_X1 U93295 ( .A(n80044), .ZN(n106593) );
  INV_X1 U93296 ( .A(n80074), .ZN(n106571) );
  INV_X1 U93297 ( .A(n80085), .ZN(n106560) );
  INV_X1 U93298 ( .A(n80095), .ZN(n106555) );
  INV_X1 U93299 ( .A(n80089), .ZN(n106557) );
  INV_X1 U93300 ( .A(n80084), .ZN(n106561) );
  INV_X1 U93301 ( .A(n80083), .ZN(n106562) );
  INV_X1 U93302 ( .A(n80082), .ZN(n106563) );
  INV_X1 U93303 ( .A(n80080), .ZN(n106565) );
  INV_X1 U93304 ( .A(n80043), .ZN(n106594) );
  INV_X1 U93305 ( .A(n82245), .ZN(n105066) );
  INV_X1 U93306 ( .A(n80172), .ZN(n106611) );
  INV_X1 U93307 ( .A(n80171), .ZN(n106612) );
  INV_X1 U93308 ( .A(n80173), .ZN(n106610) );
  INV_X1 U93309 ( .A(n80174), .ZN(n106609) );
  INV_X1 U93310 ( .A(n80161), .ZN(n106622) );
  INV_X1 U93311 ( .A(n80175), .ZN(n106608) );
  INV_X1 U93312 ( .A(n80179), .ZN(n106604) );
  INV_X1 U93313 ( .A(n80164), .ZN(n106619) );
  INV_X1 U93314 ( .A(n80165), .ZN(n106618) );
  INV_X1 U93315 ( .A(n80166), .ZN(n106617) );
  INV_X1 U93316 ( .A(n80181), .ZN(n106602) );
  INV_X1 U93317 ( .A(n80167), .ZN(n106616) );
  INV_X1 U93318 ( .A(n80180), .ZN(n106603) );
  INV_X1 U93319 ( .A(n80168), .ZN(n106615) );
  INV_X1 U93320 ( .A(n80183), .ZN(n106600) );
  INV_X1 U93321 ( .A(n80182), .ZN(n106601) );
  INV_X1 U93322 ( .A(n80178), .ZN(n106605) );
  INV_X1 U93323 ( .A(n80177), .ZN(n106606) );
  INV_X1 U93324 ( .A(n80176), .ZN(n106607) );
  INV_X1 U93325 ( .A(n80162), .ZN(n106621) );
  INV_X1 U93326 ( .A(n80169), .ZN(n106614) );
  INV_X1 U93327 ( .A(n80170), .ZN(n106613) );
  INV_X1 U93328 ( .A(n80163), .ZN(n106620) );
  INV_X1 U93329 ( .A(n80184), .ZN(n106599) );
  INV_X1 U93330 ( .A(n80037), .ZN(n106631) );
  INV_X1 U93331 ( .A(n79989), .ZN(n106653) );
  INV_X1 U93332 ( .A(n79991), .ZN(n106651) );
  INV_X1 U93333 ( .A(n79990), .ZN(n106652) );
  INV_X1 U93334 ( .A(n80028), .ZN(n106640) );
  INV_X1 U93335 ( .A(n80027), .ZN(n106641) );
  INV_X1 U93336 ( .A(n79993), .ZN(n106649) );
  INV_X1 U93337 ( .A(n79992), .ZN(n106650) );
  INV_X1 U93338 ( .A(n79995), .ZN(n106647) );
  INV_X1 U93339 ( .A(n79994), .ZN(n106648) );
  INV_X1 U93340 ( .A(n79999), .ZN(n106643) );
  INV_X1 U93341 ( .A(n79998), .ZN(n106644) );
  INV_X1 U93342 ( .A(n80000), .ZN(n106642) );
  INV_X1 U93343 ( .A(n79997), .ZN(n106645) );
  INV_X1 U93344 ( .A(n79996), .ZN(n106646) );
  INV_X1 U93345 ( .A(n80030), .ZN(n106638) );
  INV_X1 U93346 ( .A(n80031), .ZN(n106637) );
  INV_X1 U93347 ( .A(n80034), .ZN(n106634) );
  INV_X1 U93348 ( .A(n80035), .ZN(n106633) );
  INV_X1 U93349 ( .A(n80036), .ZN(n106632) );
  INV_X1 U93350 ( .A(n80032), .ZN(n106636) );
  INV_X1 U93351 ( .A(n80033), .ZN(n106635) );
  INV_X1 U93352 ( .A(n80029), .ZN(n106639) );
  INV_X1 U93353 ( .A(n80156), .ZN(n106627) );
  INV_X1 U93354 ( .A(n80158), .ZN(n106625) );
  INV_X1 U93355 ( .A(n80159), .ZN(n106624) );
  INV_X1 U93356 ( .A(n80157), .ZN(n106626) );
  INV_X1 U93357 ( .A(n80160), .ZN(n106623) );
  INV_X1 U93358 ( .A(n80155), .ZN(n106628) );
  INV_X1 U93359 ( .A(n80151), .ZN(n106630) );
  INV_X1 U93360 ( .A(n80154), .ZN(n106629) );
  INV_X1 U93361 ( .A(n80058), .ZN(n106580) );
  INV_X1 U93362 ( .A(n80057), .ZN(n106581) );
  INV_X1 U93363 ( .A(n80090), .ZN(n106556) );
  INV_X1 U93364 ( .A(n82008), .ZN(n106554) );
  INV_X1 U93365 ( .A(n100403), .ZN(n107094) );
  INV_X1 U93366 ( .A(n81847), .ZN(n107599) );
  INV_X1 U93367 ( .A(n81867), .ZN(n107616) );
  INV_X1 U93368 ( .A(n81860), .ZN(n107610) );
  INV_X1 U93369 ( .A(\DLX_Datapath/ArithLogUnit/B_add [11]), .ZN(n108507) );
  INV_X1 U93370 ( .A(\DLX_Datapath/ArithLogUnit/A_add [11]), .ZN(n108502) );
  INV_X1 U93371 ( .A(\DLX_Datapath/ArithLogUnit/B_add [27]), .ZN(n108047) );
  INV_X1 U93372 ( .A(\DLX_Datapath/ArithLogUnit/A_add [27]), .ZN(n110749) );
  INV_X1 U93373 ( .A(n81972), .ZN(n111125) );
  INV_X1 U93374 ( .A(n81833), .ZN(n107597) );
  INV_X1 U93375 ( .A(n82764), .ZN(n111144) );
  INV_X1 U93376 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [14]), .ZN(n108392) );
  INV_X1 U93377 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [12]), .ZN(n107740) );
  INV_X1 U93378 ( .A(\DLX_Datapath/ArithLogUnit/A_add [13]), .ZN(n109769) );
  INV_X1 U93379 ( .A(n81871), .ZN(n107618) );
  INV_X1 U93380 ( .A(n81872), .ZN(n107619) );
  INV_X1 U93381 ( .A(\DLX_Datapath/ArithLogUnit/A_add [5]), .ZN(n109315) );
  INV_X1 U93382 ( .A(\DLX_Datapath/ArithLogUnit/A_add [21]), .ZN(n110651) );
  INV_X1 U93383 ( .A(\DLX_Datapath/ArithLogUnit/A_add [29]), .ZN(n109772) );
  INV_X1 U93384 ( .A(n99943), .ZN(n107561) );
  INV_X1 U93385 ( .A(n100009), .ZN(n107563) );
  INV_X1 U93386 ( .A(n100040), .ZN(n107564) );
  INV_X1 U93387 ( .A(n99978), .ZN(n107562) );
  INV_X1 U93388 ( .A(n100131), .ZN(n107565) );
  INV_X1 U93389 ( .A(n100179), .ZN(n107567) );
  INV_X1 U93390 ( .A(n100158), .ZN(n107566) );
  INV_X1 U93391 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[0] ), .ZN(n107568) );
  INV_X1 U93392 ( .A(n81874), .ZN(n109892) );
  INV_X1 U93393 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[14] ), .ZN(
        n107502) );
  INV_X1 U93394 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/m_2A[8] ), .ZN(
        n107531) );
  INV_X1 U93395 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[17] ), .ZN(
        n108266) );
  INV_X1 U93396 ( .A(\DLX_Datapath/ArithLogUnit/A_add [9]), .ZN(n109764) );
  INV_X1 U93397 ( .A(\DLX_Datapath/ArithLogUnit/A_add [25]), .ZN(n110953) );
  INV_X1 U93398 ( .A(\DLX_Datapath/ArithLogUnit/A_add [30]), .ZN(n110955) );
  INV_X1 U93399 ( .A(n81822), .ZN(n107587) );
  INV_X1 U93400 ( .A(n81849), .ZN(n107600) );
  INV_X1 U93401 ( .A(n81869), .ZN(n107617) );
  INV_X1 U93402 ( .A(n81862), .ZN(n107611) );
  INV_X1 U93403 ( .A(n81858), .ZN(n107605) );
  INV_X1 U93404 ( .A(n81835), .ZN(n107598) );
  INV_X1 U93405 ( .A(n81831), .ZN(n107592) );
  CLKBUF_X1 U93406 ( .A(n79746), .Z(n105123) );
  INV_X1 U93407 ( .A(IR_in[30]), .ZN(n111141) );
  INV_X1 U93408 ( .A(\DLX_Datapath/ArithLogUnit/B_add [31]), .ZN(n107951) );
  INV_X1 U93409 ( .A(\DLX_Datapath/ArithLogUnit/A_add [31]), .ZN(n109771) );
  INV_X1 U93410 ( .A(IR_in[0]), .ZN(net67007) );
  INV_X1 U93411 ( .A(IR_in[28]), .ZN(n111143) );
  INV_X1 U93412 ( .A(\DLX_Datapath/ArithLogUnit/A_log [20]), .ZN(n110440) );
  INV_X1 U93413 ( .A(\DLX_Datapath/ArithLogUnit/A_log [16]), .ZN(n109896) );
  INV_X1 U93414 ( .A(\DLX_Datapath/ArithLogUnit/A_log [8]), .ZN(n109546) );
  INV_X1 U93415 ( .A(\DLX_Datapath/ArithLogUnit/A_log [4]), .ZN(n109205) );
  INV_X1 U93416 ( .A(\DLX_Datapath/ArithLogUnit/A_log [12]), .ZN(n107743) );
  INV_X1 U93417 ( .A(\DLX_Datapath/ArithLogUnit/A_log [24]), .ZN(n108157) );
  INV_X1 U93418 ( .A(\DLX_Datapath/ArithLogUnit/A_log [28]), .ZN(n107854) );
  INV_X1 U93419 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[3] ), .ZN(n108737) );
  INV_X1 U93420 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[5] ), .ZN(n109313) );
  INV_X1 U93421 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[7] ), .ZN(n109082) );
  INV_X1 U93422 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[9] ), .ZN(n109759) );
  INV_X1 U93423 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[1] ), .ZN(n108855) );
  INV_X1 U93424 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [7]), .ZN(n109089) );
  INV_X1 U93425 ( .A(n81846), .ZN(n109894) );
  INV_X1 U93426 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [5]), .ZN(n109310) );
  INV_X1 U93427 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [3]), .ZN(n108745) );
  INV_X1 U93428 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[2] ), .ZN(n108966) );
  INV_X1 U93429 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[4] ), .ZN(n109204) );
  INV_X1 U93430 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[6] ), .ZN(n109429) );
  INV_X1 U93431 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[8] ), .ZN(n109545) );
  INV_X1 U93432 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[10] ), .ZN(
        n108614) );
  INV_X1 U93433 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[11] ), .ZN(
        n109652) );
  INV_X1 U93434 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[12] ), .ZN(
        n107742) );
  INV_X1 U93435 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[13] ), .ZN(
        n108501) );
  INV_X1 U93436 ( .A(\DLX_Datapath/ArithLogUnit/ALU_mult/p_A[14] ), .ZN(
        n108389) );
  INV_X1 U93437 ( .A(n100292), .ZN(n106955) );
  INV_X1 U93438 ( .A(n86298), .ZN(n106941) );
  INV_X1 U93439 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [1]), .ZN(n108857) );
  INV_X1 U93440 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [9]), .ZN(n109762) );
  INV_X1 U93441 ( .A(IR_in[1]), .ZN(net67008) );
  INV_X1 U93442 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [11]), .ZN(n108505) );
  INV_X1 U93443 ( .A(\DLX_Datapath/ArithLogUnit/Cin_add ), .ZN(n107578) );
  INV_X1 U93444 ( .A(\DLX_Datapath/ArithLogUnit/A_add [19]), .ZN(n110118) );
  INV_X1 U93445 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [15]), .ZN(n108273) );
  INV_X1 U93446 ( .A(IR_in[4]), .ZN(n111158) );
  INV_X1 U93447 ( .A(\DLX_Datapath/ArithLogUnit/A_add [18]), .ZN(n110225) );
  INV_X1 U93448 ( .A(IR_in[31]), .ZN(n111123) );
  INV_X1 U93449 ( .A(IR_in[27]), .ZN(n111146) );
  INV_X1 U93450 ( .A(IR_in[26]), .ZN(n111149) );
  INV_X1 U93451 ( .A(IR_in[14]), .ZN(n111155) );
  INV_X1 U93452 ( .A(IR_in[15]), .ZN(n111154) );
  INV_X1 U93453 ( .A(IR_in[2]), .ZN(n111160) );
  INV_X1 U93454 ( .A(\DLX_Datapath/ArithLogUnit/B_add [18]), .ZN(n109781) );
  INV_X1 U93455 ( .A(\DLX_Datapath/ArithLogUnit/B_add [19]), .ZN(n109779) );
  INV_X1 U93456 ( .A(n99717), .ZN(n108268) );
  INV_X1 U93457 ( .A(n99014), .ZN(n108267) );
  INV_X1 U93458 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [2]), .ZN(n108968) );
  INV_X1 U93459 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [6]), .ZN(n109432) );
  INV_X1 U93460 ( .A(\DLX_Datapath/ArithLogUnit/A_log [31]), .ZN(n107949) );
  INV_X1 U93461 ( .A(\DLX_Datapath/ArithLogUnit/A_add [0]), .ZN(n108858) );
  INV_X1 U93462 ( .A(\DLX_Datapath/ArithLogUnit/A_log [21]), .ZN(n110650) );
  INV_X1 U93463 ( .A(\DLX_Datapath/ArithLogUnit/A_log [22]), .ZN(n110330) );
  INV_X1 U93464 ( .A(\DLX_Datapath/ArithLogUnit/A_log [23]), .ZN(n110545) );
  INV_X1 U93465 ( .A(\DLX_Datapath/ArithLogUnit/A_log [17]), .ZN(n110009) );
  INV_X1 U93466 ( .A(\DLX_Datapath/ArithLogUnit/A_log [18]), .ZN(n110224) );
  INV_X1 U93467 ( .A(\DLX_Datapath/ArithLogUnit/A_log [19]), .ZN(n110117) );
  INV_X1 U93468 ( .A(\DLX_Datapath/ArithLogUnit/A_log [9]), .ZN(n109760) );
  INV_X1 U93469 ( .A(\DLX_Datapath/ArithLogUnit/A_log [5]), .ZN(n109314) );
  INV_X1 U93470 ( .A(\DLX_Datapath/ArithLogUnit/A_log [6]), .ZN(n109430) );
  INV_X1 U93471 ( .A(\DLX_Datapath/ArithLogUnit/A_log [7]), .ZN(n109083) );
  INV_X1 U93472 ( .A(\DLX_Datapath/ArithLogUnit/A_log [2]), .ZN(n108967) );
  INV_X1 U93473 ( .A(\DLX_Datapath/ArithLogUnit/A_log [1]), .ZN(n108856) );
  INV_X1 U93474 ( .A(\DLX_Datapath/ArithLogUnit/A_log [3]), .ZN(n108738) );
  INV_X1 U93475 ( .A(\DLX_Datapath/ArithLogUnit/A_log [10]), .ZN(n109765) );
  INV_X1 U93476 ( .A(\DLX_Datapath/ArithLogUnit/A_log [11]), .ZN(n109653) );
  INV_X1 U93477 ( .A(\DLX_Datapath/ArithLogUnit/A_log [13]), .ZN(n109768) );
  INV_X1 U93478 ( .A(\DLX_Datapath/ArithLogUnit/A_log [14]), .ZN(n108390) );
  INV_X1 U93479 ( .A(\DLX_Datapath/ArithLogUnit/A_log [15]), .ZN(n108269) );
  INV_X1 U93480 ( .A(\DLX_Datapath/ArithLogUnit/A_log [25]), .ZN(n108156) );
  INV_X1 U93481 ( .A(\DLX_Datapath/ArithLogUnit/A_log [26]), .ZN(n108153) );
  INV_X1 U93482 ( .A(\DLX_Datapath/ArithLogUnit/A_log [27]), .ZN(n110748) );
  INV_X1 U93483 ( .A(\DLX_Datapath/ArithLogUnit/A_log [30]), .ZN(n108045) );
  INV_X1 U93484 ( .A(\DLX_Datapath/ArithLogUnit/A_log [29]), .ZN(n107572) );
  INV_X1 U93485 ( .A(\DLX_Datapath/ArithLogUnit/B_mul [4]), .ZN(n109202) );
  INV_X1 U93486 ( .A(\DLX_Datapath/ArithLogUnit/A_log [0]), .ZN(n107571) );
  INV_X1 U93487 ( .A(\DLX_Datapath/ArithLogUnit/B_add [0]), .ZN(n107620) );
  INV_X1 U93488 ( .A(\DLX_Datapath/ArithLogUnit/A_add [14]), .ZN(n109770) );
  INV_X1 U93489 ( .A(\DLX_Datapath/ArithLogUnit/A_add [2]), .ZN(n108969) );
  INV_X1 U93490 ( .A(\DLX_Datapath/ArithLogUnit/A_add [6]), .ZN(n109433) );
  INV_X1 U93491 ( .A(\DLX_Datapath/ArithLogUnit/A_add [22]), .ZN(n110331) );
  INV_X1 U93492 ( .A(n81875), .ZN(n109893) );
  INV_X1 U93493 ( .A(IR_in[12]), .ZN(n111156) );
  INV_X1 U93494 ( .A(IR_in[22]), .ZN(n111152) );
  INV_X1 U93495 ( .A(IR_in[29]), .ZN(n111142) );
  INV_X1 U93496 ( .A(IR_in[21]), .ZN(n111153) );
  INV_X1 U93497 ( .A(\DLX_Datapath/next_A_IDEX[1] ), .ZN(n108852) );
  INV_X1 U93498 ( .A(\DLX_Datapath/next_A_IDEX[0] ), .ZN(n107418) );
  INV_X1 U93499 ( .A(\DLX_Datapath/ArithLogUnit/B_log [21]), .ZN(n110653) );
  INV_X1 U93500 ( .A(\DLX_Datapath/ArithLogUnit/B_log [22]), .ZN(n110333) );
  INV_X1 U93501 ( .A(\DLX_Datapath/ArithLogUnit/B_log [23]), .ZN(n110227) );
  INV_X1 U93502 ( .A(\DLX_Datapath/ArithLogUnit/B_log [17]), .ZN(n110011) );
  INV_X1 U93503 ( .A(\DLX_Datapath/ArithLogUnit/B_log [18]), .ZN(n109780) );
  INV_X1 U93504 ( .A(\DLX_Datapath/ArithLogUnit/B_log [19]), .ZN(n109778) );
  INV_X1 U93505 ( .A(\DLX_Datapath/ArithLogUnit/B_log [9]), .ZN(n109763) );
  INV_X1 U93506 ( .A(\DLX_Datapath/ArithLogUnit/B_log [5]), .ZN(n109311) );
  INV_X1 U93507 ( .A(\DLX_Datapath/ArithLogUnit/B_log [6]), .ZN(n109434) );
  INV_X1 U93508 ( .A(\DLX_Datapath/ArithLogUnit/B_log [7]), .ZN(n109091) );
  INV_X1 U93509 ( .A(\DLX_Datapath/ArithLogUnit/B_log [2]), .ZN(n108970) );
  INV_X1 U93510 ( .A(\DLX_Datapath/ArithLogUnit/B_log [1]), .ZN(n108859) );
  INV_X1 U93511 ( .A(\DLX_Datapath/ArithLogUnit/B_log [3]), .ZN(n108746) );
  INV_X1 U93512 ( .A(\DLX_Datapath/ArithLogUnit/B_log [10]), .ZN(n109767) );
  INV_X1 U93513 ( .A(\DLX_Datapath/ArithLogUnit/B_log [11]), .ZN(n108506) );
  INV_X1 U93514 ( .A(\DLX_Datapath/ArithLogUnit/B_log [13]), .ZN(n109773) );
  INV_X1 U93515 ( .A(\DLX_Datapath/ArithLogUnit/B_log [14]), .ZN(n108393) );
  INV_X1 U93516 ( .A(\DLX_Datapath/ArithLogUnit/B_log [15]), .ZN(n108274) );
  INV_X1 U93517 ( .A(\DLX_Datapath/ArithLogUnit/B_log [25]), .ZN(n110954) );
  INV_X1 U93518 ( .A(\DLX_Datapath/ArithLogUnit/B_log [26]), .ZN(n108155) );
  INV_X1 U93519 ( .A(\DLX_Datapath/ArithLogUnit/B_log [27]), .ZN(n108046) );
  INV_X1 U93520 ( .A(\DLX_Datapath/ArithLogUnit/B_log [30]), .ZN(n110956) );
  INV_X1 U93521 ( .A(\DLX_Datapath/ArithLogUnit/B_log [31]), .ZN(n107950) );
  INV_X1 U93522 ( .A(\DLX_Datapath/ArithLogUnit/B_log [29]), .ZN(n107574) );
  INV_X1 U93523 ( .A(\DLX_Datapath/ArithLogUnit/B_log [0]), .ZN(n107573) );
  INV_X1 U93524 ( .A(IR_in[25]), .ZN(n111150) );
  INV_X1 U93525 ( .A(IR_in[23]), .ZN(n111151) );
  NAND2_X1 U93526 ( .A1(\DLX_Datapath/RegisterFile/N27074 ), .A2(n104328), 
        .ZN(n105064) );
  NAND2_X1 U93527 ( .A1(n82246), .A2(n105067), .ZN(n60297) );
  NOR2_X1 U93528 ( .A1(n105066), .A2(n82243), .ZN(n105067) );
  OR2_X1 U93529 ( .A1(n82329), .A2(n59478), .ZN(n105068) );
  INV_X1 U93530 ( .A(net2465245), .ZN(PC_out[2]) );
  INV_X1 U93531 ( .A(PC_out[0]), .ZN(n105072) );
  INV_X1 U93532 ( .A(\DLX_Datapath/NPC_adder/P4_SumGen/CSel_i_0/S_0[1] ), .ZN(
        n105073) );
  NOR2_X1 U93533 ( .A1(n105073), .A2(n105072), .ZN(n105074) );
  CLKBUF_X1 U93534 ( .A(n105032), .Z(n105076) );
  INV_X1 U93535 ( .A(n105052), .ZN(n81890) );
  INV_X1 U93536 ( .A(n59517), .ZN(n107106) );
  CLKBUF_X1 U93537 ( .A(n106595), .Z(n105162) );
  CLKBUF_X1 U93538 ( .A(n106595), .Z(n105163) );
  CLKBUF_X1 U93539 ( .A(n106595), .Z(n105164) );
  INV_X1 U93540 ( .A(n105151), .ZN(n106595) );
  INV_X1 U93541 ( .A(PC_out[2]), .ZN(n105078) );
  INV_X1 U93542 ( .A(IR_in[3]), .ZN(n111159) );
  INV_X1 U93543 ( .A(n104857), .ZN(n106813) );
  NAND2_X1 U93544 ( .A1(n82282), .A2(n105069), .ZN(n60294) );
  INV_X1 U93545 ( .A(n82434), .ZN(n106549) );
  INV_X1 U93546 ( .A(n82436), .ZN(n106548) );
  INV_X1 U93547 ( .A(n82437), .ZN(n106547) );
  INV_X1 U93548 ( .A(n82438), .ZN(n106546) );
  INV_X1 U93549 ( .A(n82443), .ZN(n106542) );
  INV_X1 U93550 ( .A(n82439), .ZN(n106545) );
  INV_X1 U93551 ( .A(n82440), .ZN(n106544) );
  INV_X1 U93552 ( .A(n82441), .ZN(n106543) );
  INV_X1 U93553 ( .A(n82445), .ZN(n106541) );
  INV_X1 U93554 ( .A(n82471), .ZN(n106530) );
  INV_X1 U93555 ( .A(n82451), .ZN(n106538) );
  INV_X1 U93556 ( .A(n82461), .ZN(n106534) );
  INV_X1 U93557 ( .A(n82453), .ZN(n106537) );
  INV_X1 U93558 ( .A(n82456), .ZN(n106536) );
  INV_X1 U93559 ( .A(n82459), .ZN(n106535) );
  INV_X1 U93560 ( .A(n82449), .ZN(n106539) );
  INV_X1 U93561 ( .A(n82447), .ZN(n106540) );
  INV_X1 U93562 ( .A(n82469), .ZN(n106531) );
  INV_X1 U93563 ( .A(n82464), .ZN(n106533) );
  INV_X1 U93564 ( .A(n82466), .ZN(n106532) );
  INV_X1 U93565 ( .A(n82474), .ZN(n106529) );
  INV_X1 U93566 ( .A(n82480), .ZN(n106526) );
  INV_X1 U93567 ( .A(n82498), .ZN(n106518) );
  INV_X1 U93568 ( .A(n82497), .ZN(n106519) );
  INV_X1 U93569 ( .A(n82493), .ZN(n106521) );
  INV_X1 U93570 ( .A(n82494), .ZN(n106520) );
  NAND2_X1 U93571 ( .A1(n105079), .A2(n82265), .ZN(n60295) );
  NOR2_X1 U93572 ( .A1(n105080), .A2(n82263), .ZN(n105079) );
  INV_X1 U93573 ( .A(n82491), .ZN(n106522) );
  INV_X1 U93574 ( .A(n82483), .ZN(n106525) );
  INV_X1 U93575 ( .A(n82486), .ZN(n106524) );
  INV_X1 U93576 ( .A(n82488), .ZN(n106523) );
  NAND2_X1 U93577 ( .A1(n82258), .A2(n104804), .ZN(n105081) );
  NOR2_X1 U93578 ( .A1(n105082), .A2(n104799), .ZN(n82296) );
  INV_X1 U93579 ( .A(n82479), .ZN(n106527) );
  INV_X1 U93580 ( .A(n82612), .ZN(n106769) );
  INV_X1 U93581 ( .A(n82476), .ZN(n106528) );
  INV_X1 U93582 ( .A(n82292), .ZN(n106770) );
  INV_X1 U93583 ( .A(n82300), .ZN(n110963) );
  NAND2_X1 U93584 ( .A1(n105085), .A2(n82306), .ZN(n105083) );
  NAND2_X1 U93585 ( .A1(n82309), .A2(n82308), .ZN(n105085) );
  INV_X1 U93586 ( .A(n105153), .ZN(n111132) );
  OR2_X1 U93587 ( .A1(n105086), .A2(n105087), .ZN(n82485) );
  OR2_X1 U93588 ( .A1(n59477), .A2(n82500), .ZN(n105087) );
  INV_X1 U93589 ( .A(n80136), .ZN(n106783) );
  OR2_X1 U93590 ( .A1(n82490), .A2(n59478), .ZN(n105088) );
  CLKBUF_X3 U93591 ( .A(n98091), .Z(n105124) );
  CLKBUF_X3 U93592 ( .A(n97575), .Z(n105125) );
  CLKBUF_X3 U93593 ( .A(n97062), .Z(n105127) );
  CLKBUF_X3 U93594 ( .A(n96561), .Z(n105129) );
  CLKBUF_X3 U93595 ( .A(n96014), .Z(n105131) );
  CLKBUF_X3 U93596 ( .A(n96014), .Z(n105132) );
  CLKBUF_X3 U93597 ( .A(n95452), .Z(n105133) );
  CLKBUF_X3 U93598 ( .A(n95452), .Z(n105134) );
  CLKBUF_X3 U93599 ( .A(n95170), .Z(n105135) );
  CLKBUF_X3 U93600 ( .A(n94295), .Z(n105136) );
  CLKBUF_X3 U93601 ( .A(n94295), .Z(n105137) );
  NOR2_X1 U93602 ( .A1(n109317), .A2(n59422), .ZN(n105145) );
  NOR2_X1 U93603 ( .A1(n109317), .A2(n108971), .ZN(n105146) );
  NOR2_X1 U93604 ( .A1(n59422), .A2(n59423), .ZN(n105147) );
  NOR2_X1 U93605 ( .A1(n59422), .A2(n59423), .ZN(n105148) );
  NOR2_X1 U93606 ( .A1(n108971), .A2(n59423), .ZN(n105149) );
  CLKBUF_X1 U93607 ( .A(n106745), .Z(n105170) );
  CLKBUF_X1 U93608 ( .A(n106746), .Z(n105173) );
  CLKBUF_X1 U93609 ( .A(n107022), .Z(n105206) );
  INV_X1 U93610 ( .A(n105554), .ZN(n105553) );
  CLKBUF_X1 U93611 ( .A(n94663), .Z(n105601) );
  INV_X1 U93612 ( .A(n105601), .ZN(n105602) );
  INV_X1 U93613 ( .A(n83163), .ZN(n105858) );
  INV_X1 U93614 ( .A(n83158), .ZN(n105864) );
  INV_X1 U93615 ( .A(n81651), .ZN(n105972) );
  INV_X1 U93616 ( .A(n81629), .ZN(n105993) );
  INV_X1 U93617 ( .A(n106012), .ZN(n106009) );
  INV_X1 U93618 ( .A(n81509), .ZN(n106047) );
  INV_X1 U93619 ( .A(n81501), .ZN(n106052) );
  INV_X1 U93620 ( .A(n81498), .ZN(n106057) );
  INV_X1 U93621 ( .A(n81451), .ZN(n106073) );
  INV_X1 U93622 ( .A(n81415), .ZN(n106097) );
  INV_X1 U93623 ( .A(n81408), .ZN(n106102) );
  INV_X1 U93624 ( .A(n81403), .ZN(n106107) );
  INV_X1 U93625 ( .A(n81398), .ZN(n106112) );
  INV_X1 U93626 ( .A(n81394), .ZN(n106117) );
  INV_X1 U93627 ( .A(n81383), .ZN(n106132) );
  INV_X1 U93628 ( .A(n81378), .ZN(n106139) );
  INV_X1 U93629 ( .A(n81358), .ZN(n106150) );
  INV_X1 U93630 ( .A(n81349), .ZN(n106161) );
  INV_X1 U93631 ( .A(n81345), .ZN(n106166) );
  INV_X1 U93632 ( .A(n81340), .ZN(n106174) );
  INV_X1 U93633 ( .A(n81318), .ZN(n106189) );
  INV_X1 U93634 ( .A(n81315), .ZN(n106194) );
  INV_X1 U93635 ( .A(n81310), .ZN(n106201) );
  INV_X1 U93636 ( .A(n81306), .ZN(n106207) );
  INV_X1 U93637 ( .A(n81299), .ZN(n106212) );
  INV_X1 U93638 ( .A(n81294), .ZN(n106222) );
  INV_X1 U93639 ( .A(n81284), .ZN(n106234) );
  INV_X1 U93640 ( .A(n81281), .ZN(n106239) );
  INV_X1 U93641 ( .A(n81278), .ZN(n106247) );
  INV_X1 U93642 ( .A(n81270), .ZN(n106258) );
  INV_X1 U93643 ( .A(n81267), .ZN(n106263) );
  INV_X1 U93644 ( .A(n81262), .ZN(n106270) );
  INV_X1 U93645 ( .A(n81250), .ZN(n106277) );
  INV_X1 U93646 ( .A(n81208), .ZN(n106280) );
  INV_X1 U93647 ( .A(n81199), .ZN(n106281) );
  CLKBUF_X1 U93648 ( .A(n80260), .Z(n106282) );
  CLKBUF_X1 U93649 ( .A(n80259), .Z(n106286) );
  INV_X1 U93650 ( .A(n106328), .ZN(n106327) );
  INV_X1 U93651 ( .A(n80203), .ZN(n106328) );
  INV_X1 U93652 ( .A(n80190), .ZN(n106334) );
  CLKBUF_X1 U93653 ( .A(n106361), .Z(n106367) );
  CLKBUF_X1 U93654 ( .A(\DLX_Datapath/ArithLogUnit/N178 ), .Z(n106370) );
  INV_X1 U93655 ( .A(n106511), .ZN(n106373) );
  INV_X1 U93656 ( .A(n106516), .ZN(n106374) );
  INV_X1 U93657 ( .A(n106516), .ZN(n106375) );
  INV_X1 U93658 ( .A(n106509), .ZN(n106376) );
  INV_X1 U93659 ( .A(n106515), .ZN(n106377) );
  INV_X1 U93660 ( .A(n106510), .ZN(n106378) );
  INV_X1 U93661 ( .A(n106510), .ZN(n106379) );
  INV_X1 U93662 ( .A(n106510), .ZN(n106380) );
  INV_X1 U93663 ( .A(n106510), .ZN(n106381) );
  INV_X1 U93664 ( .A(n106514), .ZN(n106382) );
  INV_X1 U93665 ( .A(n106509), .ZN(n106383) );
  INV_X1 U93666 ( .A(n106516), .ZN(n106384) );
  INV_X1 U93667 ( .A(n106510), .ZN(n106385) );
  INV_X1 U93668 ( .A(n106510), .ZN(n106386) );
  INV_X1 U93669 ( .A(n106515), .ZN(n106387) );
  INV_X1 U93670 ( .A(n106515), .ZN(n106388) );
  INV_X1 U93671 ( .A(n106515), .ZN(n106389) );
  INV_X1 U93672 ( .A(n106514), .ZN(n106390) );
  INV_X1 U93673 ( .A(n106512), .ZN(n106391) );
  INV_X1 U93674 ( .A(n106512), .ZN(n106392) );
  INV_X1 U93675 ( .A(n106512), .ZN(n106393) );
  INV_X1 U93676 ( .A(n106516), .ZN(n106394) );
  INV_X1 U93677 ( .A(n106514), .ZN(n106395) );
  INV_X1 U93678 ( .A(n106511), .ZN(n106396) );
  INV_X1 U93679 ( .A(n106513), .ZN(n106397) );
  INV_X1 U93680 ( .A(n106512), .ZN(n106398) );
  INV_X1 U93681 ( .A(n106509), .ZN(n106399) );
  INV_X1 U93682 ( .A(n106509), .ZN(n106400) );
  INV_X1 U93683 ( .A(n106512), .ZN(n106401) );
  INV_X1 U93684 ( .A(n106515), .ZN(n106402) );
  INV_X1 U93685 ( .A(n106515), .ZN(n106403) );
  INV_X1 U93686 ( .A(n106516), .ZN(n106404) );
  INV_X1 U93687 ( .A(n106510), .ZN(n106405) );
  INV_X1 U93688 ( .A(n106510), .ZN(n106406) );
  INV_X1 U93689 ( .A(n106515), .ZN(n106407) );
  INV_X1 U93690 ( .A(n106516), .ZN(n106408) );
  INV_X1 U93691 ( .A(n106512), .ZN(n106409) );
  INV_X1 U93692 ( .A(n106514), .ZN(n106410) );
  INV_X1 U93693 ( .A(n106512), .ZN(n106411) );
  INV_X1 U93694 ( .A(n106515), .ZN(n106412) );
  INV_X1 U93695 ( .A(n106510), .ZN(n106413) );
  INV_X1 U93696 ( .A(n106515), .ZN(n106414) );
  INV_X1 U93697 ( .A(n106516), .ZN(n106415) );
  INV_X1 U93698 ( .A(n106516), .ZN(n106416) );
  INV_X1 U93699 ( .A(n106516), .ZN(n106417) );
  INV_X1 U93700 ( .A(n106513), .ZN(n106418) );
  INV_X1 U93701 ( .A(n106514), .ZN(n106419) );
  INV_X1 U93702 ( .A(n106514), .ZN(n106420) );
  INV_X1 U93703 ( .A(n106514), .ZN(n106421) );
  INV_X1 U93704 ( .A(n106514), .ZN(n106422) );
  INV_X1 U93705 ( .A(n106512), .ZN(n106423) );
  INV_X1 U93706 ( .A(n106511), .ZN(n106424) );
  INV_X1 U93707 ( .A(n106513), .ZN(n106425) );
  INV_X1 U93708 ( .A(n106512), .ZN(n106426) );
  INV_X1 U93709 ( .A(n106516), .ZN(n106427) );
  INV_X1 U93710 ( .A(n106515), .ZN(n106428) );
  INV_X1 U93711 ( .A(n106513), .ZN(n106429) );
  INV_X1 U93712 ( .A(n106512), .ZN(n106430) );
  INV_X1 U93713 ( .A(n106511), .ZN(n106431) );
  INV_X1 U93714 ( .A(n106510), .ZN(n106432) );
  INV_X1 U93715 ( .A(n106510), .ZN(n106433) );
  INV_X1 U93716 ( .A(n106510), .ZN(n106434) );
  INV_X1 U93717 ( .A(n106511), .ZN(n106435) );
  INV_X1 U93718 ( .A(n106514), .ZN(n106436) );
  INV_X1 U93719 ( .A(n106510), .ZN(n106437) );
  INV_X1 U93720 ( .A(n106510), .ZN(n106438) );
  INV_X1 U93721 ( .A(n106510), .ZN(n106439) );
  INV_X1 U93722 ( .A(n106511), .ZN(n106440) );
  INV_X1 U93723 ( .A(n106513), .ZN(n106441) );
  INV_X1 U93724 ( .A(n106511), .ZN(n106442) );
  INV_X1 U93725 ( .A(n106513), .ZN(n106443) );
  INV_X1 U93726 ( .A(n106516), .ZN(n106444) );
  INV_X1 U93727 ( .A(n106510), .ZN(n106445) );
  INV_X1 U93728 ( .A(n106515), .ZN(n106446) );
  INV_X1 U93729 ( .A(n106516), .ZN(n106447) );
  INV_X1 U93730 ( .A(n106515), .ZN(n106448) );
  INV_X1 U93731 ( .A(n106514), .ZN(n106449) );
  INV_X1 U93732 ( .A(n106509), .ZN(n106450) );
  INV_X1 U93733 ( .A(n106509), .ZN(n106451) );
  INV_X1 U93734 ( .A(n106509), .ZN(n106452) );
  INV_X1 U93735 ( .A(n106509), .ZN(n106453) );
  INV_X1 U93736 ( .A(n106509), .ZN(n106454) );
  INV_X1 U93737 ( .A(n106512), .ZN(n106455) );
  INV_X1 U93738 ( .A(n106513), .ZN(n106456) );
  INV_X1 U93739 ( .A(n106511), .ZN(n106457) );
  INV_X1 U93740 ( .A(n106511), .ZN(n106458) );
  INV_X1 U93741 ( .A(n106509), .ZN(n106459) );
  INV_X1 U93742 ( .A(n106512), .ZN(n106460) );
  INV_X1 U93743 ( .A(n106509), .ZN(n106461) );
  INV_X1 U93744 ( .A(n106511), .ZN(n106462) );
  INV_X1 U93745 ( .A(n106511), .ZN(n106463) );
  INV_X1 U93746 ( .A(n106511), .ZN(n106464) );
  INV_X1 U93747 ( .A(n106512), .ZN(n106465) );
  INV_X1 U93748 ( .A(n106512), .ZN(n106466) );
  INV_X1 U93749 ( .A(n106513), .ZN(n106467) );
  INV_X1 U93750 ( .A(n106513), .ZN(n106468) );
  INV_X1 U93751 ( .A(n106513), .ZN(n106469) );
  INV_X1 U93752 ( .A(n106514), .ZN(n106470) );
  INV_X1 U93753 ( .A(n106514), .ZN(n106471) );
  INV_X1 U93754 ( .A(n106514), .ZN(n106472) );
  INV_X1 U93755 ( .A(n106511), .ZN(n106473) );
  INV_X1 U93756 ( .A(n106514), .ZN(n106474) );
  INV_X1 U93757 ( .A(n106511), .ZN(n106475) );
  INV_X1 U93758 ( .A(n106515), .ZN(n106476) );
  INV_X1 U93759 ( .A(n106516), .ZN(n106477) );
  INV_X1 U93760 ( .A(n106516), .ZN(n106478) );
  INV_X1 U93761 ( .A(n106512), .ZN(n106479) );
  INV_X1 U93762 ( .A(n106514), .ZN(n106480) );
  INV_X1 U93763 ( .A(n106514), .ZN(n106481) );
  INV_X1 U93764 ( .A(n106512), .ZN(n106482) );
  INV_X1 U93765 ( .A(n106512), .ZN(n106483) );
  INV_X1 U93766 ( .A(n106513), .ZN(n106484) );
  INV_X1 U93767 ( .A(n106512), .ZN(n106485) );
  INV_X1 U93768 ( .A(n106513), .ZN(n106486) );
  INV_X1 U93769 ( .A(n106509), .ZN(n106487) );
  INV_X1 U93770 ( .A(n106513), .ZN(n106488) );
  INV_X1 U93771 ( .A(n106512), .ZN(n106489) );
  INV_X1 U93772 ( .A(n106513), .ZN(n106490) );
  INV_X1 U93773 ( .A(n106512), .ZN(n106491) );
  INV_X1 U93774 ( .A(n106515), .ZN(n106492) );
  INV_X1 U93775 ( .A(n106513), .ZN(n106493) );
  INV_X1 U93776 ( .A(n106513), .ZN(n106494) );
  INV_X1 U93777 ( .A(n106510), .ZN(n106495) );
  INV_X1 U93778 ( .A(n106511), .ZN(n106496) );
  INV_X1 U93779 ( .A(n106513), .ZN(n106497) );
  INV_X1 U93780 ( .A(n106511), .ZN(n106498) );
  INV_X1 U93781 ( .A(n106511), .ZN(n106499) );
  INV_X1 U93782 ( .A(n106511), .ZN(n106500) );
  INV_X1 U93783 ( .A(n106512), .ZN(n106501) );
  INV_X1 U93784 ( .A(n106513), .ZN(n106502) );
  INV_X1 U93785 ( .A(n106512), .ZN(n106503) );
  INV_X1 U93786 ( .A(n106510), .ZN(n106504) );
  INV_X1 U93787 ( .A(n106512), .ZN(n106505) );
  INV_X1 U93788 ( .A(n106513), .ZN(n106506) );
  INV_X1 U93789 ( .A(n106512), .ZN(n106507) );
  INV_X1 U93790 ( .A(n106514), .ZN(n106508) );
  INV_X1 U93791 ( .A(Rst), .ZN(n106509) );
  INV_X1 U93792 ( .A(Rst), .ZN(n106510) );
  INV_X1 U93793 ( .A(Rst), .ZN(n106511) );
  INV_X1 U93794 ( .A(Rst), .ZN(n106512) );
  INV_X1 U93795 ( .A(Rst), .ZN(n106513) );
  INV_X1 U93796 ( .A(Rst), .ZN(n106514) );
  INV_X1 U93797 ( .A(Rst), .ZN(n106515) );
  INV_X1 U93798 ( .A(Rst), .ZN(n106516) );
endmodule

